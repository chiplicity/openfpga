magic
tech EFS8A
magscale 1 2
timestamp 1603801337
<< locali >>
rect 7665 12631 7699 12937
rect 6009 11543 6043 11645
rect 3893 8347 3927 8585
rect 11529 8347 11563 8449
rect 7021 2363 7055 2465
<< viali >>
rect 25053 23817 25087 23851
rect 13553 23681 13587 23715
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 13068 23613 13102 23647
rect 24660 23613 24694 23647
rect 1547 23477 1581 23511
rect 13139 23477 13173 23511
rect 24731 23477 24765 23511
rect 25053 22729 25087 22763
rect 24660 22525 24694 22559
rect 24731 22389 24765 22423
rect 12976 21437 13010 21471
rect 13461 21369 13495 21403
rect 13047 21301 13081 21335
rect 1476 20961 1510 20995
rect 2488 20961 2522 20995
rect 24660 20961 24694 20995
rect 1547 20825 1581 20859
rect 2559 20757 2593 20791
rect 24731 20757 24765 20791
rect 3249 20553 3283 20587
rect 24685 20553 24719 20587
rect 1547 20485 1581 20519
rect 1476 20349 1510 20383
rect 2237 20349 2271 20383
rect 2488 20349 2522 20383
rect 2973 20281 3007 20315
rect 1869 20213 1903 20247
rect 2559 20213 2593 20247
rect 1444 19873 1478 19907
rect 4144 19873 4178 19907
rect 2421 19805 2455 19839
rect 1547 19669 1581 19703
rect 4215 19669 4249 19703
rect 2237 19465 2271 19499
rect 1444 19261 1478 19295
rect 1869 19261 1903 19295
rect 2488 19261 2522 19295
rect 2973 19261 3007 19295
rect 3500 19261 3534 19295
rect 3893 19261 3927 19295
rect 4512 19261 4546 19295
rect 1547 19193 1581 19227
rect 2559 19125 2593 19159
rect 3571 19125 3605 19159
rect 4353 19125 4387 19159
rect 4583 19125 4617 19159
rect 4997 19125 5031 19159
rect 1476 18785 1510 18819
rect 2488 18785 2522 18819
rect 4112 18785 4146 18819
rect 5156 18785 5190 18819
rect 5227 18649 5261 18683
rect 1547 18581 1581 18615
rect 2559 18581 2593 18615
rect 4215 18581 4249 18615
rect 1961 18377 1995 18411
rect 3341 18377 3375 18411
rect 4261 18309 4295 18343
rect 5181 18241 5215 18275
rect 1444 18173 1478 18207
rect 2488 18173 2522 18207
rect 2881 18173 2915 18207
rect 3500 18173 3534 18207
rect 4480 18173 4514 18207
rect 5508 18173 5542 18207
rect 6929 18173 6963 18207
rect 2237 18105 2271 18139
rect 5595 18105 5629 18139
rect 7481 18105 7515 18139
rect 1547 18037 1581 18071
rect 2559 18037 2593 18071
rect 3571 18037 3605 18071
rect 3893 18037 3927 18071
rect 4583 18037 4617 18071
rect 5917 18037 5951 18071
rect 7113 18037 7147 18071
rect 1961 17697 1995 17731
rect 2145 17697 2179 17731
rect 4420 17697 4454 17731
rect 6168 17697 6202 17731
rect 8284 17697 8318 17731
rect 9756 17697 9790 17731
rect 2237 17629 2271 17663
rect 7205 17629 7239 17663
rect 10701 17629 10735 17663
rect 2789 17493 2823 17527
rect 4491 17493 4525 17527
rect 6239 17493 6273 17527
rect 8355 17493 8389 17527
rect 9827 17493 9861 17527
rect 6193 17289 6227 17323
rect 3065 17221 3099 17255
rect 1961 17085 1995 17119
rect 2145 17085 2179 17119
rect 3284 17085 3318 17119
rect 3709 17085 3743 17119
rect 4972 17085 5006 17119
rect 7180 17085 7214 17119
rect 8125 17085 8159 17119
rect 9648 17085 9682 17119
rect 10425 17085 10459 17119
rect 10676 17085 10710 17119
rect 11069 17085 11103 17119
rect 13068 17085 13102 17119
rect 13461 17085 13495 17119
rect 15025 17085 15059 17119
rect 15485 17085 15519 17119
rect 2789 17017 2823 17051
rect 7573 17017 7607 17051
rect 9045 17017 9079 17051
rect 9735 17017 9769 17051
rect 1777 16949 1811 16983
rect 3387 16949 3421 16983
rect 4445 16949 4479 16983
rect 5043 16949 5077 16983
rect 5365 16949 5399 16983
rect 7251 16949 7285 16983
rect 8309 16949 8343 16983
rect 8677 16949 8711 16983
rect 10057 16949 10091 16983
rect 10747 16949 10781 16983
rect 13139 16949 13173 16983
rect 15209 16949 15243 16983
rect 1777 16745 1811 16779
rect 4721 16745 4755 16779
rect 9781 16745 9815 16779
rect 13277 16745 13311 16779
rect 15485 16745 15519 16779
rect 16221 16745 16255 16779
rect 16497 16745 16531 16779
rect 2237 16677 2271 16711
rect 2329 16677 2363 16711
rect 8631 16677 8665 16711
rect 10793 16677 10827 16711
rect 4128 16609 4162 16643
rect 4215 16609 4249 16643
rect 5140 16609 5174 16643
rect 5227 16609 5261 16643
rect 6561 16609 6595 16643
rect 8528 16609 8562 16643
rect 9229 16609 9263 16643
rect 9965 16609 9999 16643
rect 10241 16609 10275 16643
rect 11713 16609 11747 16643
rect 11989 16609 12023 16643
rect 12173 16609 12207 16643
rect 13001 16609 13035 16643
rect 13553 16609 13587 16643
rect 15301 16609 15335 16643
rect 16313 16609 16347 16643
rect 2881 16541 2915 16575
rect 6745 16405 6779 16439
rect 12449 16405 12483 16439
rect 14197 16405 14231 16439
rect 3617 16201 3651 16235
rect 4629 16201 4663 16235
rect 8953 16201 8987 16235
rect 10149 16201 10183 16235
rect 12173 16201 12207 16235
rect 25053 16201 25087 16235
rect 2605 16065 2639 16099
rect 2881 16065 2915 16099
rect 4813 16065 4847 16099
rect 5089 16065 5123 16099
rect 14657 16065 14691 16099
rect 16221 16065 16255 16099
rect 7180 15997 7214 16031
rect 8160 15997 8194 16031
rect 8585 15997 8619 16031
rect 9137 15997 9171 16031
rect 9689 15997 9723 16031
rect 10701 15997 10735 16031
rect 11253 15997 11287 16031
rect 12541 15997 12575 16031
rect 13001 15997 13035 16031
rect 14289 15997 14323 16031
rect 14565 15997 14599 16031
rect 18061 15997 18095 16031
rect 24660 15997 24694 16031
rect 1501 15929 1535 15963
rect 2329 15929 2363 15963
rect 2697 15929 2731 15963
rect 4905 15929 4939 15963
rect 10517 15929 10551 15963
rect 11437 15929 11471 15963
rect 13461 15929 13495 15963
rect 15945 15929 15979 15963
rect 16313 15929 16347 15963
rect 16865 15929 16899 15963
rect 1961 15861 1995 15895
rect 4169 15861 4203 15895
rect 5825 15861 5859 15895
rect 6653 15861 6687 15895
rect 7251 15861 7285 15895
rect 7665 15861 7699 15895
rect 8263 15861 8297 15895
rect 9413 15861 9447 15895
rect 11805 15861 11839 15895
rect 12541 15861 12575 15895
rect 14013 15861 14047 15895
rect 15393 15861 15427 15895
rect 17141 15861 17175 15895
rect 18245 15861 18279 15895
rect 18613 15861 18647 15895
rect 19073 15861 19107 15895
rect 24731 15861 24765 15895
rect 1685 15657 1719 15691
rect 3157 15657 3191 15691
rect 9137 15657 9171 15691
rect 11805 15657 11839 15691
rect 2329 15589 2363 15623
rect 2881 15589 2915 15623
rect 3525 15589 3559 15623
rect 4261 15589 4295 15623
rect 6101 15589 6135 15623
rect 6193 15589 6227 15623
rect 10333 15589 10367 15623
rect 13829 15589 13863 15623
rect 16313 15589 16347 15623
rect 17785 15589 17819 15623
rect 17877 15589 17911 15623
rect 8033 15521 8067 15555
rect 8493 15521 8527 15555
rect 11897 15521 11931 15555
rect 12265 15521 12299 15555
rect 2053 15453 2087 15487
rect 2237 15453 2271 15487
rect 4169 15453 4203 15487
rect 4813 15453 4847 15487
rect 6377 15453 6411 15487
rect 7021 15453 7055 15487
rect 8769 15453 8803 15487
rect 10241 15453 10275 15487
rect 13737 15453 13771 15487
rect 16221 15453 16255 15487
rect 16865 15453 16899 15487
rect 18061 15453 18095 15487
rect 19441 15453 19475 15487
rect 21557 15453 21591 15487
rect 9873 15385 9907 15419
rect 10793 15385 10827 15419
rect 13093 15385 13127 15419
rect 14289 15385 14323 15419
rect 11437 15317 11471 15351
rect 13369 15317 13403 15351
rect 14657 15317 14691 15351
rect 15761 15317 15795 15351
rect 1961 15113 1995 15147
rect 5733 15113 5767 15147
rect 10241 15113 10275 15147
rect 12265 15113 12299 15147
rect 13645 15113 13679 15147
rect 15209 15113 15243 15147
rect 17417 15113 17451 15147
rect 2329 15045 2363 15079
rect 3709 15045 3743 15079
rect 4077 15045 4111 15079
rect 19625 15045 19659 15079
rect 2789 14977 2823 15011
rect 4353 14977 4387 15011
rect 5273 14977 5307 15011
rect 6929 14977 6963 15011
rect 7205 14977 7239 15011
rect 10885 14977 10919 15011
rect 12633 14977 12667 15011
rect 14197 14977 14231 15011
rect 16037 14977 16071 15011
rect 17785 14977 17819 15011
rect 1476 14909 1510 14943
rect 8861 14909 8895 14943
rect 9413 14909 9447 14943
rect 18061 14909 18095 14943
rect 19073 14909 19107 14943
rect 20152 14909 20186 14943
rect 21316 14909 21350 14943
rect 21741 14909 21775 14943
rect 23832 14909 23866 14943
rect 24777 14909 24811 14943
rect 2881 14841 2915 14875
rect 3433 14841 3467 14875
rect 4445 14841 4479 14875
rect 4997 14841 5031 14875
rect 7021 14841 7055 14875
rect 9597 14841 9631 14875
rect 10977 14841 11011 14875
rect 11529 14841 11563 14875
rect 12725 14841 12759 14875
rect 13277 14841 13311 14875
rect 14289 14841 14323 14875
rect 14841 14841 14875 14875
rect 15761 14841 15795 14875
rect 15853 14841 15887 14875
rect 1547 14773 1581 14807
rect 6101 14773 6135 14807
rect 6653 14773 6687 14807
rect 8033 14773 8067 14807
rect 8677 14773 8711 14807
rect 10701 14773 10735 14807
rect 11897 14773 11931 14807
rect 15485 14773 15519 14807
rect 16681 14773 16715 14807
rect 18245 14773 18279 14807
rect 18521 14773 18555 14807
rect 19257 14773 19291 14807
rect 20223 14773 20257 14807
rect 20545 14773 20579 14807
rect 21419 14773 21453 14807
rect 22293 14773 22327 14807
rect 23903 14773 23937 14807
rect 24317 14773 24351 14807
rect 1961 14569 1995 14603
rect 2973 14569 3007 14603
rect 3249 14569 3283 14603
rect 3893 14569 3927 14603
rect 6929 14569 6963 14603
rect 7941 14569 7975 14603
rect 9137 14569 9171 14603
rect 12357 14569 12391 14603
rect 14105 14569 14139 14603
rect 14381 14569 14415 14603
rect 15439 14569 15473 14603
rect 16221 14569 16255 14603
rect 17969 14569 18003 14603
rect 2374 14501 2408 14535
rect 4261 14501 4295 14535
rect 4813 14501 4847 14535
rect 6330 14501 6364 14535
rect 10051 14501 10085 14535
rect 11758 14501 11792 14535
rect 13547 14501 13581 14535
rect 16497 14501 16531 14535
rect 2053 14433 2087 14467
rect 8309 14433 8343 14467
rect 8585 14433 8619 14467
rect 9689 14433 9723 14467
rect 11437 14433 11471 14467
rect 13185 14433 13219 14467
rect 15368 14433 15402 14467
rect 17877 14433 17911 14467
rect 18337 14433 18371 14467
rect 19568 14433 19602 14467
rect 20948 14433 20982 14467
rect 21992 14433 22026 14467
rect 23984 14433 24018 14467
rect 24996 14433 25030 14467
rect 4169 14365 4203 14399
rect 6009 14365 6043 14399
rect 8769 14365 8803 14399
rect 16405 14365 16439 14399
rect 17049 14365 17083 14399
rect 22937 14365 22971 14399
rect 10885 14297 10919 14331
rect 5181 14229 5215 14263
rect 10609 14229 10643 14263
rect 11253 14229 11287 14263
rect 12725 14229 12759 14263
rect 13001 14229 13035 14263
rect 19671 14229 19705 14263
rect 21051 14229 21085 14263
rect 22063 14229 22097 14263
rect 24087 14229 24121 14263
rect 25099 14229 25133 14263
rect 2973 14025 3007 14059
rect 4629 14025 4663 14059
rect 7757 14025 7791 14059
rect 8125 14025 8159 14059
rect 8493 14025 8527 14059
rect 8723 14025 8757 14059
rect 11805 14025 11839 14059
rect 13369 14025 13403 14059
rect 15393 14025 15427 14059
rect 16405 14025 16439 14059
rect 16681 14025 16715 14059
rect 17417 14025 17451 14059
rect 20085 14025 20119 14059
rect 21465 14025 21499 14059
rect 22109 14025 22143 14059
rect 25421 14025 25455 14059
rect 3617 13957 3651 13991
rect 10609 13957 10643 13991
rect 10885 13957 10919 13991
rect 14013 13957 14047 13991
rect 17141 13957 17175 13991
rect 19809 13957 19843 13991
rect 25053 13957 25087 13991
rect 2053 13889 2087 13923
rect 3939 13889 3973 13923
rect 5273 13889 5307 13923
rect 5917 13889 5951 13923
rect 9689 13889 9723 13923
rect 12449 13889 12483 13923
rect 15025 13889 15059 13923
rect 15485 13889 15519 13923
rect 24731 13889 24765 13923
rect 3836 13821 3870 13855
rect 4261 13821 4295 13855
rect 6833 13821 6867 13855
rect 8620 13821 8654 13855
rect 9045 13821 9079 13855
rect 17785 13821 17819 13855
rect 18153 13821 18187 13855
rect 18797 13821 18831 13855
rect 19625 13821 19659 13855
rect 20453 13821 20487 13855
rect 20688 13821 20722 13855
rect 20775 13821 20809 13855
rect 21716 13821 21750 13855
rect 22569 13821 22603 13855
rect 23949 13821 23983 13855
rect 24644 13821 24678 13855
rect 2374 13753 2408 13787
rect 3249 13753 3283 13787
rect 5365 13753 5399 13787
rect 6285 13753 6319 13787
rect 6653 13753 6687 13787
rect 7199 13753 7233 13787
rect 9597 13753 9631 13787
rect 10051 13753 10085 13787
rect 12770 13753 12804 13787
rect 13645 13753 13679 13787
rect 14197 13753 14231 13787
rect 15806 13753 15840 13787
rect 1961 13685 1995 13719
rect 5089 13685 5123 13719
rect 11437 13685 11471 13719
rect 12173 13685 12207 13719
rect 21097 13685 21131 13719
rect 21787 13685 21821 13719
rect 25605 13685 25639 13719
rect 3065 13481 3099 13515
rect 4537 13481 4571 13515
rect 5089 13481 5123 13515
rect 6377 13481 6411 13515
rect 6653 13481 6687 13515
rect 7297 13481 7331 13515
rect 9505 13481 9539 13515
rect 16957 13481 16991 13515
rect 17325 13481 17359 13515
rect 18613 13481 18647 13515
rect 19211 13481 19245 13515
rect 2466 13413 2500 13447
rect 5819 13413 5853 13447
rect 10241 13413 10275 13447
rect 10333 13413 10367 13447
rect 13829 13413 13863 13447
rect 16129 13413 16163 13447
rect 17693 13413 17727 13447
rect 4144 13345 4178 13379
rect 7481 13345 7515 13379
rect 7665 13345 7699 13379
rect 12541 13345 12575 13379
rect 19140 13345 19174 13379
rect 20980 13345 21014 13379
rect 22636 13345 22670 13379
rect 23616 13345 23650 13379
rect 24628 13345 24662 13379
rect 2145 13277 2179 13311
rect 5457 13277 5491 13311
rect 10885 13277 10919 13311
rect 12817 13277 12851 13311
rect 13737 13277 13771 13311
rect 14013 13277 14047 13311
rect 16037 13277 16071 13311
rect 16313 13277 16347 13311
rect 17601 13277 17635 13311
rect 18245 13277 18279 13311
rect 4215 13209 4249 13243
rect 24731 13209 24765 13243
rect 1777 13141 1811 13175
rect 7113 13141 7147 13175
rect 9873 13141 9907 13175
rect 15485 13141 15519 13175
rect 21051 13141 21085 13175
rect 22707 13141 22741 13175
rect 23719 13141 23753 13175
rect 3249 12937 3283 12971
rect 4537 12937 4571 12971
rect 6101 12937 6135 12971
rect 7665 12937 7699 12971
rect 7941 12937 7975 12971
rect 8907 12937 8941 12971
rect 11161 12937 11195 12971
rect 13737 12937 13771 12971
rect 15301 12937 15335 12971
rect 16773 12937 16807 12971
rect 17601 12937 17635 12971
rect 20177 12937 20211 12971
rect 21649 12937 21683 12971
rect 23397 12937 23431 12971
rect 23857 12937 23891 12971
rect 24409 12937 24443 12971
rect 25145 12937 25179 12971
rect 4077 12869 4111 12903
rect 3525 12801 3559 12835
rect 5089 12801 5123 12835
rect 7297 12801 7331 12835
rect 1869 12733 1903 12767
rect 2237 12733 2271 12767
rect 2421 12733 2455 12767
rect 6653 12733 6687 12767
rect 7021 12733 7055 12767
rect 7389 12733 7423 12767
rect 3617 12665 3651 12699
rect 5181 12665 5215 12699
rect 5733 12665 5767 12699
rect 10885 12869 10919 12903
rect 11483 12801 11517 12835
rect 14565 12801 14599 12835
rect 15853 12801 15887 12835
rect 16313 12801 16347 12835
rect 18521 12801 18555 12835
rect 8804 12733 8838 12767
rect 9229 12733 9263 12767
rect 11380 12733 11414 12767
rect 12265 12733 12299 12767
rect 12541 12733 12575 12767
rect 17233 12733 17267 12767
rect 18061 12733 18095 12767
rect 18153 12733 18187 12767
rect 18337 12733 18371 12767
rect 19692 12733 19726 12767
rect 20856 12733 20890 12767
rect 21281 12733 21315 12767
rect 22636 12733 22670 12767
rect 24593 12733 24627 12767
rect 9873 12665 9907 12699
rect 9965 12665 9999 12699
rect 10517 12665 10551 12699
rect 11897 12665 11931 12699
rect 13185 12665 13219 12699
rect 14289 12665 14323 12699
rect 14381 12665 14415 12699
rect 15945 12665 15979 12699
rect 23121 12665 23155 12699
rect 2697 12597 2731 12631
rect 4905 12597 4939 12631
rect 7665 12597 7699 12631
rect 8585 12597 8619 12631
rect 9689 12597 9723 12631
rect 14105 12597 14139 12631
rect 15577 12597 15611 12631
rect 19165 12597 19199 12631
rect 19763 12597 19797 12631
rect 20959 12597 20993 12631
rect 22707 12597 22741 12631
rect 24777 12597 24811 12631
rect 3065 12393 3099 12427
rect 3525 12393 3559 12427
rect 5549 12393 5583 12427
rect 5733 12393 5767 12427
rect 9505 12393 9539 12427
rect 10609 12393 10643 12427
rect 13737 12393 13771 12427
rect 14657 12393 14691 12427
rect 18613 12393 18647 12427
rect 2145 12325 2179 12359
rect 2237 12325 2271 12359
rect 4261 12325 4295 12359
rect 10051 12325 10085 12359
rect 12449 12325 12483 12359
rect 13001 12325 13035 12359
rect 16221 12325 16255 12359
rect 17785 12325 17819 12359
rect 5917 12257 5951 12291
rect 6101 12257 6135 12291
rect 6837 12257 6871 12291
rect 7205 12257 7239 12291
rect 7757 12257 7791 12291
rect 8033 12257 8067 12291
rect 14197 12257 14231 12291
rect 19257 12257 19291 12291
rect 20948 12257 20982 12291
rect 22268 12257 22302 12291
rect 23740 12257 23774 12291
rect 24752 12257 24786 12291
rect 2789 12189 2823 12223
rect 4169 12189 4203 12223
rect 4813 12189 4847 12223
rect 8125 12189 8159 12223
rect 9689 12189 9723 12223
rect 10885 12189 10919 12223
rect 12357 12189 12391 12223
rect 16129 12189 16163 12223
rect 16773 12189 16807 12223
rect 17693 12189 17727 12223
rect 17969 12189 18003 12223
rect 14381 12121 14415 12155
rect 22339 12121 22373 12155
rect 1777 12053 1811 12087
rect 12081 12053 12115 12087
rect 15853 12053 15887 12087
rect 17509 12053 17543 12087
rect 19441 12053 19475 12087
rect 21051 12053 21085 12087
rect 23811 12053 23845 12087
rect 24823 12053 24857 12087
rect 1593 11849 1627 11883
rect 2053 11849 2087 11883
rect 5273 11849 5307 11883
rect 6561 11849 6595 11883
rect 10609 11849 10643 11883
rect 15945 11849 15979 11883
rect 16221 11849 16255 11883
rect 16681 11849 16715 11883
rect 19073 11849 19107 11883
rect 19441 11849 19475 11883
rect 22293 11849 22327 11883
rect 25145 11849 25179 11883
rect 3157 11781 3191 11815
rect 5641 11781 5675 11815
rect 5917 11781 5951 11815
rect 8309 11781 8343 11815
rect 10333 11781 10367 11815
rect 11437 11781 11471 11815
rect 24501 11781 24535 11815
rect 2237 11713 2271 11747
rect 3801 11713 3835 11747
rect 6929 11713 6963 11747
rect 9413 11713 9447 11747
rect 12725 11713 12759 11747
rect 15025 11713 15059 11747
rect 18153 11713 18187 11747
rect 18429 11713 18463 11747
rect 19717 11713 19751 11747
rect 5733 11645 5767 11679
rect 6009 11645 6043 11679
rect 8436 11645 8470 11679
rect 11253 11645 11287 11679
rect 14289 11645 14323 11679
rect 16773 11645 16807 11679
rect 17233 11645 17267 11679
rect 21281 11645 21315 11679
rect 23719 11645 23753 11679
rect 24133 11645 24167 11679
rect 24752 11645 24786 11679
rect 25513 11645 25547 11679
rect 2329 11577 2363 11611
rect 2881 11577 2915 11611
rect 3893 11577 3927 11611
rect 4445 11577 4479 11611
rect 7021 11577 7055 11611
rect 7573 11577 7607 11611
rect 8539 11577 8573 11611
rect 9734 11577 9768 11611
rect 13046 11577 13080 11611
rect 14933 11577 14967 11611
rect 15346 11577 15380 11611
rect 17877 11577 17911 11611
rect 18245 11577 18279 11611
rect 19809 11577 19843 11611
rect 20361 11577 20395 11611
rect 3617 11509 3651 11543
rect 4721 11509 4755 11543
rect 6009 11509 6043 11543
rect 6285 11509 6319 11543
rect 7849 11509 7883 11543
rect 8953 11509 8987 11543
rect 9321 11509 9355 11543
rect 11713 11509 11747 11543
rect 12265 11509 12299 11543
rect 13645 11509 13679 11543
rect 16957 11509 16991 11543
rect 20913 11509 20947 11543
rect 21649 11509 21683 11543
rect 23811 11509 23845 11543
rect 24823 11509 24857 11543
rect 1547 11305 1581 11339
rect 2237 11305 2271 11339
rect 3801 11305 3835 11339
rect 4261 11305 4295 11339
rect 5733 11305 5767 11339
rect 7389 11305 7423 11339
rect 9505 11305 9539 11339
rect 12541 11305 12575 11339
rect 12817 11305 12851 11339
rect 15025 11305 15059 11339
rect 16313 11305 16347 11339
rect 18153 11305 18187 11339
rect 18429 11305 18463 11339
rect 19993 11305 20027 11339
rect 21281 11305 21315 11339
rect 2513 11237 2547 11271
rect 2605 11237 2639 11271
rect 4813 11237 4847 11271
rect 5365 11237 5399 11271
rect 6555 11237 6589 11271
rect 8217 11237 8251 11271
rect 10010 11237 10044 11271
rect 11983 11237 12017 11271
rect 13185 11237 13219 11271
rect 13829 11237 13863 11271
rect 14381 11237 14415 11271
rect 15485 11237 15519 11271
rect 17554 11237 17588 11271
rect 18889 11237 18923 11271
rect 19165 11237 19199 11271
rect 19717 11237 19751 11271
rect 21741 11237 21775 11271
rect 1476 11169 1510 11203
rect 7113 11169 7147 11203
rect 9689 11169 9723 11203
rect 11621 11169 11655 11203
rect 23616 11169 23650 11203
rect 24593 11169 24627 11203
rect 4721 11101 4755 11135
rect 6193 11101 6227 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 8769 11101 8803 11135
rect 13737 11101 13771 11135
rect 15393 11101 15427 11135
rect 15669 11101 15703 11135
rect 17049 11101 17083 11135
rect 17233 11101 17267 11135
rect 19073 11101 19107 11135
rect 20361 11101 20395 11135
rect 21649 11101 21683 11135
rect 3065 11033 3099 11067
rect 6101 11033 6135 11067
rect 22201 11033 22235 11067
rect 23719 11033 23753 11067
rect 10609 10965 10643 10999
rect 24777 10965 24811 10999
rect 1685 10761 1719 10795
rect 3065 10761 3099 10795
rect 4813 10761 4847 10795
rect 9689 10761 9723 10795
rect 11989 10761 12023 10795
rect 13277 10761 13311 10795
rect 15393 10761 15427 10795
rect 16037 10761 16071 10795
rect 17141 10761 17175 10795
rect 21005 10761 21039 10795
rect 21465 10761 21499 10795
rect 22569 10761 22603 10795
rect 23029 10761 23063 10795
rect 24685 10761 24719 10795
rect 3341 10693 3375 10727
rect 4537 10693 4571 10727
rect 10609 10693 10643 10727
rect 20729 10693 20763 10727
rect 5273 10625 5307 10659
rect 5917 10625 5951 10659
rect 10057 10625 10091 10659
rect 14105 10625 14139 10659
rect 15025 10625 15059 10659
rect 18153 10625 18187 10659
rect 21649 10625 21683 10659
rect 21925 10625 21959 10659
rect 2145 10557 2179 10591
rect 3893 10557 3927 10591
rect 6653 10557 6687 10591
rect 7113 10557 7147 10591
rect 7389 10557 7423 10591
rect 8309 10557 8343 10591
rect 8677 10557 8711 10591
rect 8861 10557 8895 10591
rect 16221 10557 16255 10591
rect 18061 10557 18095 10591
rect 18337 10557 18371 10591
rect 19809 10557 19843 10591
rect 23489 10557 23523 10591
rect 23765 10557 23799 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 2053 10489 2087 10523
rect 2466 10489 2500 10523
rect 5365 10489 5399 10523
rect 10149 10489 10183 10523
rect 12725 10489 12759 10523
rect 13553 10489 13587 10523
rect 13829 10489 13863 10523
rect 13921 10489 13955 10523
rect 16542 10489 16576 10523
rect 17417 10489 17451 10523
rect 20171 10489 20205 10523
rect 21741 10489 21775 10523
rect 24409 10489 24443 10523
rect 3709 10421 3743 10455
rect 4077 10421 4111 10455
rect 6193 10421 6227 10455
rect 6929 10421 6963 10455
rect 7849 10421 7883 10455
rect 8493 10421 8527 10455
rect 11069 10421 11103 10455
rect 11713 10421 11747 10455
rect 15761 10421 15795 10455
rect 17785 10421 17819 10455
rect 18521 10421 18555 10455
rect 19349 10421 19383 10455
rect 19717 10421 19751 10455
rect 25421 10421 25455 10455
rect 2881 10217 2915 10251
rect 3157 10217 3191 10251
rect 3893 10217 3927 10251
rect 5549 10217 5583 10251
rect 7665 10217 7699 10251
rect 8585 10217 8619 10251
rect 9413 10217 9447 10251
rect 10701 10217 10735 10251
rect 11529 10217 11563 10251
rect 13369 10217 13403 10251
rect 14381 10217 14415 10251
rect 15393 10217 15427 10251
rect 17509 10217 17543 10251
rect 18797 10217 18831 10251
rect 21557 10217 21591 10251
rect 24317 10217 24351 10251
rect 2323 10149 2357 10183
rect 4261 10149 4295 10183
rect 4813 10149 4847 10183
rect 6187 10149 6221 10183
rect 7113 10149 7147 10183
rect 9873 10149 9907 10183
rect 12541 10149 12575 10183
rect 21925 10149 21959 10183
rect 23489 10149 23523 10183
rect 24961 10149 24995 10183
rect 25053 10149 25087 10183
rect 5273 10081 5307 10115
rect 6745 10081 6779 10115
rect 7757 10081 7791 10115
rect 8125 10081 8159 10115
rect 11345 10081 11379 10115
rect 13829 10081 13863 10115
rect 13988 10081 14022 10115
rect 15301 10081 15335 10115
rect 15761 10081 15795 10115
rect 16957 10081 16991 10115
rect 17141 10081 17175 10115
rect 19809 10081 19843 10115
rect 19993 10081 20027 10115
rect 1961 10013 1995 10047
rect 4169 10013 4203 10047
rect 5825 10013 5859 10047
rect 9781 10013 9815 10047
rect 11897 10013 11931 10047
rect 12449 10013 12483 10047
rect 21833 10013 21867 10047
rect 23397 10013 23431 10047
rect 23673 10013 23707 10047
rect 25237 10013 25271 10047
rect 10333 9945 10367 9979
rect 13001 9945 13035 9979
rect 18521 9945 18555 9979
rect 22385 9945 22419 9979
rect 12173 9877 12207 9911
rect 14059 9877 14093 9911
rect 16405 9877 16439 9911
rect 18061 9877 18095 9911
rect 20453 9877 20487 9911
rect 8217 9673 8251 9707
rect 13921 9673 13955 9707
rect 15301 9673 15335 9707
rect 24961 9673 24995 9707
rect 3065 9605 3099 9639
rect 3801 9605 3835 9639
rect 4537 9605 4571 9639
rect 9229 9605 9263 9639
rect 10333 9605 10367 9639
rect 11391 9605 11425 9639
rect 11805 9605 11839 9639
rect 13093 9605 13127 9639
rect 15669 9605 15703 9639
rect 19533 9605 19567 9639
rect 21373 9605 21407 9639
rect 21741 9605 21775 9639
rect 23397 9605 23431 9639
rect 2145 9537 2179 9571
rect 3433 9537 3467 9571
rect 5273 9537 5307 9571
rect 5917 9537 5951 9571
rect 12541 9537 12575 9571
rect 13553 9537 13587 9571
rect 16037 9537 16071 9571
rect 17785 9537 17819 9571
rect 19901 9537 19935 9571
rect 20361 9537 20395 9571
rect 23765 9537 23799 9571
rect 24409 9537 24443 9571
rect 3893 9469 3927 9503
rect 6653 9469 6687 9503
rect 7113 9469 7147 9503
rect 7389 9469 7423 9503
rect 8744 9469 8778 9503
rect 10793 9469 10827 9503
rect 11320 9469 11354 9503
rect 14289 9469 14323 9503
rect 14473 9469 14507 9503
rect 15577 9469 15611 9503
rect 15853 9469 15887 9503
rect 16589 9469 16623 9503
rect 18245 9469 18279 9503
rect 18613 9469 18647 9503
rect 18981 9469 19015 9503
rect 19349 9469 19383 9503
rect 20453 9469 20487 9503
rect 22477 9469 22511 9503
rect 25237 9469 25271 9503
rect 25789 9469 25823 9503
rect 1685 9401 1719 9435
rect 2053 9401 2087 9435
rect 2507 9401 2541 9435
rect 5365 9401 5399 9435
rect 9781 9401 9815 9435
rect 9873 9401 9907 9435
rect 11161 9401 11195 9435
rect 12633 9401 12667 9435
rect 17049 9401 17083 9435
rect 17417 9401 17451 9435
rect 20815 9401 20849 9435
rect 22385 9401 22419 9435
rect 23857 9401 23891 9435
rect 4077 9333 4111 9367
rect 5089 9333 5123 9367
rect 6193 9333 6227 9367
rect 6929 9333 6963 9367
rect 7849 9333 7883 9367
rect 8815 9333 8849 9367
rect 9505 9333 9539 9367
rect 12081 9333 12115 9367
rect 14105 9333 14139 9367
rect 22661 9333 22695 9367
rect 25421 9333 25455 9367
rect 1869 9129 1903 9163
rect 2605 9129 2639 9163
rect 4261 9129 4295 9163
rect 5825 9129 5859 9163
rect 6193 9129 6227 9163
rect 7297 9129 7331 9163
rect 9505 9129 9539 9163
rect 11897 9129 11931 9163
rect 14381 9129 14415 9163
rect 15761 9129 15795 9163
rect 19809 9129 19843 9163
rect 20177 9129 20211 9163
rect 21373 9129 21407 9163
rect 23305 9129 23339 9163
rect 23765 9129 23799 9163
rect 25053 9129 25087 9163
rect 5226 9061 5260 9095
rect 6837 9061 6871 9095
rect 8211 9061 8245 9095
rect 10010 9061 10044 9095
rect 12310 9061 12344 9095
rect 13185 9061 13219 9095
rect 14749 9061 14783 9095
rect 21786 9061 21820 9095
rect 24133 9061 24167 9095
rect 24225 9061 24259 9095
rect 1869 8993 1903 9027
rect 2053 8993 2087 9027
rect 11989 8993 12023 9027
rect 14197 8993 14231 9027
rect 15117 8993 15151 9027
rect 15945 8993 15979 9027
rect 16405 8993 16439 9027
rect 16589 8993 16623 9027
rect 16865 8993 16899 9027
rect 18245 8993 18279 9027
rect 18797 8993 18831 9027
rect 18981 8993 19015 9027
rect 19349 8993 19383 9027
rect 22385 8993 22419 9027
rect 4905 8925 4939 8959
rect 7757 8925 7791 8959
rect 7849 8925 7883 8959
rect 9689 8925 9723 8959
rect 14105 8925 14139 8959
rect 17969 8925 18003 8959
rect 19533 8925 19567 8959
rect 21465 8925 21499 8959
rect 24409 8925 24443 8959
rect 8769 8789 8803 8823
rect 10609 8789 10643 8823
rect 12909 8789 12943 8823
rect 15577 8789 15611 8823
rect 17601 8789 17635 8823
rect 3893 8585 3927 8619
rect 3985 8585 4019 8619
rect 5549 8585 5583 8619
rect 6561 8585 6595 8619
rect 7021 8585 7055 8619
rect 9321 8585 9355 8619
rect 9597 8585 9631 8619
rect 10701 8585 10735 8619
rect 13645 8585 13679 8619
rect 20637 8585 20671 8619
rect 23489 8585 23523 8619
rect 25513 8585 25547 8619
rect 3709 8449 3743 8483
rect 1869 8381 1903 8415
rect 2237 8381 2271 8415
rect 2421 8381 2455 8415
rect 2973 8381 3007 8415
rect 5917 8517 5951 8551
rect 14197 8517 14231 8551
rect 17509 8517 17543 8551
rect 19901 8517 19935 8551
rect 25237 8517 25271 8551
rect 4261 8449 4295 8483
rect 4905 8449 4939 8483
rect 9781 8449 9815 8483
rect 10977 8449 11011 8483
rect 11529 8449 11563 8483
rect 11989 8449 12023 8483
rect 12541 8449 12575 8483
rect 13001 8449 13035 8483
rect 14565 8449 14599 8483
rect 19625 8449 19659 8483
rect 21465 8449 21499 8483
rect 22661 8449 22695 8483
rect 24501 8449 24535 8483
rect 5733 8381 5767 8415
rect 6837 8381 6871 8415
rect 8033 8381 8067 8415
rect 8953 8381 8987 8415
rect 11621 8381 11655 8415
rect 14105 8381 14139 8415
rect 14381 8381 14415 8415
rect 15117 8381 15151 8415
rect 15945 8381 15979 8415
rect 16405 8381 16439 8415
rect 16589 8381 16623 8415
rect 16957 8381 16991 8415
rect 18245 8381 18279 8415
rect 18797 8381 18831 8415
rect 18981 8381 19015 8415
rect 19533 8381 19567 8415
rect 20453 8381 20487 8415
rect 22385 8381 22419 8415
rect 3893 8313 3927 8347
rect 4353 8313 4387 8347
rect 6285 8313 6319 8347
rect 8355 8313 8389 8347
rect 10102 8313 10136 8347
rect 11529 8313 11563 8347
rect 12633 8313 12667 8347
rect 14013 8313 14047 8347
rect 15577 8313 15611 8347
rect 17785 8313 17819 8347
rect 20269 8313 20303 8347
rect 21786 8313 21820 8347
rect 24225 8313 24259 8347
rect 24317 8313 24351 8347
rect 2237 8245 2271 8279
rect 5181 8245 5215 8279
rect 7481 8245 7515 8279
rect 7849 8245 7883 8279
rect 15945 8245 15979 8279
rect 20913 8245 20947 8279
rect 21281 8245 21315 8279
rect 24041 8245 24075 8279
rect 1685 8041 1719 8075
rect 4169 8041 4203 8075
rect 5733 8041 5767 8075
rect 7297 8041 7331 8075
rect 9505 8041 9539 8075
rect 11989 8041 12023 8075
rect 12449 8041 12483 8075
rect 14013 8041 14047 8075
rect 16405 8041 16439 8075
rect 17049 8041 17083 8075
rect 19441 8041 19475 8075
rect 21925 8041 21959 8075
rect 2558 7973 2592 8007
rect 9781 7973 9815 8007
rect 9873 7973 9907 8007
rect 12817 7973 12851 8007
rect 14749 7973 14783 8007
rect 15117 7973 15151 8007
rect 16681 7973 16715 8007
rect 21097 7973 21131 8007
rect 22661 7973 22695 8007
rect 24041 7973 24075 8007
rect 2237 7905 2271 7939
rect 4169 7905 4203 7939
rect 4537 7905 4571 7939
rect 5917 7905 5951 7939
rect 6193 7905 6227 7939
rect 7481 7905 7515 7939
rect 7665 7905 7699 7939
rect 8401 7905 8435 7939
rect 11437 7905 11471 7939
rect 14197 7905 14231 7939
rect 15301 7905 15335 7939
rect 15577 7905 15611 7939
rect 16865 7905 16899 7939
rect 17417 7905 17451 7939
rect 18245 7905 18279 7939
rect 18705 7905 18739 7939
rect 19073 7905 19107 7939
rect 19533 7905 19567 7939
rect 24133 7905 24167 7939
rect 2053 7837 2087 7871
rect 10149 7837 10183 7871
rect 10701 7837 10735 7871
rect 12725 7837 12759 7871
rect 13369 7837 13403 7871
rect 15761 7837 15795 7871
rect 21005 7837 21039 7871
rect 22569 7837 22603 7871
rect 6837 7769 6871 7803
rect 11621 7769 11655 7803
rect 15393 7769 15427 7803
rect 18061 7769 18095 7803
rect 21557 7769 21591 7803
rect 23121 7769 23155 7803
rect 3157 7701 3191 7735
rect 8861 7701 8895 7735
rect 13737 7701 13771 7735
rect 14381 7701 14415 7735
rect 17785 7701 17819 7735
rect 20177 7701 20211 7735
rect 1593 7497 1627 7531
rect 4721 7497 4755 7531
rect 6193 7497 6227 7531
rect 7941 7497 7975 7531
rect 8309 7497 8343 7531
rect 9781 7497 9815 7531
rect 11437 7497 11471 7531
rect 13553 7497 13587 7531
rect 15853 7497 15887 7531
rect 16129 7497 16163 7531
rect 18337 7497 18371 7531
rect 24685 7497 24719 7531
rect 2053 7429 2087 7463
rect 6561 7429 6595 7463
rect 10885 7429 10919 7463
rect 12541 7429 12575 7463
rect 14105 7429 14139 7463
rect 21097 7429 21131 7463
rect 3617 7361 3651 7395
rect 4905 7361 4939 7395
rect 10333 7361 10367 7395
rect 14657 7361 14691 7395
rect 15485 7361 15519 7395
rect 19349 7361 19383 7395
rect 21741 7361 21775 7395
rect 22293 7361 22327 7395
rect 23765 7361 23799 7395
rect 24041 7361 24075 7395
rect 1409 7293 1443 7327
rect 6837 7293 6871 7327
rect 7297 7293 7331 7327
rect 8401 7293 8435 7327
rect 8861 7293 8895 7327
rect 12449 7293 12483 7327
rect 12725 7293 12759 7327
rect 14013 7293 14047 7327
rect 14289 7293 14323 7327
rect 16589 7293 16623 7327
rect 19165 7293 19199 7327
rect 20177 7293 20211 7327
rect 25237 7293 25271 7327
rect 25789 7293 25823 7327
rect 2973 7225 3007 7259
rect 3065 7225 3099 7259
rect 5226 7225 5260 7259
rect 10149 7225 10183 7259
rect 10425 7225 10459 7259
rect 11897 7225 11931 7259
rect 17141 7225 17175 7259
rect 20498 7225 20532 7259
rect 21373 7225 21407 7259
rect 22017 7225 22051 7259
rect 22109 7225 22143 7259
rect 23489 7225 23523 7259
rect 23857 7225 23891 7259
rect 2329 7157 2363 7191
rect 2789 7157 2823 7191
rect 4169 7157 4203 7191
rect 5825 7157 5859 7191
rect 6929 7157 6963 7191
rect 8493 7157 8527 7191
rect 12265 7157 12299 7191
rect 12909 7157 12943 7191
rect 13829 7157 13863 7191
rect 15117 7157 15151 7191
rect 17417 7157 17451 7191
rect 17877 7157 17911 7191
rect 19625 7157 19659 7191
rect 20085 7157 20119 7191
rect 22937 7157 22971 7191
rect 25421 7157 25455 7191
rect 2053 6953 2087 6987
rect 3893 6953 3927 6987
rect 5089 6953 5123 6987
rect 5641 6953 5675 6987
rect 6929 6953 6963 6987
rect 7297 6953 7331 6987
rect 9781 6953 9815 6987
rect 13185 6953 13219 6987
rect 14013 6953 14047 6987
rect 16957 6953 16991 6987
rect 17417 6953 17451 6987
rect 20729 6953 20763 6987
rect 21649 6953 21683 6987
rect 22017 6953 22051 6987
rect 23305 6953 23339 6987
rect 23765 6953 23799 6987
rect 2329 6885 2363 6919
rect 4261 6885 4295 6919
rect 6054 6885 6088 6919
rect 7665 6885 7699 6919
rect 13737 6885 13771 6919
rect 22471 6885 22505 6919
rect 24133 6885 24167 6919
rect 5733 6817 5767 6851
rect 6653 6817 6687 6851
rect 9505 6817 9539 6851
rect 9965 6817 9999 6851
rect 10149 6817 10183 6851
rect 12173 6817 12207 6851
rect 12449 6817 12483 6851
rect 14197 6817 14231 6851
rect 14657 6817 14691 6851
rect 15853 6817 15887 6851
rect 16037 6817 16071 6851
rect 16589 6817 16623 6851
rect 16865 6817 16899 6851
rect 18153 6817 18187 6851
rect 18613 6817 18647 6851
rect 18705 6817 18739 6851
rect 19073 6817 19107 6851
rect 19993 6817 20027 6851
rect 21005 6817 21039 6851
rect 22109 6817 22143 6851
rect 2237 6749 2271 6783
rect 2881 6749 2915 6783
rect 3157 6749 3191 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 7573 6749 7607 6783
rect 7849 6749 7883 6783
rect 11713 6749 11747 6783
rect 12633 6749 12667 6783
rect 15117 6749 15151 6783
rect 24041 6749 24075 6783
rect 24685 6749 24719 6783
rect 12265 6681 12299 6715
rect 14381 6681 14415 6715
rect 19257 6681 19291 6715
rect 1593 6613 1627 6647
rect 8769 6613 8803 6647
rect 10885 6613 10919 6647
rect 12081 6613 12115 6647
rect 17693 6613 17727 6647
rect 19625 6613 19659 6647
rect 21189 6613 21223 6647
rect 23029 6613 23063 6647
rect 4261 6409 4295 6443
rect 4721 6409 4755 6443
rect 7849 6409 7883 6443
rect 10057 6409 10091 6443
rect 13461 6409 13495 6443
rect 13921 6409 13955 6443
rect 17509 6409 17543 6443
rect 17785 6409 17819 6443
rect 21281 6409 21315 6443
rect 21741 6409 21775 6443
rect 22661 6409 22695 6443
rect 23489 6409 23523 6443
rect 25329 6409 25363 6443
rect 3617 6341 3651 6375
rect 6193 6341 6227 6375
rect 10885 6341 10919 6375
rect 16681 6341 16715 6375
rect 5733 6273 5767 6307
rect 11253 6273 11287 6307
rect 11897 6273 11931 6307
rect 16313 6273 16347 6307
rect 19809 6273 19843 6307
rect 24409 6273 24443 6307
rect 2329 6205 2363 6239
rect 3249 6205 3283 6239
rect 4077 6205 4111 6239
rect 6837 6205 6871 6239
rect 7297 6205 7331 6239
rect 8769 6205 8803 6239
rect 10793 6205 10827 6239
rect 11069 6205 11103 6239
rect 12449 6205 12483 6239
rect 12541 6205 12575 6239
rect 12725 6205 12759 6239
rect 14013 6205 14047 6239
rect 14565 6205 14599 6239
rect 15577 6205 15611 6239
rect 15669 6205 15703 6239
rect 15853 6205 15887 6239
rect 18245 6205 18279 6239
rect 18521 6205 18555 6239
rect 18889 6205 18923 6239
rect 19349 6205 19383 6239
rect 20361 6205 20395 6239
rect 22477 6205 22511 6239
rect 23029 6205 23063 6239
rect 2145 6137 2179 6171
rect 2650 6137 2684 6171
rect 5273 6137 5307 6171
rect 5365 6137 5399 6171
rect 9131 6137 9165 6171
rect 10701 6137 10735 6171
rect 15117 6137 15151 6171
rect 20723 6137 20757 6171
rect 24501 6137 24535 6171
rect 25053 6137 25087 6171
rect 1869 6069 1903 6103
rect 3985 6069 4019 6103
rect 5089 6069 5123 6103
rect 6561 6069 6595 6103
rect 6929 6069 6963 6103
rect 8217 6069 8251 6103
rect 8677 6069 8711 6103
rect 9689 6069 9723 6103
rect 12265 6069 12299 6103
rect 12909 6069 12943 6103
rect 14105 6069 14139 6103
rect 15485 6069 15519 6103
rect 17049 6069 17083 6103
rect 19257 6069 19291 6103
rect 20269 6069 20303 6103
rect 22201 6069 22235 6103
rect 24133 6069 24167 6103
rect 1869 5865 1903 5899
rect 2881 5865 2915 5899
rect 5825 5865 5859 5899
rect 7297 5865 7331 5899
rect 9413 5865 9447 5899
rect 10885 5865 10919 5899
rect 11529 5865 11563 5899
rect 12817 5865 12851 5899
rect 13553 5865 13587 5899
rect 14657 5865 14691 5899
rect 17141 5865 17175 5899
rect 17601 5865 17635 5899
rect 19441 5865 19475 5899
rect 19809 5865 19843 5899
rect 23121 5865 23155 5899
rect 2282 5797 2316 5831
rect 3525 5797 3559 5831
rect 4261 5797 4295 5831
rect 6330 5797 6364 5831
rect 8217 5797 8251 5831
rect 9873 5797 9907 5831
rect 19165 5797 19199 5831
rect 20361 5797 20395 5831
rect 22522 5797 22556 5831
rect 24409 5797 24443 5831
rect 24961 5797 24995 5831
rect 3801 5729 3835 5763
rect 6009 5729 6043 5763
rect 11897 5729 11931 5763
rect 13829 5729 13863 5763
rect 15577 5729 15611 5763
rect 15853 5729 15887 5763
rect 16405 5729 16439 5763
rect 16773 5729 16807 5763
rect 17693 5729 17727 5763
rect 18153 5729 18187 5763
rect 18613 5729 18647 5763
rect 18981 5729 19015 5763
rect 20913 5729 20947 5763
rect 21833 5729 21867 5763
rect 22201 5729 22235 5763
rect 1961 5661 1995 5695
rect 4169 5661 4203 5695
rect 4813 5661 4847 5695
rect 5181 5661 5215 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 9781 5661 9815 5695
rect 10057 5661 10091 5695
rect 14381 5661 14415 5695
rect 15025 5661 15059 5695
rect 16865 5661 16899 5695
rect 24317 5661 24351 5695
rect 8677 5593 8711 5627
rect 12541 5593 12575 5627
rect 21465 5593 21499 5627
rect 6929 5525 6963 5559
rect 9137 5525 9171 5559
rect 21097 5525 21131 5559
rect 24041 5525 24075 5559
rect 1593 5321 1627 5355
rect 2053 5321 2087 5355
rect 3709 5321 3743 5355
rect 5733 5321 5767 5355
rect 7941 5321 7975 5355
rect 9781 5321 9815 5355
rect 13645 5321 13679 5355
rect 19073 5321 19107 5355
rect 19441 5321 19475 5355
rect 22753 5321 22787 5355
rect 7481 5253 7515 5287
rect 11897 5253 11931 5287
rect 15669 5253 15703 5287
rect 17785 5253 17819 5287
rect 24961 5253 24995 5287
rect 2973 5185 3007 5219
rect 4445 5185 4479 5219
rect 4813 5185 4847 5219
rect 6009 5185 6043 5219
rect 6929 5185 6963 5219
rect 9137 5185 9171 5219
rect 10057 5185 10091 5219
rect 10701 5185 10735 5219
rect 12449 5185 12483 5219
rect 16865 5185 16899 5219
rect 18153 5185 18187 5219
rect 18521 5185 18555 5219
rect 21189 5185 21223 5219
rect 25329 5185 25363 5219
rect 1409 5117 1443 5151
rect 12265 5117 12299 5151
rect 13001 5117 13035 5151
rect 14289 5117 14323 5151
rect 14381 5117 14415 5151
rect 14565 5117 14599 5151
rect 15853 5117 15887 5151
rect 15945 5117 15979 5151
rect 16129 5117 16163 5151
rect 18061 5117 18095 5151
rect 18337 5117 18371 5151
rect 20269 5117 20303 5151
rect 20729 5117 20763 5151
rect 2697 5049 2731 5083
rect 2789 5049 2823 5083
rect 4537 5049 4571 5083
rect 6561 5049 6595 5083
rect 7021 5049 7055 5083
rect 8493 5049 8527 5083
rect 8585 5049 8619 5083
rect 10149 5049 10183 5083
rect 14105 5049 14139 5083
rect 15301 5049 15335 5083
rect 20361 5049 20395 5083
rect 21510 5049 21544 5083
rect 22385 5049 22419 5083
rect 23489 5049 23523 5083
rect 24409 5049 24443 5083
rect 24501 5049 24535 5083
rect 2513 4981 2547 5015
rect 4261 4981 4295 5015
rect 8309 4981 8343 5015
rect 11345 4981 11379 5015
rect 14749 4981 14783 5015
rect 16313 4981 16347 5015
rect 17509 4981 17543 5015
rect 21005 4981 21039 5015
rect 22109 4981 22143 5015
rect 24225 4981 24259 5015
rect 1593 4777 1627 4811
rect 1961 4777 1995 4811
rect 3249 4777 3283 4811
rect 3801 4777 3835 4811
rect 5089 4777 5123 4811
rect 6239 4777 6273 4811
rect 8401 4777 8435 4811
rect 9965 4777 9999 4811
rect 10425 4777 10459 4811
rect 13277 4777 13311 4811
rect 15393 4777 15427 4811
rect 17049 4777 17083 4811
rect 17509 4777 17543 4811
rect 20269 4777 20303 4811
rect 20729 4777 20763 4811
rect 23489 4777 23523 4811
rect 24317 4777 24351 4811
rect 25053 4777 25087 4811
rect 2237 4709 2271 4743
rect 2329 4709 2363 4743
rect 2881 4709 2915 4743
rect 4261 4709 4295 4743
rect 4813 4709 4847 4743
rect 7021 4709 7055 4743
rect 7205 4709 7239 4743
rect 7297 4709 7331 4743
rect 10701 4709 10735 4743
rect 10793 4709 10827 4743
rect 15117 4709 15151 4743
rect 19026 4709 19060 4743
rect 21097 4709 21131 4743
rect 22661 4709 22695 4743
rect 6136 4641 6170 4675
rect 12817 4641 12851 4675
rect 14105 4641 14139 4675
rect 15577 4641 15611 4675
rect 15945 4641 15979 4675
rect 16313 4641 16347 4675
rect 16589 4641 16623 4675
rect 17601 4641 17635 4675
rect 18153 4641 18187 4675
rect 24133 4641 24167 4675
rect 4169 4573 4203 4607
rect 7481 4573 7515 4607
rect 11345 4573 11379 4607
rect 11621 4573 11655 4607
rect 14657 4573 14691 4607
rect 18705 4573 18739 4607
rect 21005 4573 21039 4607
rect 21281 4573 21315 4607
rect 22293 4573 22327 4607
rect 22569 4573 22603 4607
rect 9413 4505 9447 4539
rect 14289 4505 14323 4539
rect 19625 4505 19659 4539
rect 19993 4505 20027 4539
rect 21925 4505 21959 4539
rect 23121 4505 23155 4539
rect 9137 4437 9171 4471
rect 11989 4437 12023 4471
rect 12633 4437 12667 4471
rect 13645 4437 13679 4471
rect 14013 4437 14047 4471
rect 17785 4437 17819 4471
rect 18521 4437 18555 4471
rect 4169 4233 4203 4267
rect 4445 4233 4479 4267
rect 6193 4233 6227 4267
rect 13461 4233 13495 4267
rect 13921 4233 13955 4267
rect 17877 4233 17911 4267
rect 21373 4233 21407 4267
rect 23029 4233 23063 4267
rect 23397 4233 23431 4267
rect 24685 4233 24719 4267
rect 16865 4165 16899 4199
rect 1961 4097 1995 4131
rect 2789 4097 2823 4131
rect 3065 4097 3099 4131
rect 3709 4097 3743 4131
rect 6561 4097 6595 4131
rect 7573 4097 7607 4131
rect 7849 4097 7883 4131
rect 9137 4097 9171 4131
rect 9781 4097 9815 4131
rect 12541 4097 12575 4131
rect 14289 4097 14323 4131
rect 17509 4097 17543 4131
rect 20453 4097 20487 4131
rect 21097 4097 21131 4131
rect 22109 4097 22143 4131
rect 22385 4097 22419 4131
rect 25789 4097 25823 4131
rect 1409 4029 1443 4063
rect 1869 4029 1903 4063
rect 2421 4029 2455 4063
rect 5089 4029 5123 4063
rect 5825 4029 5859 4063
rect 10149 4029 10183 4063
rect 10609 4029 10643 4063
rect 11897 4029 11931 4063
rect 14657 4029 14691 4063
rect 15025 4029 15059 4063
rect 15393 4029 15427 4063
rect 15853 4029 15887 4063
rect 16129 4029 16163 4063
rect 16497 4029 16531 4063
rect 18061 4029 18095 4063
rect 18521 4029 18555 4063
rect 18889 4029 18923 4063
rect 19349 4029 19383 4063
rect 23765 4029 23799 4063
rect 25237 4029 25271 4063
rect 3157 3961 3191 3995
rect 7297 3961 7331 3995
rect 7665 3961 7699 3995
rect 8493 3961 8527 3995
rect 8953 3961 8987 3995
rect 9229 3961 9263 3995
rect 10517 3961 10551 3995
rect 10971 3961 11005 3995
rect 12265 3961 12299 3995
rect 12903 3961 12937 3995
rect 19533 3961 19567 3995
rect 20545 3961 20579 3995
rect 22201 3961 22235 3995
rect 23673 3961 23707 3995
rect 5457 3893 5491 3927
rect 11529 3893 11563 3927
rect 15209 3893 15243 3927
rect 19901 3893 19935 3927
rect 20177 3893 20211 3927
rect 21925 3893 21959 3927
rect 25421 3893 25455 3927
rect 1593 3689 1627 3723
rect 2237 3689 2271 3723
rect 2697 3689 2731 3723
rect 3157 3689 3191 3723
rect 3433 3689 3467 3723
rect 9827 3689 9861 3723
rect 10333 3689 10367 3723
rect 12081 3689 12115 3723
rect 15117 3689 15151 3723
rect 15393 3689 15427 3723
rect 17141 3689 17175 3723
rect 17509 3689 17543 3723
rect 19809 3689 19843 3723
rect 20453 3689 20487 3723
rect 22109 3689 22143 3723
rect 23489 3689 23523 3723
rect 6009 3621 6043 3655
rect 6561 3621 6595 3655
rect 7751 3621 7785 3655
rect 11161 3621 11195 3655
rect 11713 3621 11747 3655
rect 12725 3621 12759 3655
rect 14749 3621 14783 3655
rect 21097 3621 21131 3655
rect 22569 3621 22603 3655
rect 22661 3621 22695 3655
rect 24041 3621 24075 3655
rect 1409 3553 1443 3587
rect 2973 3553 3007 3587
rect 4261 3553 4295 3587
rect 4537 3553 4571 3587
rect 4997 3553 5031 3587
rect 7389 3553 7423 3587
rect 9724 3553 9758 3587
rect 14105 3553 14139 3587
rect 15301 3553 15335 3587
rect 15945 3553 15979 3587
rect 16221 3553 16255 3587
rect 16681 3553 16715 3587
rect 17693 3553 17727 3587
rect 18337 3553 18371 3587
rect 18521 3553 18555 3587
rect 18889 3553 18923 3587
rect 24685 3553 24719 3587
rect 5917 3485 5951 3519
rect 9229 3485 9263 3519
rect 11069 3485 11103 3519
rect 12633 3485 12667 3519
rect 13093 3485 13127 3519
rect 13645 3485 13679 3519
rect 19165 3485 19199 3519
rect 21005 3485 21039 3519
rect 21281 3485 21315 3519
rect 23029 3485 23063 3519
rect 4353 3417 4387 3451
rect 14289 3417 14323 3451
rect 19441 3417 19475 3451
rect 5365 3349 5399 3383
rect 7113 3349 7147 3383
rect 8309 3349 8343 3383
rect 8861 3349 8895 3383
rect 10701 3349 10735 3383
rect 12449 3349 12483 3383
rect 14013 3349 14047 3383
rect 1593 3145 1627 3179
rect 2053 3145 2087 3179
rect 2329 3145 2363 3179
rect 3157 3145 3191 3179
rect 4629 3145 4663 3179
rect 6561 3145 6595 3179
rect 8217 3145 8251 3179
rect 8677 3145 8711 3179
rect 9781 3145 9815 3179
rect 10057 3145 10091 3179
rect 10517 3145 10551 3179
rect 12265 3145 12299 3179
rect 13461 3145 13495 3179
rect 15393 3145 15427 3179
rect 17693 3145 17727 3179
rect 19809 3145 19843 3179
rect 21649 3145 21683 3179
rect 24685 3145 24719 3179
rect 25421 3145 25455 3179
rect 2789 3077 2823 3111
rect 5089 3077 5123 3111
rect 7849 3077 7883 3111
rect 13093 3077 13127 3111
rect 13829 3077 13863 3111
rect 14105 3077 14139 3111
rect 23489 3077 23523 3111
rect 4353 3009 4387 3043
rect 5917 3009 5951 3043
rect 6193 3009 6227 3043
rect 7297 3009 7331 3043
rect 8861 3009 8895 3043
rect 10701 3009 10735 3043
rect 11345 3009 11379 3043
rect 12541 3009 12575 3043
rect 14749 3009 14783 3043
rect 17417 3009 17451 3043
rect 20453 3009 20487 3043
rect 22109 3009 22143 3043
rect 24041 3009 24075 3043
rect 1409 2941 1443 2975
rect 2605 2941 2639 2975
rect 3525 2941 3559 2975
rect 4077 2941 4111 2975
rect 5365 2941 5399 2975
rect 7021 2941 7055 2975
rect 14013 2941 14047 2975
rect 14289 2941 14323 2975
rect 15761 2941 15795 2975
rect 16037 2941 16071 2975
rect 16405 2941 16439 2975
rect 16773 2941 16807 2975
rect 18061 2941 18095 2975
rect 18521 2941 18555 2975
rect 18889 2941 18923 2975
rect 19257 2941 19291 2975
rect 22477 2941 22511 2975
rect 25237 2941 25271 2975
rect 25789 2941 25823 2975
rect 7389 2873 7423 2907
rect 9182 2873 9216 2907
rect 10793 2873 10827 2907
rect 12633 2873 12667 2907
rect 20774 2873 20808 2907
rect 23765 2873 23799 2907
rect 23857 2873 23891 2907
rect 11713 2805 11747 2839
rect 16773 2805 16807 2839
rect 19257 2805 19291 2839
rect 20269 2805 20303 2839
rect 21373 2805 21407 2839
rect 22661 2805 22695 2839
rect 23121 2805 23155 2839
rect 2513 2601 2547 2635
rect 5181 2601 5215 2635
rect 6377 2601 6411 2635
rect 6745 2601 6779 2635
rect 7251 2601 7285 2635
rect 9505 2601 9539 2635
rect 10425 2601 10459 2635
rect 12449 2601 12483 2635
rect 13645 2601 13679 2635
rect 14105 2601 14139 2635
rect 14933 2601 14967 2635
rect 15301 2601 15335 2635
rect 16589 2601 16623 2635
rect 17785 2601 17819 2635
rect 19625 2601 19659 2635
rect 21005 2601 21039 2635
rect 22569 2601 22603 2635
rect 23765 2601 23799 2635
rect 25421 2601 25455 2635
rect 2053 2533 2087 2567
rect 8217 2533 8251 2567
rect 8309 2533 8343 2567
rect 10793 2533 10827 2567
rect 11069 2533 11103 2567
rect 11621 2533 11655 2567
rect 12633 2533 12667 2567
rect 18153 2533 18187 2567
rect 18791 2533 18825 2567
rect 21373 2533 21407 2567
rect 22201 2533 22235 2567
rect 24041 2533 24075 2567
rect 1409 2465 1443 2499
rect 4261 2465 4295 2499
rect 4813 2465 4847 2499
rect 5917 2465 5951 2499
rect 7021 2465 7055 2499
rect 7148 2465 7182 2499
rect 8861 2465 8895 2499
rect 9873 2465 9907 2499
rect 12725 2465 12759 2499
rect 14289 2465 14323 2499
rect 15577 2465 15611 2499
rect 17325 2465 17359 2499
rect 19349 2465 19383 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 24133 2465 24167 2499
rect 25053 2465 25087 2499
rect 25672 2465 25706 2499
rect 6009 2397 6043 2431
rect 7941 2397 7975 2431
rect 9229 2397 9263 2431
rect 10977 2397 11011 2431
rect 11897 2397 11931 2431
rect 16129 2397 16163 2431
rect 17417 2397 17451 2431
rect 18429 2397 18463 2431
rect 21281 2397 21315 2431
rect 21557 2397 21591 2431
rect 7021 2329 7055 2363
rect 7573 2329 7607 2363
rect 25743 2329 25777 2363
rect 1593 2261 1627 2295
rect 4445 2261 4479 2295
rect 10057 2261 10091 2295
rect 14473 2261 14507 2295
rect 15761 2261 15795 2295
rect 23029 2261 23063 2295
rect 26157 2261 26191 2295
rect 26433 2261 26467 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 24762 23808 24768 23860
rect 24820 23848 24826 23860
rect 25041 23851 25099 23857
rect 25041 23848 25053 23851
rect 24820 23820 25053 23848
rect 24820 23808 24826 23820
rect 25041 23817 25053 23820
rect 25087 23817 25099 23851
rect 25041 23811 25099 23817
rect 13538 23712 13544 23724
rect 13499 23684 13544 23712
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 1394 23604 1400 23656
rect 1452 23653 1458 23656
rect 1452 23647 1490 23653
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1452 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 13056 23647 13114 23653
rect 13056 23613 13068 23647
rect 13102 23644 13114 23647
rect 13556 23644 13584 23672
rect 13102 23616 13584 23644
rect 24648 23647 24706 23653
rect 13102 23613 13114 23616
rect 13056 23607 13114 23613
rect 24648 23613 24660 23647
rect 24694 23644 24706 23647
rect 24762 23644 24768 23656
rect 24694 23616 24768 23644
rect 24694 23613 24706 23616
rect 24648 23607 24706 23613
rect 1452 23604 1458 23607
rect 24762 23604 24768 23616
rect 24820 23604 24826 23656
rect 1535 23511 1593 23517
rect 1535 23477 1547 23511
rect 1581 23508 1593 23511
rect 1762 23508 1768 23520
rect 1581 23480 1768 23508
rect 1581 23477 1593 23480
rect 1535 23471 1593 23477
rect 1762 23468 1768 23480
rect 1820 23468 1826 23520
rect 13127 23511 13185 23517
rect 13127 23477 13139 23511
rect 13173 23508 13185 23511
rect 13354 23508 13360 23520
rect 13173 23480 13360 23508
rect 13173 23477 13185 23480
rect 13127 23471 13185 23477
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 23474 23468 23480 23520
rect 23532 23508 23538 23520
rect 24719 23511 24777 23517
rect 24719 23508 24731 23511
rect 23532 23480 24731 23508
rect 23532 23468 23538 23480
rect 24719 23477 24731 23480
rect 24765 23477 24777 23511
rect 24719 23471 24777 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 24670 22720 24676 22772
rect 24728 22760 24734 22772
rect 25041 22763 25099 22769
rect 25041 22760 25053 22763
rect 24728 22732 25053 22760
rect 24728 22720 24734 22732
rect 25041 22729 25053 22732
rect 25087 22729 25099 22763
rect 25041 22723 25099 22729
rect 24670 22565 24676 22568
rect 24648 22559 24676 22565
rect 24648 22525 24660 22559
rect 24648 22519 24676 22525
rect 24670 22516 24676 22519
rect 24728 22516 24734 22568
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 24719 22423 24777 22429
rect 24719 22420 24731 22423
rect 23716 22392 24731 22420
rect 23716 22380 23722 22392
rect 24719 22389 24731 22392
rect 24765 22389 24777 22423
rect 24719 22383 24777 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 12964 21471 13022 21477
rect 12964 21437 12976 21471
rect 13010 21468 13022 21471
rect 13010 21440 13492 21468
rect 13010 21437 13022 21440
rect 12964 21431 13022 21437
rect 13464 21412 13492 21440
rect 13446 21400 13452 21412
rect 13407 21372 13452 21400
rect 13446 21360 13452 21372
rect 13504 21360 13510 21412
rect 13035 21335 13093 21341
rect 13035 21301 13047 21335
rect 13081 21332 13093 21335
rect 13538 21332 13544 21344
rect 13081 21304 13544 21332
rect 13081 21301 13093 21304
rect 13035 21295 13093 21301
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1464 20995 1522 21001
rect 1464 20961 1476 20995
rect 1510 20992 1522 20995
rect 1854 20992 1860 21004
rect 1510 20964 1860 20992
rect 1510 20961 1522 20964
rect 1464 20955 1522 20961
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 2476 20995 2534 21001
rect 2476 20961 2488 20995
rect 2522 20992 2534 20995
rect 2682 20992 2688 21004
rect 2522 20964 2688 20992
rect 2522 20961 2534 20964
rect 2476 20955 2534 20961
rect 2682 20952 2688 20964
rect 2740 20992 2746 21004
rect 2774 20992 2780 21004
rect 2740 20964 2780 20992
rect 2740 20952 2746 20964
rect 2774 20952 2780 20964
rect 2832 20952 2838 21004
rect 24670 21001 24676 21004
rect 24648 20995 24676 21001
rect 24648 20961 24660 20995
rect 24648 20955 24676 20961
rect 24670 20952 24676 20955
rect 24728 20952 24734 21004
rect 1535 20859 1593 20865
rect 1535 20825 1547 20859
rect 1581 20856 1593 20859
rect 2130 20856 2136 20868
rect 1581 20828 2136 20856
rect 1581 20825 1593 20828
rect 1535 20819 1593 20825
rect 2130 20816 2136 20828
rect 2188 20816 2194 20868
rect 2547 20791 2605 20797
rect 2547 20757 2559 20791
rect 2593 20788 2605 20791
rect 3418 20788 3424 20800
rect 2593 20760 3424 20788
rect 2593 20757 2605 20760
rect 2547 20751 2605 20757
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 24719 20791 24777 20797
rect 24719 20788 24731 20791
rect 23532 20760 24731 20788
rect 23532 20748 23538 20760
rect 24719 20757 24731 20760
rect 24765 20757 24777 20791
rect 24719 20751 24777 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 3237 20587 3295 20593
rect 3237 20584 3249 20587
rect 2832 20556 3249 20584
rect 2832 20544 2838 20556
rect 3237 20553 3249 20556
rect 3283 20553 3295 20587
rect 24670 20584 24676 20596
rect 24631 20556 24676 20584
rect 3237 20547 3295 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 1535 20519 1593 20525
rect 1535 20485 1547 20519
rect 1581 20516 1593 20519
rect 2038 20516 2044 20528
rect 1581 20488 2044 20516
rect 1581 20485 1593 20488
rect 1535 20479 1593 20485
rect 2038 20476 2044 20488
rect 2096 20476 2102 20528
rect 2491 20420 3004 20448
rect 1464 20383 1522 20389
rect 1464 20349 1476 20383
rect 1510 20380 1522 20383
rect 1578 20380 1584 20392
rect 1510 20352 1584 20380
rect 1510 20349 1522 20352
rect 1464 20343 1522 20349
rect 1578 20340 1584 20352
rect 1636 20380 1642 20392
rect 2491 20389 2519 20420
rect 2225 20383 2283 20389
rect 2225 20380 2237 20383
rect 1636 20352 2237 20380
rect 1636 20340 1642 20352
rect 2225 20349 2237 20352
rect 2271 20349 2283 20383
rect 2225 20343 2283 20349
rect 2476 20383 2534 20389
rect 2476 20349 2488 20383
rect 2522 20349 2534 20383
rect 2476 20343 2534 20349
rect 2976 20321 3004 20420
rect 2961 20315 3019 20321
rect 1596 20284 1992 20312
rect 1596 20256 1624 20284
rect 1578 20204 1584 20256
rect 1636 20204 1642 20256
rect 1854 20244 1860 20256
rect 1815 20216 1860 20244
rect 1854 20204 1860 20216
rect 1912 20204 1918 20256
rect 1964 20244 1992 20284
rect 2961 20281 2973 20315
rect 3007 20312 3019 20315
rect 3142 20312 3148 20324
rect 3007 20284 3148 20312
rect 3007 20281 3019 20284
rect 2961 20275 3019 20281
rect 3142 20272 3148 20284
rect 3200 20272 3206 20324
rect 2547 20247 2605 20253
rect 2547 20244 2559 20247
rect 1964 20216 2559 20244
rect 2547 20213 2559 20216
rect 2593 20213 2605 20247
rect 2547 20207 2605 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1394 19864 1400 19916
rect 1452 19913 1458 19916
rect 1452 19907 1490 19913
rect 1478 19873 1490 19907
rect 1452 19867 1490 19873
rect 4132 19907 4190 19913
rect 4132 19873 4144 19907
rect 4178 19904 4190 19907
rect 4338 19904 4344 19916
rect 4178 19876 4344 19904
rect 4178 19873 4190 19876
rect 4132 19867 4190 19873
rect 1452 19864 1458 19867
rect 4338 19864 4344 19876
rect 4396 19864 4402 19916
rect 2409 19839 2467 19845
rect 2409 19805 2421 19839
rect 2455 19836 2467 19839
rect 2498 19836 2504 19848
rect 2455 19808 2504 19836
rect 2455 19805 2467 19808
rect 2409 19799 2467 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 1535 19703 1593 19709
rect 1535 19669 1547 19703
rect 1581 19700 1593 19703
rect 2314 19700 2320 19712
rect 1581 19672 2320 19700
rect 1581 19669 1593 19672
rect 1535 19663 1593 19669
rect 2314 19660 2320 19672
rect 2372 19660 2378 19712
rect 4203 19703 4261 19709
rect 4203 19669 4215 19703
rect 4249 19700 4261 19703
rect 4982 19700 4988 19712
rect 4249 19672 4988 19700
rect 4249 19669 4261 19672
rect 4203 19663 4261 19669
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1394 19456 1400 19508
rect 1452 19496 1458 19508
rect 2225 19499 2283 19505
rect 2225 19496 2237 19499
rect 1452 19468 2237 19496
rect 1452 19456 1458 19468
rect 2225 19465 2237 19468
rect 2271 19465 2283 19499
rect 2225 19459 2283 19465
rect 1394 19252 1400 19304
rect 1452 19301 1458 19304
rect 1452 19295 1490 19301
rect 1478 19292 1490 19295
rect 1857 19295 1915 19301
rect 1857 19292 1869 19295
rect 1478 19264 1869 19292
rect 1478 19261 1490 19264
rect 1452 19255 1490 19261
rect 1857 19261 1869 19264
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 2476 19295 2534 19301
rect 2476 19261 2488 19295
rect 2522 19292 2534 19295
rect 2958 19292 2964 19304
rect 2522 19264 2964 19292
rect 2522 19261 2534 19264
rect 2476 19255 2534 19261
rect 1452 19252 1458 19255
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 3488 19295 3546 19301
rect 3488 19261 3500 19295
rect 3534 19292 3546 19295
rect 3602 19292 3608 19304
rect 3534 19264 3608 19292
rect 3534 19261 3546 19264
rect 3488 19255 3546 19261
rect 3602 19252 3608 19264
rect 3660 19292 3666 19304
rect 3881 19295 3939 19301
rect 3881 19292 3893 19295
rect 3660 19264 3893 19292
rect 3660 19252 3666 19264
rect 3881 19261 3893 19264
rect 3927 19261 3939 19295
rect 3881 19255 3939 19261
rect 4500 19295 4558 19301
rect 4500 19261 4512 19295
rect 4546 19292 4558 19295
rect 5074 19292 5080 19304
rect 4546 19264 5080 19292
rect 4546 19261 4558 19264
rect 4500 19255 4558 19261
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 1535 19227 1593 19233
rect 1535 19193 1547 19227
rect 1581 19224 1593 19227
rect 2130 19224 2136 19236
rect 1581 19196 2136 19224
rect 1581 19193 1593 19196
rect 1535 19187 1593 19193
rect 2130 19184 2136 19196
rect 2188 19184 2194 19236
rect 2406 19116 2412 19168
rect 2464 19156 2470 19168
rect 2547 19159 2605 19165
rect 2547 19156 2559 19159
rect 2464 19128 2559 19156
rect 2464 19116 2470 19128
rect 2547 19125 2559 19128
rect 2593 19125 2605 19159
rect 2547 19119 2605 19125
rect 3142 19116 3148 19168
rect 3200 19156 3206 19168
rect 3559 19159 3617 19165
rect 3559 19156 3571 19159
rect 3200 19128 3571 19156
rect 3200 19116 3206 19128
rect 3559 19125 3571 19128
rect 3605 19125 3617 19159
rect 4338 19156 4344 19168
rect 4299 19128 4344 19156
rect 3559 19119 3617 19125
rect 4338 19116 4344 19128
rect 4396 19116 4402 19168
rect 4522 19116 4528 19168
rect 4580 19165 4586 19168
rect 4580 19159 4629 19165
rect 4580 19125 4583 19159
rect 4617 19125 4629 19159
rect 4580 19119 4629 19125
rect 4985 19159 5043 19165
rect 4985 19125 4997 19159
rect 5031 19156 5043 19159
rect 5074 19156 5080 19168
rect 5031 19128 5080 19156
rect 5031 19125 5043 19128
rect 4985 19119 5043 19125
rect 4580 19116 4586 19119
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1464 18819 1522 18825
rect 1464 18785 1476 18819
rect 1510 18816 1522 18819
rect 1946 18816 1952 18828
rect 1510 18788 1952 18816
rect 1510 18785 1522 18788
rect 1464 18779 1522 18785
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 2476 18819 2534 18825
rect 2476 18785 2488 18819
rect 2522 18816 2534 18819
rect 2682 18816 2688 18828
rect 2522 18788 2688 18816
rect 2522 18785 2534 18788
rect 2476 18779 2534 18785
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 3326 18776 3332 18828
rect 3384 18816 3390 18828
rect 5166 18825 5172 18828
rect 4100 18819 4158 18825
rect 4100 18816 4112 18819
rect 3384 18788 4112 18816
rect 3384 18776 3390 18788
rect 4100 18785 4112 18788
rect 4146 18816 4158 18819
rect 5144 18819 5172 18825
rect 4146 18788 5028 18816
rect 4146 18785 4158 18788
rect 4100 18779 4158 18785
rect 5000 18748 5028 18788
rect 5144 18785 5156 18819
rect 5144 18779 5172 18785
rect 5166 18776 5172 18779
rect 5224 18776 5230 18828
rect 5442 18748 5448 18760
rect 5000 18720 5448 18748
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 3878 18640 3884 18692
rect 3936 18680 3942 18692
rect 5215 18683 5273 18689
rect 5215 18680 5227 18683
rect 3936 18652 5227 18680
rect 3936 18640 3942 18652
rect 5215 18649 5227 18652
rect 5261 18649 5273 18683
rect 5215 18643 5273 18649
rect 1535 18615 1593 18621
rect 1535 18581 1547 18615
rect 1581 18612 1593 18615
rect 1670 18612 1676 18624
rect 1581 18584 1676 18612
rect 1581 18581 1593 18584
rect 1535 18575 1593 18581
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 2547 18615 2605 18621
rect 2547 18612 2559 18615
rect 2188 18584 2559 18612
rect 2188 18572 2194 18584
rect 2547 18581 2559 18584
rect 2593 18581 2605 18615
rect 2547 18575 2605 18581
rect 4154 18572 4160 18624
rect 4212 18621 4218 18624
rect 4212 18615 4261 18621
rect 4212 18581 4215 18615
rect 4249 18581 4261 18615
rect 4212 18575 4261 18581
rect 4212 18572 4218 18575
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1946 18408 1952 18420
rect 1859 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18408 2010 18420
rect 2590 18408 2596 18420
rect 2004 18380 2596 18408
rect 2004 18368 2010 18380
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 3326 18408 3332 18420
rect 3287 18380 3332 18408
rect 3326 18368 3332 18380
rect 3384 18368 3390 18420
rect 1302 18300 1308 18352
rect 1360 18340 1366 18352
rect 4249 18343 4307 18349
rect 4249 18340 4261 18343
rect 1360 18312 4261 18340
rect 1360 18300 1366 18312
rect 4249 18309 4261 18312
rect 4295 18340 4307 18343
rect 8110 18340 8116 18352
rect 4295 18312 8116 18340
rect 4295 18309 4307 18312
rect 4249 18303 4307 18309
rect 1210 18164 1216 18216
rect 1268 18204 1274 18216
rect 1432 18207 1490 18213
rect 1432 18204 1444 18207
rect 1268 18176 1444 18204
rect 1268 18164 1274 18176
rect 1432 18173 1444 18176
rect 1478 18173 1490 18207
rect 1432 18167 1490 18173
rect 2476 18207 2534 18213
rect 2476 18173 2488 18207
rect 2522 18204 2534 18207
rect 2590 18204 2596 18216
rect 2522 18176 2596 18204
rect 2522 18173 2534 18176
rect 2476 18167 2534 18173
rect 1447 18136 1475 18167
rect 2590 18164 2596 18176
rect 2648 18204 2654 18216
rect 2869 18207 2927 18213
rect 2869 18204 2881 18207
rect 2648 18176 2881 18204
rect 2648 18164 2654 18176
rect 2869 18173 2881 18176
rect 2915 18173 2927 18207
rect 2869 18167 2927 18173
rect 3488 18207 3546 18213
rect 3488 18173 3500 18207
rect 3534 18204 3546 18207
rect 4264 18204 4292 18303
rect 8110 18300 8116 18312
rect 8168 18300 8174 18352
rect 5166 18272 5172 18284
rect 5079 18244 5172 18272
rect 5166 18232 5172 18244
rect 5224 18272 5230 18284
rect 8570 18272 8576 18284
rect 5224 18244 8576 18272
rect 5224 18232 5230 18244
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 4468 18207 4526 18213
rect 4468 18204 4480 18207
rect 3534 18176 3832 18204
rect 4264 18176 4480 18204
rect 3534 18173 3546 18176
rect 3488 18167 3546 18173
rect 2225 18139 2283 18145
rect 2225 18136 2237 18139
rect 1447 18108 2237 18136
rect 2225 18105 2237 18108
rect 2271 18105 2283 18139
rect 2225 18099 2283 18105
rect 3804 18080 3832 18176
rect 4468 18173 4480 18176
rect 4514 18173 4526 18207
rect 4468 18167 4526 18173
rect 5496 18207 5554 18213
rect 5496 18173 5508 18207
rect 5542 18204 5554 18207
rect 6917 18207 6975 18213
rect 5542 18176 6132 18204
rect 5542 18173 5554 18176
rect 5496 18167 5554 18173
rect 5583 18139 5641 18145
rect 5583 18105 5595 18139
rect 5629 18136 5641 18139
rect 5994 18136 6000 18148
rect 5629 18108 6000 18136
rect 5629 18105 5641 18108
rect 5583 18099 5641 18105
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 1578 18077 1584 18080
rect 1535 18071 1584 18077
rect 1535 18037 1547 18071
rect 1581 18037 1584 18071
rect 1535 18031 1584 18037
rect 1578 18028 1584 18031
rect 1636 18028 1642 18080
rect 2590 18077 2596 18080
rect 2547 18071 2596 18077
rect 2547 18037 2559 18071
rect 2593 18037 2596 18071
rect 2547 18031 2596 18037
rect 2590 18028 2596 18031
rect 2648 18028 2654 18080
rect 3510 18028 3516 18080
rect 3568 18077 3574 18080
rect 3568 18071 3617 18077
rect 3568 18037 3571 18071
rect 3605 18037 3617 18071
rect 3568 18031 3617 18037
rect 3568 18028 3574 18031
rect 3786 18028 3792 18080
rect 3844 18068 3850 18080
rect 3881 18071 3939 18077
rect 3881 18068 3893 18071
rect 3844 18040 3893 18068
rect 3844 18028 3850 18040
rect 3881 18037 3893 18040
rect 3927 18037 3939 18071
rect 3881 18031 3939 18037
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 4571 18071 4629 18077
rect 4571 18068 4583 18071
rect 4488 18040 4583 18068
rect 4488 18028 4494 18040
rect 4571 18037 4583 18040
rect 4617 18037 4629 18071
rect 4571 18031 4629 18037
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 6104 18068 6132 18176
rect 6917 18173 6929 18207
rect 6963 18173 6975 18207
rect 6917 18167 6975 18173
rect 6932 18136 6960 18167
rect 7466 18136 7472 18148
rect 6932 18108 7472 18136
rect 7466 18096 7472 18108
rect 7524 18096 7530 18148
rect 6178 18068 6184 18080
rect 5951 18040 6184 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 7101 18071 7159 18077
rect 7101 18068 7113 18071
rect 6972 18040 7113 18068
rect 6972 18028 6978 18040
rect 7101 18037 7113 18040
rect 7147 18068 7159 18071
rect 7650 18068 7656 18080
rect 7147 18040 7656 18068
rect 7147 18037 7159 18040
rect 7101 18031 7159 18037
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1946 17728 1952 17740
rect 1907 17700 1952 17728
rect 1946 17688 1952 17700
rect 2004 17688 2010 17740
rect 2133 17731 2191 17737
rect 2133 17728 2145 17731
rect 2056 17700 2145 17728
rect 1394 17620 1400 17672
rect 1452 17660 1458 17672
rect 2056 17660 2084 17700
rect 2133 17697 2145 17700
rect 2179 17697 2191 17731
rect 2133 17691 2191 17697
rect 4408 17731 4466 17737
rect 4408 17697 4420 17731
rect 4454 17728 4466 17731
rect 4798 17728 4804 17740
rect 4454 17700 4804 17728
rect 4454 17697 4466 17700
rect 4408 17691 4466 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 6156 17731 6214 17737
rect 6156 17697 6168 17731
rect 6202 17728 6214 17731
rect 6270 17728 6276 17740
rect 6202 17700 6276 17728
rect 6202 17697 6214 17700
rect 6156 17691 6214 17697
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 8272 17731 8330 17737
rect 8272 17697 8284 17731
rect 8318 17728 8330 17731
rect 8938 17728 8944 17740
rect 8318 17700 8944 17728
rect 8318 17697 8330 17700
rect 8272 17691 8330 17697
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9744 17731 9802 17737
rect 9744 17697 9756 17731
rect 9790 17728 9802 17731
rect 9950 17728 9956 17740
rect 9790 17700 9956 17728
rect 9790 17697 9802 17700
rect 9744 17691 9802 17697
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 2222 17660 2228 17672
rect 1452 17632 2084 17660
rect 2183 17632 2228 17660
rect 1452 17620 1458 17632
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 6454 17620 6460 17672
rect 6512 17660 6518 17672
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 6512 17632 7205 17660
rect 6512 17620 6518 17632
rect 7193 17629 7205 17632
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17660 10747 17663
rect 10962 17660 10968 17672
rect 10735 17632 10968 17660
rect 10735 17629 10747 17632
rect 10689 17623 10747 17629
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 2682 17484 2688 17536
rect 2740 17524 2746 17536
rect 2777 17527 2835 17533
rect 2777 17524 2789 17527
rect 2740 17496 2789 17524
rect 2740 17484 2746 17496
rect 2777 17493 2789 17496
rect 2823 17524 2835 17527
rect 3694 17524 3700 17536
rect 2823 17496 3700 17524
rect 2823 17493 2835 17496
rect 2777 17487 2835 17493
rect 3694 17484 3700 17496
rect 3752 17484 3758 17536
rect 4479 17527 4537 17533
rect 4479 17493 4491 17527
rect 4525 17524 4537 17527
rect 4706 17524 4712 17536
rect 4525 17496 4712 17524
rect 4525 17493 4537 17496
rect 4479 17487 4537 17493
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 6086 17484 6092 17536
rect 6144 17524 6150 17536
rect 6227 17527 6285 17533
rect 6227 17524 6239 17527
rect 6144 17496 6239 17524
rect 6144 17484 6150 17496
rect 6227 17493 6239 17496
rect 6273 17493 6285 17527
rect 6227 17487 6285 17493
rect 8294 17484 8300 17536
rect 8352 17533 8358 17536
rect 9858 17533 9864 17536
rect 8352 17527 8401 17533
rect 8352 17493 8355 17527
rect 8389 17493 8401 17527
rect 8352 17487 8401 17493
rect 9815 17527 9864 17533
rect 9815 17493 9827 17527
rect 9861 17493 9864 17527
rect 9815 17487 9864 17493
rect 8352 17484 8358 17487
rect 9858 17484 9864 17487
rect 9916 17484 9922 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 6270 17320 6276 17332
rect 6227 17292 6276 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 3053 17255 3111 17261
rect 3053 17252 3065 17255
rect 2056 17224 3065 17252
rect 1394 17144 1400 17196
rect 1452 17184 1458 17196
rect 2056 17184 2084 17224
rect 3053 17221 3065 17224
rect 3099 17252 3111 17255
rect 6914 17252 6920 17264
rect 3099 17224 6920 17252
rect 3099 17221 3111 17224
rect 3053 17215 3111 17221
rect 6914 17212 6920 17224
rect 6972 17212 6978 17264
rect 1452 17156 2084 17184
rect 1452 17144 1458 17156
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17085 2007 17119
rect 2056 17116 2084 17156
rect 2133 17119 2191 17125
rect 2133 17116 2145 17119
rect 2056 17088 2145 17116
rect 1949 17079 2007 17085
rect 2133 17085 2145 17088
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 1964 17048 1992 17079
rect 3234 17076 3240 17128
rect 3292 17125 3298 17128
rect 3292 17119 3330 17125
rect 3318 17116 3330 17119
rect 3697 17119 3755 17125
rect 3697 17116 3709 17119
rect 3318 17088 3709 17116
rect 3318 17085 3330 17088
rect 3292 17079 3330 17085
rect 3697 17085 3709 17088
rect 3743 17085 3755 17119
rect 3697 17079 3755 17085
rect 4960 17119 5018 17125
rect 4960 17085 4972 17119
rect 5006 17116 5018 17119
rect 7168 17119 7226 17125
rect 5006 17088 5396 17116
rect 5006 17085 5018 17088
rect 4960 17079 5018 17085
rect 3292 17076 3298 17079
rect 2777 17051 2835 17057
rect 2777 17048 2789 17051
rect 1964 17020 2789 17048
rect 2777 17017 2789 17020
rect 2823 17048 2835 17051
rect 2958 17048 2964 17060
rect 2823 17020 2964 17048
rect 2823 17017 2835 17020
rect 2777 17011 2835 17017
rect 2958 17008 2964 17020
rect 3016 17008 3022 17060
rect 5368 16992 5396 17088
rect 7168 17085 7180 17119
rect 7214 17116 7226 17119
rect 8113 17119 8171 17125
rect 7214 17088 7420 17116
rect 7214 17085 7226 17088
rect 7168 17079 7226 17085
rect 7392 17060 7420 17088
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 9636 17119 9694 17125
rect 9636 17085 9648 17119
rect 9682 17116 9694 17119
rect 10042 17116 10048 17128
rect 9682 17088 10048 17116
rect 9682 17085 9694 17088
rect 9636 17079 9694 17085
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 7561 17051 7619 17057
rect 7561 17048 7573 17051
rect 7432 17020 7573 17048
rect 7432 17008 7438 17020
rect 7561 17017 7573 17020
rect 7607 17017 7619 17051
rect 8128 17048 8156 17079
rect 10042 17076 10048 17088
rect 10100 17116 10106 17128
rect 10413 17119 10471 17125
rect 10413 17116 10425 17119
rect 10100 17088 10425 17116
rect 10100 17076 10106 17088
rect 10413 17085 10425 17088
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 10664 17119 10722 17125
rect 10664 17085 10676 17119
rect 10710 17116 10722 17119
rect 11057 17119 11115 17125
rect 11057 17116 11069 17119
rect 10710 17088 11069 17116
rect 10710 17085 10722 17088
rect 10664 17079 10722 17085
rect 11057 17085 11069 17088
rect 11103 17116 11115 17119
rect 11146 17116 11152 17128
rect 11103 17088 11152 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 13078 17125 13084 17128
rect 13056 17119 13084 17125
rect 13056 17085 13068 17119
rect 13136 17116 13142 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13136 17088 13461 17116
rect 13056 17079 13084 17085
rect 13078 17076 13084 17079
rect 13136 17076 13142 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 14734 17076 14740 17128
rect 14792 17116 14798 17128
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 14792 17088 15025 17116
rect 14792 17076 14798 17088
rect 15013 17085 15025 17088
rect 15059 17116 15071 17119
rect 15473 17119 15531 17125
rect 15473 17116 15485 17119
rect 15059 17088 15485 17116
rect 15059 17085 15071 17088
rect 15013 17079 15071 17085
rect 15473 17085 15485 17088
rect 15519 17085 15531 17119
rect 15473 17079 15531 17085
rect 9030 17048 9036 17060
rect 8128 17020 9036 17048
rect 7561 17011 7619 17017
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 9723 17051 9781 17057
rect 9723 17017 9735 17051
rect 9769 17048 9781 17051
rect 10870 17048 10876 17060
rect 9769 17020 10876 17048
rect 9769 17017 9781 17020
rect 9723 17011 9781 17017
rect 10870 17008 10876 17020
rect 10928 17008 10934 17060
rect 1765 16983 1823 16989
rect 1765 16949 1777 16983
rect 1811 16980 1823 16983
rect 1854 16980 1860 16992
rect 1811 16952 1860 16980
rect 1811 16949 1823 16952
rect 1765 16943 1823 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 3375 16983 3433 16989
rect 3375 16949 3387 16983
rect 3421 16980 3433 16983
rect 3970 16980 3976 16992
rect 3421 16952 3976 16980
rect 3421 16949 3433 16952
rect 3375 16943 3433 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4433 16983 4491 16989
rect 4433 16949 4445 16983
rect 4479 16980 4491 16983
rect 4798 16980 4804 16992
rect 4479 16952 4804 16980
rect 4479 16949 4491 16952
rect 4433 16943 4491 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 5031 16983 5089 16989
rect 5031 16980 5043 16983
rect 4948 16952 5043 16980
rect 4948 16940 4954 16952
rect 5031 16949 5043 16952
rect 5077 16949 5089 16983
rect 5350 16980 5356 16992
rect 5311 16952 5356 16980
rect 5031 16943 5089 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 7239 16983 7297 16989
rect 7239 16949 7251 16983
rect 7285 16980 7297 16983
rect 7466 16980 7472 16992
rect 7285 16952 7472 16980
rect 7285 16949 7297 16952
rect 7239 16943 7297 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 8297 16983 8355 16989
rect 8297 16949 8309 16983
rect 8343 16980 8355 16983
rect 8386 16980 8392 16992
rect 8343 16952 8392 16980
rect 8343 16949 8355 16952
rect 8297 16943 8355 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 8665 16983 8723 16989
rect 8665 16949 8677 16983
rect 8711 16980 8723 16983
rect 8938 16980 8944 16992
rect 8711 16952 8944 16980
rect 8711 16949 8723 16952
rect 8665 16943 8723 16949
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9950 16940 9956 16992
rect 10008 16980 10014 16992
rect 10045 16983 10103 16989
rect 10045 16980 10057 16983
rect 10008 16952 10057 16980
rect 10008 16940 10014 16952
rect 10045 16949 10057 16952
rect 10091 16949 10103 16983
rect 10045 16943 10103 16949
rect 10735 16983 10793 16989
rect 10735 16949 10747 16983
rect 10781 16980 10793 16983
rect 11238 16980 11244 16992
rect 10781 16952 11244 16980
rect 10781 16949 10793 16952
rect 10735 16943 10793 16949
rect 11238 16940 11244 16952
rect 11296 16940 11302 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 13127 16983 13185 16989
rect 13127 16980 13139 16983
rect 12860 16952 13139 16980
rect 12860 16940 12866 16952
rect 13127 16949 13139 16952
rect 13173 16949 13185 16983
rect 13127 16943 13185 16949
rect 15197 16983 15255 16989
rect 15197 16949 15209 16983
rect 15243 16980 15255 16983
rect 16298 16980 16304 16992
rect 15243 16952 16304 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1765 16779 1823 16785
rect 1765 16745 1777 16779
rect 1811 16776 1823 16779
rect 1946 16776 1952 16788
rect 1811 16748 1952 16776
rect 1811 16745 1823 16748
rect 1765 16739 1823 16745
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2038 16736 2044 16788
rect 2096 16736 2102 16788
rect 4706 16776 4712 16788
rect 4667 16748 4712 16776
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 9766 16776 9772 16788
rect 9727 16748 9772 16776
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 13262 16776 13268 16788
rect 13223 16748 13268 16776
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 15473 16779 15531 16785
rect 15473 16745 15485 16779
rect 15519 16776 15531 16779
rect 15930 16776 15936 16788
rect 15519 16748 15936 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 16206 16776 16212 16788
rect 16167 16748 16212 16776
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16485 16779 16543 16785
rect 16485 16745 16497 16779
rect 16531 16745 16543 16779
rect 16485 16739 16543 16745
rect 2056 16708 2084 16736
rect 2225 16711 2283 16717
rect 2225 16708 2237 16711
rect 2056 16680 2237 16708
rect 2056 16584 2084 16680
rect 2225 16677 2237 16680
rect 2271 16677 2283 16711
rect 2225 16671 2283 16677
rect 2317 16711 2375 16717
rect 2317 16677 2329 16711
rect 2363 16708 2375 16711
rect 2682 16708 2688 16720
rect 2363 16680 2688 16708
rect 2363 16677 2375 16680
rect 2317 16671 2375 16677
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 8202 16668 8208 16720
rect 8260 16708 8266 16720
rect 8619 16711 8677 16717
rect 8619 16708 8631 16711
rect 8260 16680 8631 16708
rect 8260 16668 8266 16680
rect 8619 16677 8631 16680
rect 8665 16677 8677 16711
rect 8619 16671 8677 16677
rect 10781 16711 10839 16717
rect 10781 16677 10793 16711
rect 10827 16708 10839 16711
rect 10827 16680 13584 16708
rect 10827 16677 10839 16680
rect 10781 16671 10839 16677
rect 4116 16643 4174 16649
rect 4116 16609 4128 16643
rect 4162 16640 4174 16643
rect 4203 16643 4261 16649
rect 4162 16609 4175 16640
rect 4116 16603 4175 16609
rect 4203 16609 4215 16643
rect 4249 16640 4261 16643
rect 4338 16640 4344 16652
rect 4249 16612 4344 16640
rect 4249 16609 4261 16612
rect 4203 16603 4261 16609
rect 2038 16532 2044 16584
rect 2096 16532 2102 16584
rect 2866 16572 2872 16584
rect 2827 16544 2872 16572
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 4147 16572 4175 16603
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 5258 16649 5264 16652
rect 5128 16643 5186 16649
rect 5128 16609 5140 16643
rect 5174 16640 5186 16643
rect 5215 16643 5264 16649
rect 5174 16609 5187 16640
rect 5128 16603 5187 16609
rect 5215 16609 5227 16643
rect 5261 16609 5264 16643
rect 5215 16603 5264 16609
rect 4614 16572 4620 16584
rect 4147 16544 4620 16572
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 5159 16572 5187 16603
rect 5258 16600 5264 16603
rect 5316 16600 5322 16652
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 6822 16640 6828 16652
rect 6595 16612 6828 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 8478 16600 8484 16652
rect 8536 16649 8542 16652
rect 8536 16643 8574 16649
rect 8562 16609 8574 16643
rect 8536 16603 8574 16609
rect 9217 16643 9275 16649
rect 9217 16609 9229 16643
rect 9263 16640 9275 16643
rect 9582 16640 9588 16652
rect 9263 16612 9588 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 8536 16600 8542 16603
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10134 16640 10140 16652
rect 9999 16612 10140 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16640 10287 16643
rect 10796 16640 10824 16671
rect 10275 16612 10824 16640
rect 11701 16643 11759 16649
rect 10275 16609 10287 16612
rect 10229 16603 10287 16609
rect 11701 16609 11713 16643
rect 11747 16640 11759 16643
rect 11882 16640 11888 16652
rect 11747 16612 11888 16640
rect 11747 16609 11759 16612
rect 11701 16603 11759 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 11992 16649 12020 16680
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 12161 16643 12219 16649
rect 12161 16609 12173 16643
rect 12207 16640 12219 16643
rect 12342 16640 12348 16652
rect 12207 16612 12348 16640
rect 12207 16609 12219 16612
rect 12161 16603 12219 16609
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 13556 16649 13584 16680
rect 16114 16668 16120 16720
rect 16172 16708 16178 16720
rect 16500 16708 16528 16739
rect 16172 16680 16528 16708
rect 16172 16668 16178 16680
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16609 13047 16643
rect 12989 16603 13047 16609
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13630 16640 13636 16652
rect 13587 16612 13636 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 5534 16572 5540 16584
rect 5159 16544 5540 16572
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 13004 16572 13032 16603
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16640 16359 16643
rect 16942 16640 16948 16652
rect 16347 16612 16948 16640
rect 16347 16609 16359 16612
rect 16301 16603 16359 16609
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 12308 16544 13032 16572
rect 12308 16532 12314 16544
rect 6730 16436 6736 16448
rect 6691 16408 6736 16436
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 14185 16439 14243 16445
rect 12492 16408 12537 16436
rect 12492 16396 12498 16408
rect 14185 16405 14197 16439
rect 14231 16436 14243 16439
rect 14366 16436 14372 16448
rect 14231 16408 14372 16436
rect 14231 16405 14243 16408
rect 14185 16399 14243 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2682 16192 2688 16244
rect 2740 16232 2746 16244
rect 3605 16235 3663 16241
rect 3605 16232 3617 16235
rect 2740 16204 3617 16232
rect 2740 16192 2746 16204
rect 3605 16201 3617 16204
rect 3651 16232 3663 16235
rect 4617 16235 4675 16241
rect 4617 16232 4629 16235
rect 3651 16204 4629 16232
rect 3651 16201 3663 16204
rect 3605 16195 3663 16201
rect 4617 16201 4629 16204
rect 4663 16232 4675 16235
rect 4663 16204 5488 16232
rect 4663 16201 4675 16204
rect 4617 16195 4675 16201
rect 4706 16124 4712 16176
rect 4764 16124 4770 16176
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 2332 16068 2605 16096
rect 2332 15969 2360 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2866 16096 2872 16108
rect 2827 16068 2872 16096
rect 2593 16059 2651 16065
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 4724 16096 4752 16124
rect 4801 16099 4859 16105
rect 4801 16096 4813 16099
rect 4724 16068 4813 16096
rect 4801 16065 4813 16068
rect 4847 16065 4859 16099
rect 5074 16096 5080 16108
rect 5035 16068 5080 16096
rect 4801 16059 4859 16065
rect 5074 16056 5080 16068
rect 5132 16056 5138 16108
rect 4614 15988 4620 16040
rect 4672 15988 4678 16040
rect 1489 15963 1547 15969
rect 1489 15929 1501 15963
rect 1535 15960 1547 15963
rect 2317 15963 2375 15969
rect 2317 15960 2329 15963
rect 1535 15932 2329 15960
rect 1535 15929 1547 15932
rect 1489 15923 1547 15929
rect 2317 15929 2329 15932
rect 2363 15929 2375 15963
rect 2682 15960 2688 15972
rect 2643 15932 2688 15960
rect 2317 15923 2375 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1452 15864 1961 15892
rect 1452 15852 1458 15864
rect 1949 15861 1961 15864
rect 1995 15861 2007 15895
rect 1949 15855 2007 15861
rect 4157 15895 4215 15901
rect 4157 15861 4169 15895
rect 4203 15892 4215 15895
rect 4632 15892 4660 15988
rect 4893 15963 4951 15969
rect 4893 15929 4905 15963
rect 4939 15960 4951 15963
rect 5460 15960 5488 16204
rect 8478 16192 8484 16244
rect 8536 16232 8542 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 8536 16204 8953 16232
rect 8536 16192 8542 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 10134 16232 10140 16244
rect 10095 16204 10140 16232
rect 8941 16195 8999 16201
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 24762 16192 24768 16244
rect 24820 16232 24826 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 24820 16204 25053 16232
rect 24820 16192 24826 16204
rect 25041 16201 25053 16204
rect 25087 16201 25099 16235
rect 25041 16195 25099 16201
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 12434 16096 12440 16108
rect 9640 16068 12440 16096
rect 9640 16056 9646 16068
rect 7168 16031 7226 16037
rect 7168 15997 7180 16031
rect 7214 16028 7226 16031
rect 7214 16000 7696 16028
rect 7214 15997 7226 16000
rect 7168 15991 7226 15997
rect 6270 15960 6276 15972
rect 4939 15932 6276 15960
rect 4939 15929 4951 15932
rect 4893 15923 4951 15929
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 5626 15892 5632 15904
rect 4203 15864 5632 15892
rect 4203 15861 4215 15864
rect 4157 15855 4215 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 5813 15895 5871 15901
rect 5813 15892 5825 15895
rect 5776 15864 5825 15892
rect 5776 15852 5782 15864
rect 5813 15861 5825 15864
rect 5859 15892 5871 15895
rect 6546 15892 6552 15904
rect 5859 15864 6552 15892
rect 5859 15861 5871 15864
rect 5813 15855 5871 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 6822 15892 6828 15904
rect 6687 15864 6828 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7282 15901 7288 15904
rect 7239 15895 7288 15901
rect 7239 15861 7251 15895
rect 7285 15861 7288 15895
rect 7239 15855 7288 15861
rect 7282 15852 7288 15855
rect 7340 15852 7346 15904
rect 7668 15901 7696 16000
rect 8110 15988 8116 16040
rect 8168 16037 8174 16040
rect 8168 16031 8206 16037
rect 8194 16028 8206 16031
rect 8573 16031 8631 16037
rect 8573 16028 8585 16031
rect 8194 16000 8585 16028
rect 8194 15997 8206 16000
rect 8168 15991 8206 15997
rect 8573 15997 8585 16000
rect 8619 15997 8631 16031
rect 9122 16028 9128 16040
rect 9083 16000 9128 16028
rect 8573 15991 8631 15997
rect 8168 15988 8174 15991
rect 9122 15988 9128 16000
rect 9180 15988 9186 16040
rect 9692 16037 9720 16068
rect 12434 16056 12440 16068
rect 12492 16096 12498 16108
rect 14642 16096 14648 16108
rect 12492 16068 14412 16096
rect 14603 16068 14648 16096
rect 12492 16056 12498 16068
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 15997 10747 16031
rect 10689 15991 10747 15997
rect 11241 16031 11299 16037
rect 11241 15997 11253 16031
rect 11287 16028 11299 16031
rect 11330 16028 11336 16040
rect 11287 16000 11336 16028
rect 11287 15997 11299 16000
rect 11241 15991 11299 15997
rect 9140 15960 9168 15988
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 9140 15932 10517 15960
rect 10505 15929 10517 15932
rect 10551 15960 10563 15963
rect 10704 15960 10732 15991
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 12158 16028 12164 16040
rect 11572 16000 12164 16028
rect 11572 15988 11578 16000
rect 12158 15988 12164 16000
rect 12216 16028 12222 16040
rect 13004 16037 13032 16068
rect 14384 16040 14412 16068
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 16206 16096 16212 16108
rect 16167 16068 16212 16096
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 12529 16031 12587 16037
rect 12529 16028 12541 16031
rect 12216 16000 12541 16028
rect 12216 15988 12222 16000
rect 12529 15997 12541 16000
rect 12575 15997 12587 16031
rect 12529 15991 12587 15997
rect 12989 16031 13047 16037
rect 12989 15997 13001 16031
rect 13035 15997 13047 16031
rect 14274 16028 14280 16040
rect 14235 16000 14280 16028
rect 12989 15991 13047 15997
rect 11422 15960 11428 15972
rect 10551 15932 10732 15960
rect 11383 15932 11428 15960
rect 10551 15929 10563 15932
rect 10505 15923 10563 15929
rect 11422 15920 11428 15932
rect 11480 15920 11486 15972
rect 12544 15960 12572 15991
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 14366 15988 14372 16040
rect 14424 16028 14430 16040
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 14424 16000 14565 16028
rect 14424 15988 14430 16000
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 24648 16031 24706 16037
rect 18095 16000 18644 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 12544 15932 13461 15960
rect 13449 15929 13461 15932
rect 13495 15929 13507 15963
rect 13449 15923 13507 15929
rect 13814 15920 13820 15972
rect 13872 15960 13878 15972
rect 15933 15963 15991 15969
rect 15933 15960 15945 15963
rect 13872 15932 15945 15960
rect 13872 15920 13878 15932
rect 15933 15929 15945 15932
rect 15979 15960 15991 15963
rect 16301 15963 16359 15969
rect 16301 15960 16313 15963
rect 15979 15932 16313 15960
rect 15979 15929 15991 15932
rect 15933 15923 15991 15929
rect 16301 15929 16313 15932
rect 16347 15929 16359 15963
rect 16850 15960 16856 15972
rect 16811 15932 16856 15960
rect 16301 15923 16359 15929
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15892 7711 15895
rect 7926 15892 7932 15904
rect 7699 15864 7932 15892
rect 7699 15861 7711 15864
rect 7653 15855 7711 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 8251 15895 8309 15901
rect 8251 15892 8263 15895
rect 8168 15864 8263 15892
rect 8168 15852 8174 15864
rect 8251 15861 8263 15864
rect 8297 15861 8309 15895
rect 9398 15892 9404 15904
rect 9359 15864 9404 15892
rect 8251 15855 8309 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 11793 15895 11851 15901
rect 11793 15861 11805 15895
rect 11839 15892 11851 15895
rect 11882 15892 11888 15904
rect 11839 15864 11888 15892
rect 11839 15861 11851 15864
rect 11793 15855 11851 15861
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12529 15895 12587 15901
rect 12529 15861 12541 15895
rect 12575 15892 12587 15895
rect 12618 15892 12624 15904
rect 12575 15864 12624 15892
rect 12575 15861 12587 15864
rect 12529 15855 12587 15861
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 14001 15895 14059 15901
rect 14001 15861 14013 15895
rect 14047 15892 14059 15895
rect 14274 15892 14280 15904
rect 14047 15864 14280 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 14274 15852 14280 15864
rect 14332 15892 14338 15904
rect 14458 15892 14464 15904
rect 14332 15864 14464 15892
rect 14332 15852 14338 15864
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15381 15895 15439 15901
rect 15381 15892 15393 15895
rect 15344 15864 15393 15892
rect 15344 15852 15350 15864
rect 15381 15861 15393 15864
rect 15427 15892 15439 15895
rect 15746 15892 15752 15904
rect 15427 15864 15752 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 16942 15852 16948 15904
rect 17000 15892 17006 15904
rect 17129 15895 17187 15901
rect 17129 15892 17141 15895
rect 17000 15864 17141 15892
rect 17000 15852 17006 15864
rect 17129 15861 17141 15864
rect 17175 15861 17187 15895
rect 17129 15855 17187 15861
rect 18233 15895 18291 15901
rect 18233 15861 18245 15895
rect 18279 15892 18291 15895
rect 18506 15892 18512 15904
rect 18279 15864 18512 15892
rect 18279 15861 18291 15864
rect 18233 15855 18291 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 18616 15901 18644 16000
rect 24648 15997 24660 16031
rect 24694 16028 24706 16031
rect 24762 16028 24768 16040
rect 24694 16000 24768 16028
rect 24694 15997 24706 16000
rect 24648 15991 24706 15997
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 18601 15895 18659 15901
rect 18601 15861 18613 15895
rect 18647 15892 18659 15895
rect 18782 15892 18788 15904
rect 18647 15864 18788 15892
rect 18647 15861 18659 15864
rect 18601 15855 18659 15861
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 19058 15892 19064 15904
rect 19019 15864 19064 15892
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 24719 15895 24777 15901
rect 24719 15892 24731 15895
rect 23532 15864 24731 15892
rect 23532 15852 23538 15864
rect 24719 15861 24731 15864
rect 24765 15861 24777 15895
rect 24719 15855 24777 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1210 15648 1216 15700
rect 1268 15688 1274 15700
rect 1486 15688 1492 15700
rect 1268 15660 1492 15688
rect 1268 15648 1274 15660
rect 1486 15648 1492 15660
rect 1544 15648 1550 15700
rect 1673 15691 1731 15697
rect 1673 15657 1685 15691
rect 1719 15688 1731 15691
rect 2038 15688 2044 15700
rect 1719 15660 2044 15688
rect 1719 15657 1731 15660
rect 1673 15651 1731 15657
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 2682 15648 2688 15700
rect 2740 15688 2746 15700
rect 2958 15688 2964 15700
rect 2740 15660 2964 15688
rect 2740 15648 2746 15660
rect 2958 15648 2964 15660
rect 3016 15688 3022 15700
rect 3145 15691 3203 15697
rect 3145 15688 3157 15691
rect 3016 15660 3157 15688
rect 3016 15648 3022 15660
rect 3145 15657 3157 15660
rect 3191 15688 3203 15691
rect 3191 15660 4292 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 2314 15620 2320 15632
rect 2275 15592 2320 15620
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 2866 15620 2872 15632
rect 2827 15592 2872 15620
rect 2866 15580 2872 15592
rect 2924 15620 2930 15632
rect 4264 15629 4292 15660
rect 5166 15648 5172 15700
rect 5224 15688 5230 15700
rect 5626 15688 5632 15700
rect 5224 15660 5632 15688
rect 5224 15648 5230 15660
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 11790 15688 11796 15700
rect 11751 15660 11796 15688
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 3513 15623 3571 15629
rect 3513 15620 3525 15623
rect 2924 15592 3525 15620
rect 2924 15580 2930 15592
rect 3513 15589 3525 15592
rect 3559 15589 3571 15623
rect 3513 15583 3571 15589
rect 4249 15623 4307 15629
rect 4249 15589 4261 15623
rect 4295 15589 4307 15623
rect 6086 15620 6092 15632
rect 6047 15592 6092 15620
rect 4249 15583 4307 15589
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 6270 15620 6276 15632
rect 6227 15592 6276 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 6270 15580 6276 15592
rect 6328 15580 6334 15632
rect 10226 15580 10232 15632
rect 10284 15620 10290 15632
rect 10321 15623 10379 15629
rect 10321 15620 10333 15623
rect 10284 15592 10333 15620
rect 10284 15580 10290 15592
rect 10321 15589 10333 15592
rect 10367 15589 10379 15623
rect 13814 15620 13820 15632
rect 13775 15592 13820 15620
rect 10321 15583 10379 15589
rect 13814 15580 13820 15592
rect 13872 15580 13878 15632
rect 15838 15580 15844 15632
rect 15896 15620 15902 15632
rect 16301 15623 16359 15629
rect 16301 15620 16313 15623
rect 15896 15592 16313 15620
rect 15896 15580 15902 15592
rect 16301 15589 16313 15592
rect 16347 15589 16359 15623
rect 17770 15620 17776 15632
rect 17731 15592 17776 15620
rect 16301 15583 16359 15589
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 17862 15580 17868 15632
rect 17920 15620 17926 15632
rect 17920 15592 17965 15620
rect 17920 15580 17926 15592
rect 7834 15512 7840 15564
rect 7892 15552 7898 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7892 15524 8033 15552
rect 7892 15512 7898 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15521 8539 15555
rect 11882 15552 11888 15564
rect 11843 15524 11888 15552
rect 8481 15515 8539 15521
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2225 15487 2283 15493
rect 2225 15484 2237 15487
rect 2087 15456 2237 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 2225 15453 2237 15456
rect 2271 15484 2283 15487
rect 2406 15484 2412 15496
rect 2271 15456 2412 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4246 15484 4252 15496
rect 4203 15456 4252 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 4172 15416 4200 15447
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 4798 15484 4804 15496
rect 4759 15456 4804 15484
rect 4798 15444 4804 15456
rect 4856 15484 4862 15496
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 4856 15456 6377 15484
rect 4856 15444 4862 15456
rect 6365 15453 6377 15456
rect 6411 15484 6423 15487
rect 6914 15484 6920 15496
rect 6411 15456 6920 15484
rect 6411 15453 6423 15456
rect 6365 15447 6423 15453
rect 6914 15444 6920 15456
rect 6972 15484 6978 15496
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6972 15456 7021 15484
rect 6972 15444 6978 15456
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 4120 15388 4200 15416
rect 4120 15376 4126 15388
rect 8018 15376 8024 15428
rect 8076 15416 8082 15428
rect 8496 15416 8524 15515
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 12250 15552 12256 15564
rect 12211 15524 12256 15552
rect 12250 15512 12256 15524
rect 12308 15552 12314 15564
rect 12434 15552 12440 15564
rect 12308 15524 12440 15552
rect 12308 15512 12314 15524
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 9674 15484 9680 15496
rect 8803 15456 9680 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 10152 15456 10241 15484
rect 10152 15428 10180 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 13722 15484 13728 15496
rect 13683 15456 13728 15484
rect 10229 15447 10287 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 16206 15484 16212 15496
rect 16119 15456 16212 15484
rect 16206 15444 16212 15456
rect 16264 15484 16270 15496
rect 16482 15484 16488 15496
rect 16264 15456 16488 15484
rect 16264 15444 16270 15456
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 16850 15484 16856 15496
rect 16763 15456 16856 15484
rect 16850 15444 16856 15456
rect 16908 15484 16914 15496
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 16908 15456 18061 15484
rect 16908 15444 16914 15456
rect 18049 15453 18061 15456
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 20070 15484 20076 15496
rect 19475 15456 20076 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15484 21603 15487
rect 21726 15484 21732 15496
rect 21591 15456 21732 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 21726 15444 21732 15456
rect 21784 15444 21790 15496
rect 9861 15419 9919 15425
rect 9861 15416 9873 15419
rect 8076 15388 9873 15416
rect 8076 15376 8082 15388
rect 9861 15385 9873 15388
rect 9907 15385 9919 15419
rect 9861 15379 9919 15385
rect 9876 15348 9904 15379
rect 10134 15376 10140 15428
rect 10192 15376 10198 15428
rect 10781 15419 10839 15425
rect 10781 15385 10793 15419
rect 10827 15416 10839 15419
rect 11054 15416 11060 15428
rect 10827 15388 11060 15416
rect 10827 15385 10839 15388
rect 10781 15379 10839 15385
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 13081 15419 13139 15425
rect 13081 15416 13093 15419
rect 11440 15388 13093 15416
rect 11330 15348 11336 15360
rect 9876 15320 11336 15348
rect 11330 15308 11336 15320
rect 11388 15348 11394 15360
rect 11440 15357 11468 15388
rect 13081 15385 13093 15388
rect 13127 15416 13139 15419
rect 13630 15416 13636 15428
rect 13127 15388 13636 15416
rect 13127 15385 13139 15388
rect 13081 15379 13139 15385
rect 13630 15376 13636 15388
rect 13688 15416 13694 15428
rect 13906 15416 13912 15428
rect 13688 15388 13912 15416
rect 13688 15376 13694 15388
rect 13906 15376 13912 15388
rect 13964 15376 13970 15428
rect 14277 15419 14335 15425
rect 14277 15385 14289 15419
rect 14323 15385 14335 15419
rect 14277 15379 14335 15385
rect 11425 15351 11483 15357
rect 11425 15348 11437 15351
rect 11388 15320 11437 15348
rect 11388 15308 11394 15320
rect 11425 15317 11437 15320
rect 11471 15317 11483 15351
rect 11425 15311 11483 15317
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13357 15351 13415 15357
rect 13357 15348 13369 15351
rect 12768 15320 13369 15348
rect 12768 15308 12774 15320
rect 13357 15317 13369 15320
rect 13403 15317 13415 15351
rect 14292 15348 14320 15379
rect 14550 15348 14556 15360
rect 14292 15320 14556 15348
rect 13357 15311 13415 15317
rect 14550 15308 14556 15320
rect 14608 15348 14614 15360
rect 14645 15351 14703 15357
rect 14645 15348 14657 15351
rect 14608 15320 14657 15348
rect 14608 15308 14614 15320
rect 14645 15317 14657 15320
rect 14691 15317 14703 15351
rect 14645 15311 14703 15317
rect 15749 15351 15807 15357
rect 15749 15317 15761 15351
rect 15795 15348 15807 15351
rect 15838 15348 15844 15360
rect 15795 15320 15844 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 15838 15308 15844 15320
rect 15896 15308 15902 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2774 15144 2780 15156
rect 1995 15116 2780 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 1464 14943 1522 14949
rect 1464 14909 1476 14943
rect 1510 14940 1522 14943
rect 1964 14940 1992 15107
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 6086 15144 6092 15156
rect 5767 15116 6092 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 10226 15144 10232 15156
rect 10187 15116 10232 15144
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 12250 15144 12256 15156
rect 12211 15116 12256 15144
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 13630 15144 13636 15156
rect 13591 15116 13636 15144
rect 13630 15104 13636 15116
rect 13688 15104 13694 15156
rect 15197 15147 15255 15153
rect 15197 15113 15209 15147
rect 15243 15144 15255 15147
rect 15286 15144 15292 15156
rect 15243 15116 15292 15144
rect 15243 15113 15255 15116
rect 15197 15107 15255 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 17405 15147 17463 15153
rect 17405 15113 17417 15147
rect 17451 15144 17463 15147
rect 17770 15144 17776 15156
rect 17451 15116 17776 15144
rect 17451 15113 17463 15116
rect 17405 15107 17463 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 2314 15076 2320 15088
rect 2275 15048 2320 15076
rect 2314 15036 2320 15048
rect 2372 15036 2378 15088
rect 2958 15036 2964 15088
rect 3016 15076 3022 15088
rect 3697 15079 3755 15085
rect 3697 15076 3709 15079
rect 3016 15048 3709 15076
rect 3016 15036 3022 15048
rect 3697 15045 3709 15048
rect 3743 15076 3755 15079
rect 4065 15079 4123 15085
rect 4065 15076 4077 15079
rect 3743 15048 4077 15076
rect 3743 15045 3755 15048
rect 3697 15039 3755 15045
rect 4065 15045 4077 15048
rect 4111 15045 4123 15079
rect 4065 15039 4123 15045
rect 19613 15079 19671 15085
rect 19613 15045 19625 15079
rect 19659 15076 19671 15079
rect 20162 15076 20168 15088
rect 19659 15048 20168 15076
rect 19659 15045 19671 15048
rect 19613 15039 19671 15045
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 2866 15008 2872 15020
rect 2823 14980 2872 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 1510 14912 1992 14940
rect 1510 14909 1522 14912
rect 1464 14903 1522 14909
rect 2869 14875 2927 14881
rect 2869 14841 2881 14875
rect 2915 14872 2927 14875
rect 3234 14872 3240 14884
rect 2915 14844 3240 14872
rect 2915 14841 2927 14844
rect 2869 14835 2927 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 3421 14875 3479 14881
rect 3421 14841 3433 14875
rect 3467 14841 3479 14875
rect 4080 14872 4108 15039
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4430 15008 4436 15020
rect 4387 14980 4436 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4430 14968 4436 14980
rect 4488 15008 4494 15020
rect 5261 15011 5319 15017
rect 5261 15008 5273 15011
rect 4488 14980 5273 15008
rect 4488 14968 4494 14980
rect 5261 14977 5273 14980
rect 5307 14977 5319 15011
rect 6914 15008 6920 15020
rect 6875 14980 6920 15008
rect 5261 14971 5319 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7190 15008 7196 15020
rect 7151 14980 7196 15008
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 9582 15008 9588 15020
rect 9416 14980 9588 15008
rect 9416 14949 9444 14980
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 15008 10931 15011
rect 11238 15008 11244 15020
rect 10919 14980 11244 15008
rect 10919 14977 10931 14980
rect 10873 14971 10931 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 12621 15011 12679 15017
rect 12621 15008 12633 15011
rect 11532 14980 12633 15008
rect 8849 14943 8907 14949
rect 8849 14940 8861 14943
rect 8680 14912 8861 14940
rect 4433 14875 4491 14881
rect 4433 14872 4445 14875
rect 4080 14844 4445 14872
rect 3421 14835 3479 14841
rect 4433 14841 4445 14844
rect 4479 14841 4491 14875
rect 4433 14835 4491 14841
rect 4985 14875 5043 14881
rect 4985 14841 4997 14875
rect 5031 14872 5043 14875
rect 5074 14872 5080 14884
rect 5031 14844 5080 14872
rect 5031 14841 5043 14844
rect 4985 14835 5043 14841
rect 1535 14807 1593 14813
rect 1535 14773 1547 14807
rect 1581 14804 1593 14807
rect 2406 14804 2412 14816
rect 1581 14776 2412 14804
rect 1581 14773 1593 14776
rect 1535 14767 1593 14773
rect 2406 14764 2412 14776
rect 2464 14764 2470 14816
rect 3436 14804 3464 14835
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 7064 14844 7109 14872
rect 7064 14832 7070 14844
rect 3878 14804 3884 14816
rect 3436 14776 3884 14804
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 6086 14804 6092 14816
rect 6047 14776 6092 14804
rect 6086 14764 6092 14776
rect 6144 14804 6150 14816
rect 6270 14804 6276 14816
rect 6144 14776 6276 14804
rect 6144 14764 6150 14776
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 6641 14807 6699 14813
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 7024 14804 7052 14832
rect 6687 14776 7052 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 7834 14764 7840 14816
rect 7892 14804 7898 14816
rect 8680 14813 8708 14912
rect 8849 14909 8861 14912
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 9585 14875 9643 14881
rect 9585 14872 9597 14875
rect 9548 14844 9597 14872
rect 9548 14832 9554 14844
rect 9585 14841 9597 14844
rect 9631 14841 9643 14875
rect 9585 14835 9643 14841
rect 10965 14875 11023 14881
rect 10965 14841 10977 14875
rect 11011 14841 11023 14875
rect 10965 14835 11023 14841
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7892 14776 8033 14804
rect 7892 14764 7898 14776
rect 8021 14773 8033 14776
rect 8067 14804 8079 14807
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8067 14776 8677 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 10980 14804 11008 14835
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11532 14881 11560 14980
rect 12621 14977 12633 14980
rect 12667 15008 12679 15011
rect 12710 15008 12716 15020
rect 12667 14980 12716 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 15008 14243 15011
rect 14550 15008 14556 15020
rect 14231 14980 14556 15008
rect 14231 14977 14243 14980
rect 14185 14971 14243 14977
rect 14550 14968 14556 14980
rect 14608 15008 14614 15020
rect 16025 15011 16083 15017
rect 16025 15008 16037 15011
rect 14608 14980 16037 15008
rect 14608 14968 14614 14980
rect 16025 14977 16037 14980
rect 16071 14977 16083 15011
rect 16025 14971 16083 14977
rect 17773 15011 17831 15017
rect 17773 14977 17785 15011
rect 17819 15008 17831 15011
rect 17862 15008 17868 15020
rect 17819 14980 17868 15008
rect 17819 14977 17831 14980
rect 17773 14971 17831 14977
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 19061 14943 19119 14949
rect 18095 14912 18552 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 11112 14844 11529 14872
rect 11112 14832 11118 14844
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 12250 14872 12256 14884
rect 11517 14835 11575 14841
rect 11624 14844 12256 14872
rect 11624 14804 11652 14844
rect 12250 14832 12256 14844
rect 12308 14832 12314 14884
rect 12710 14832 12716 14884
rect 12768 14872 12774 14884
rect 13265 14875 13323 14881
rect 12768 14844 12813 14872
rect 12768 14832 12774 14844
rect 13265 14841 13277 14875
rect 13311 14872 13323 14875
rect 14277 14875 14335 14881
rect 13311 14844 14228 14872
rect 13311 14841 13323 14844
rect 13265 14835 13323 14841
rect 11882 14804 11888 14816
rect 10735 14776 11652 14804
rect 11843 14776 11888 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 14200 14804 14228 14844
rect 14277 14841 14289 14875
rect 14323 14872 14335 14875
rect 14366 14872 14372 14884
rect 14323 14844 14372 14872
rect 14323 14841 14335 14844
rect 14277 14835 14335 14841
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 14826 14872 14832 14884
rect 14787 14844 14832 14872
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 15749 14875 15807 14881
rect 15749 14872 15761 14875
rect 15488 14844 15761 14872
rect 14844 14804 14872 14832
rect 14200 14776 14872 14804
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 15488 14813 15516 14844
rect 15749 14841 15761 14844
rect 15795 14841 15807 14875
rect 15749 14835 15807 14841
rect 15838 14832 15844 14884
rect 15896 14872 15902 14884
rect 15896 14844 15941 14872
rect 15896 14832 15902 14844
rect 15473 14807 15531 14813
rect 15473 14804 15485 14807
rect 15436 14776 15485 14804
rect 15436 14764 15442 14776
rect 15473 14773 15485 14776
rect 15519 14773 15531 14807
rect 15856 14804 15884 14832
rect 18524 14816 18552 14912
rect 19061 14909 19073 14943
rect 19107 14940 19119 14943
rect 19628 14940 19656 15039
rect 20162 15036 20168 15048
rect 20220 15036 20226 15088
rect 19107 14912 19656 14940
rect 20140 14943 20198 14949
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 20140 14909 20152 14943
rect 20186 14940 20198 14943
rect 20186 14912 20576 14940
rect 20186 14909 20198 14912
rect 20140 14903 20198 14909
rect 20548 14816 20576 14912
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 21304 14943 21362 14949
rect 21304 14940 21316 14943
rect 20772 14912 21316 14940
rect 20772 14900 20778 14912
rect 21304 14909 21316 14912
rect 21350 14940 21362 14943
rect 21729 14943 21787 14949
rect 21729 14940 21741 14943
rect 21350 14912 21741 14940
rect 21350 14909 21362 14912
rect 21304 14903 21362 14909
rect 21729 14909 21741 14912
rect 21775 14909 21787 14943
rect 21729 14903 21787 14909
rect 23820 14943 23878 14949
rect 23820 14909 23832 14943
rect 23866 14940 23878 14943
rect 23866 14909 23888 14940
rect 23820 14903 23888 14909
rect 23860 14872 23888 14903
rect 23934 14900 23940 14952
rect 23992 14940 23998 14952
rect 24765 14943 24823 14949
rect 24765 14940 24777 14943
rect 23992 14912 24777 14940
rect 23992 14900 23998 14912
rect 24765 14909 24777 14912
rect 24811 14909 24823 14943
rect 24765 14903 24823 14909
rect 23860 14844 24348 14872
rect 16669 14807 16727 14813
rect 16669 14804 16681 14807
rect 15856 14776 16681 14804
rect 15473 14767 15531 14773
rect 16669 14773 16681 14776
rect 16715 14773 16727 14807
rect 16669 14767 16727 14773
rect 18233 14807 18291 14813
rect 18233 14773 18245 14807
rect 18279 14804 18291 14807
rect 18322 14804 18328 14816
rect 18279 14776 18328 14804
rect 18279 14773 18291 14776
rect 18233 14767 18291 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 18506 14804 18512 14816
rect 18467 14776 18512 14804
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 18966 14764 18972 14816
rect 19024 14804 19030 14816
rect 20254 14813 20260 14816
rect 19245 14807 19303 14813
rect 19245 14804 19257 14807
rect 19024 14776 19257 14804
rect 19024 14764 19030 14776
rect 19245 14773 19257 14776
rect 19291 14773 19303 14807
rect 19245 14767 19303 14773
rect 20211 14807 20260 14813
rect 20211 14773 20223 14807
rect 20257 14773 20260 14807
rect 20211 14767 20260 14773
rect 20254 14764 20260 14767
rect 20312 14764 20318 14816
rect 20530 14804 20536 14816
rect 20491 14776 20536 14804
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 21450 14813 21456 14816
rect 21407 14807 21456 14813
rect 21407 14773 21419 14807
rect 21453 14773 21456 14807
rect 21407 14767 21456 14773
rect 21450 14764 21456 14767
rect 21508 14764 21514 14816
rect 22278 14804 22284 14816
rect 22239 14776 22284 14804
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 23891 14807 23949 14813
rect 23891 14773 23903 14807
rect 23937 14804 23949 14807
rect 24118 14804 24124 14816
rect 23937 14776 24124 14804
rect 23937 14773 23949 14776
rect 23891 14767 23949 14773
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 24320 14813 24348 14844
rect 24305 14807 24363 14813
rect 24305 14773 24317 14807
rect 24351 14804 24363 14807
rect 24946 14804 24952 14816
rect 24351 14776 24952 14804
rect 24351 14773 24363 14776
rect 24305 14767 24363 14773
rect 24946 14764 24952 14776
rect 25004 14764 25010 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1949 14603 2007 14609
rect 1949 14569 1961 14603
rect 1995 14600 2007 14603
rect 2222 14600 2228 14612
rect 1995 14572 2228 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 3234 14600 3240 14612
rect 3195 14572 3240 14600
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4062 14600 4068 14612
rect 3927 14572 4068 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 6086 14560 6092 14612
rect 6144 14600 6150 14612
rect 6917 14603 6975 14609
rect 6917 14600 6929 14603
rect 6144 14572 6929 14600
rect 6144 14560 6150 14572
rect 6917 14569 6929 14572
rect 6963 14569 6975 14603
rect 6917 14563 6975 14569
rect 7929 14603 7987 14609
rect 7929 14569 7941 14603
rect 7975 14600 7987 14603
rect 8018 14600 8024 14612
rect 7975 14572 8024 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 9125 14603 9183 14609
rect 9125 14569 9137 14603
rect 9171 14600 9183 14603
rect 9582 14600 9588 14612
rect 9171 14572 9588 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 2362 14535 2420 14541
rect 2362 14501 2374 14535
rect 2408 14501 2420 14535
rect 4246 14532 4252 14544
rect 4207 14504 4252 14532
rect 2362 14495 2420 14501
rect 1854 14424 1860 14476
rect 1912 14464 1918 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1912 14436 2053 14464
rect 1912 14424 1918 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2377 14464 2405 14495
rect 4246 14492 4252 14504
rect 4304 14492 4310 14544
rect 4798 14532 4804 14544
rect 4759 14504 4804 14532
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 6270 14492 6276 14544
rect 6328 14541 6334 14544
rect 6328 14535 6376 14541
rect 6328 14501 6330 14535
rect 6364 14501 6376 14535
rect 8662 14532 8668 14544
rect 6328 14495 6376 14501
rect 8312 14504 8668 14532
rect 6328 14492 6334 14495
rect 8312 14476 8340 14504
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 8294 14464 8300 14476
rect 2041 14427 2099 14433
rect 2332 14436 2405 14464
rect 8207 14436 8300 14464
rect 2332 14408 2360 14436
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8536 14436 8585 14464
rect 8536 14424 8542 14436
rect 8573 14433 8585 14436
rect 8619 14464 8631 14467
rect 9140 14464 9168 14563
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 12345 14603 12403 14609
rect 12345 14600 12357 14603
rect 12308 14572 12357 14600
rect 12308 14560 12314 14572
rect 12345 14569 12357 14572
rect 12391 14569 12403 14603
rect 12345 14563 12403 14569
rect 14093 14603 14151 14609
rect 14093 14569 14105 14603
rect 14139 14600 14151 14603
rect 14366 14600 14372 14612
rect 14139 14572 14372 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15427 14603 15485 14609
rect 15427 14600 15439 14603
rect 15344 14572 15439 14600
rect 15344 14560 15350 14572
rect 15427 14569 15439 14572
rect 15473 14569 15485 14603
rect 16206 14600 16212 14612
rect 16167 14572 16212 14600
rect 15427 14563 15485 14569
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 17954 14600 17960 14612
rect 17915 14572 17960 14600
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 10039 14535 10097 14541
rect 10039 14501 10051 14535
rect 10085 14532 10097 14535
rect 10226 14532 10232 14544
rect 10085 14504 10232 14532
rect 10085 14501 10097 14504
rect 10039 14495 10097 14501
rect 10226 14492 10232 14504
rect 10284 14532 10290 14544
rect 13538 14541 13544 14544
rect 11746 14535 11804 14541
rect 11746 14532 11758 14535
rect 10284 14504 11758 14532
rect 10284 14492 10290 14504
rect 11746 14501 11758 14504
rect 11792 14501 11804 14535
rect 13535 14532 13544 14541
rect 13499 14504 13544 14532
rect 11746 14495 11804 14501
rect 13535 14495 13544 14504
rect 13538 14492 13544 14495
rect 13596 14492 13602 14544
rect 16482 14532 16488 14544
rect 16443 14504 16488 14532
rect 16482 14492 16488 14504
rect 16540 14492 16546 14544
rect 9674 14464 9680 14476
rect 8619 14436 9168 14464
rect 9635 14436 9680 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9674 14424 9680 14436
rect 9732 14464 9738 14476
rect 10870 14464 10876 14476
rect 9732 14436 10876 14464
rect 9732 14424 9738 14436
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11422 14464 11428 14476
rect 11383 14436 11428 14464
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 13262 14464 13268 14476
rect 13219 14436 13268 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 15356 14467 15414 14473
rect 15356 14433 15368 14467
rect 15402 14464 15414 14467
rect 15470 14464 15476 14476
rect 15402 14436 15476 14464
rect 15402 14433 15414 14436
rect 15356 14427 15414 14433
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 17402 14424 17408 14476
rect 17460 14464 17466 14476
rect 17865 14467 17923 14473
rect 17865 14464 17877 14467
rect 17460 14436 17877 14464
rect 17460 14424 17466 14436
rect 17865 14433 17877 14436
rect 17911 14433 17923 14467
rect 17865 14427 17923 14433
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 18196 14436 18337 14464
rect 18196 14424 18202 14436
rect 18325 14433 18337 14436
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 19518 14424 19524 14476
rect 19576 14473 19582 14476
rect 19576 14467 19614 14473
rect 19602 14433 19614 14467
rect 19576 14427 19614 14433
rect 19576 14424 19582 14427
rect 20898 14424 20904 14476
rect 20956 14473 20962 14476
rect 22002 14473 22008 14476
rect 20956 14467 20994 14473
rect 20982 14433 20994 14467
rect 20956 14427 20994 14433
rect 21980 14467 22008 14473
rect 21980 14433 21992 14467
rect 21980 14427 22008 14433
rect 20956 14424 20962 14427
rect 22002 14424 22008 14427
rect 22060 14424 22066 14476
rect 23934 14424 23940 14476
rect 23992 14473 23998 14476
rect 23992 14467 24030 14473
rect 24018 14433 24030 14467
rect 23992 14427 24030 14433
rect 23992 14424 23998 14427
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 24984 14467 25042 14473
rect 24984 14464 24996 14467
rect 24912 14436 24996 14464
rect 24912 14424 24918 14436
rect 24984 14433 24996 14436
rect 25030 14433 25042 14467
rect 24984 14427 25042 14433
rect 2314 14356 2320 14408
rect 2372 14356 2378 14408
rect 4154 14396 4160 14408
rect 4115 14368 4160 14396
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14396 6055 14399
rect 6638 14396 6644 14408
rect 6043 14368 6644 14396
rect 6043 14365 6055 14368
rect 5997 14359 6055 14365
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 9306 14396 9312 14408
rect 8803 14368 9312 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 16850 14396 16856 14408
rect 16439 14368 16856 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17034 14396 17040 14408
rect 16995 14368 17040 14396
rect 17034 14356 17040 14368
rect 17092 14356 17098 14408
rect 22186 14356 22192 14408
rect 22244 14396 22250 14408
rect 22925 14399 22983 14405
rect 22925 14396 22937 14399
rect 22244 14368 22937 14396
rect 22244 14356 22250 14368
rect 22925 14365 22937 14368
rect 22971 14365 22983 14399
rect 22925 14359 22983 14365
rect 10134 14288 10140 14340
rect 10192 14328 10198 14340
rect 10873 14331 10931 14337
rect 10873 14328 10885 14331
rect 10192 14300 10885 14328
rect 10192 14288 10198 14300
rect 10873 14297 10885 14300
rect 10919 14297 10931 14331
rect 10873 14291 10931 14297
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 5169 14263 5227 14269
rect 5169 14260 5181 14263
rect 5132 14232 5181 14260
rect 5132 14220 5138 14232
rect 5169 14229 5181 14232
rect 5215 14229 5227 14263
rect 5169 14223 5227 14229
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 10686 14260 10692 14272
rect 10643 14232 10692 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11238 14260 11244 14272
rect 11199 14232 11244 14260
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 12710 14260 12716 14272
rect 12671 14232 12716 14260
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 12986 14260 12992 14272
rect 12947 14232 12992 14260
rect 12986 14220 12992 14232
rect 13044 14220 13050 14272
rect 19659 14263 19717 14269
rect 19659 14229 19671 14263
rect 19705 14260 19717 14263
rect 20714 14260 20720 14272
rect 19705 14232 20720 14260
rect 19705 14229 19717 14232
rect 19659 14223 19717 14229
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 21039 14263 21097 14269
rect 21039 14229 21051 14263
rect 21085 14260 21097 14263
rect 21542 14260 21548 14272
rect 21085 14232 21548 14260
rect 21085 14229 21097 14232
rect 21039 14223 21097 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22002 14220 22008 14272
rect 22060 14269 22066 14272
rect 22060 14263 22109 14269
rect 22060 14229 22063 14263
rect 22097 14260 22109 14263
rect 22097 14232 22153 14260
rect 22097 14229 22109 14232
rect 22060 14223 22109 14229
rect 22060 14220 22066 14223
rect 23198 14220 23204 14272
rect 23256 14260 23262 14272
rect 24075 14263 24133 14269
rect 24075 14260 24087 14263
rect 23256 14232 24087 14260
rect 23256 14220 23262 14232
rect 24075 14229 24087 14232
rect 24121 14229 24133 14263
rect 24075 14223 24133 14229
rect 25087 14263 25145 14269
rect 25087 14229 25099 14263
rect 25133 14260 25145 14263
rect 25314 14260 25320 14272
rect 25133 14232 25320 14260
rect 25133 14229 25145 14232
rect 25087 14223 25145 14229
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14056 3019 14059
rect 3234 14056 3240 14068
rect 3007 14028 3240 14056
rect 3007 14025 3019 14028
rect 2961 14019 3019 14025
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 4617 14059 4675 14065
rect 4617 14056 4629 14059
rect 4304 14028 4629 14056
rect 4304 14016 4310 14028
rect 4617 14025 4629 14028
rect 4663 14025 4675 14059
rect 4617 14019 4675 14025
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7745 14059 7803 14065
rect 7745 14056 7757 14059
rect 7064 14028 7757 14056
rect 7064 14016 7070 14028
rect 7745 14025 7757 14028
rect 7791 14025 7803 14059
rect 7745 14019 7803 14025
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8294 14056 8300 14068
rect 8159 14028 8300 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8478 14056 8484 14068
rect 8439 14028 8484 14056
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 8711 14059 8769 14065
rect 8711 14025 8723 14059
rect 8757 14056 8769 14059
rect 11238 14056 11244 14068
rect 8757 14028 11244 14056
rect 8757 14025 8769 14028
rect 8711 14019 8769 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 11480 14028 11805 14056
rect 11480 14016 11486 14028
rect 11793 14025 11805 14028
rect 11839 14025 11851 14059
rect 11793 14019 11851 14025
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 12768 14028 13369 14056
rect 12768 14016 12774 14028
rect 13357 14025 13369 14028
rect 13403 14025 13415 14059
rect 13357 14019 13415 14025
rect 15381 14059 15439 14065
rect 15381 14025 15393 14059
rect 15427 14056 15439 14059
rect 15470 14056 15476 14068
rect 15427 14028 15476 14056
rect 15427 14025 15439 14028
rect 15381 14019 15439 14025
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 16393 14059 16451 14065
rect 16393 14025 16405 14059
rect 16439 14056 16451 14059
rect 16482 14056 16488 14068
rect 16439 14028 16488 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 16482 14016 16488 14028
rect 16540 14056 16546 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16540 14028 16681 14056
rect 16540 14016 16546 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 16669 14019 16727 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 19610 14016 19616 14068
rect 19668 14056 19674 14068
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 19668 14028 20085 14056
rect 19668 14016 19674 14028
rect 20073 14025 20085 14028
rect 20119 14025 20131 14059
rect 20073 14019 20131 14025
rect 20898 14016 20904 14068
rect 20956 14056 20962 14068
rect 21358 14056 21364 14068
rect 20956 14028 21364 14056
rect 20956 14016 20962 14028
rect 21358 14016 21364 14028
rect 21416 14056 21422 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21416 14028 21465 14056
rect 21416 14016 21422 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 21910 14016 21916 14068
rect 21968 14056 21974 14068
rect 22097 14059 22155 14065
rect 22097 14056 22109 14059
rect 21968 14028 22109 14056
rect 21968 14016 21974 14028
rect 22097 14025 22109 14028
rect 22143 14025 22155 14059
rect 22097 14019 22155 14025
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25409 14059 25467 14065
rect 25409 14056 25421 14059
rect 24912 14028 25421 14056
rect 24912 14016 24918 14028
rect 25409 14025 25421 14028
rect 25455 14025 25467 14059
rect 25409 14019 25467 14025
rect 1854 13948 1860 14000
rect 1912 13988 1918 14000
rect 3605 13991 3663 13997
rect 3605 13988 3617 13991
rect 1912 13960 3617 13988
rect 1912 13948 1918 13960
rect 3605 13957 3617 13960
rect 3651 13957 3663 13991
rect 10594 13988 10600 14000
rect 10555 13960 10600 13988
rect 3605 13951 3663 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 10870 13988 10876 14000
rect 10831 13960 10876 13988
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 13262 13948 13268 14000
rect 13320 13988 13326 14000
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 13320 13960 14013 13988
rect 13320 13948 13326 13960
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 17129 13991 17187 13997
rect 17129 13988 17141 13991
rect 16632 13960 17141 13988
rect 16632 13948 16638 13960
rect 17129 13957 17141 13960
rect 17175 13988 17187 13991
rect 18138 13988 18144 14000
rect 17175 13960 18144 13988
rect 17175 13957 17187 13960
rect 17129 13951 17187 13957
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 19518 13948 19524 14000
rect 19576 13988 19582 14000
rect 19797 13991 19855 13997
rect 19797 13988 19809 13991
rect 19576 13960 19809 13988
rect 19576 13948 19582 13960
rect 19797 13957 19809 13960
rect 19843 13957 19855 13991
rect 19797 13951 19855 13957
rect 24210 13948 24216 14000
rect 24268 13988 24274 14000
rect 25041 13991 25099 13997
rect 25041 13988 25053 13991
rect 24268 13960 25053 13988
rect 24268 13948 24274 13960
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2222 13920 2228 13932
rect 2087 13892 2228 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 3927 13923 3985 13929
rect 3927 13889 3939 13923
rect 3973 13920 3985 13923
rect 4062 13920 4068 13932
rect 3973 13892 4068 13920
rect 3973 13889 3985 13892
rect 3927 13883 3985 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 5074 13920 5080 13932
rect 4356 13892 5080 13920
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 3824 13855 3882 13861
rect 3824 13852 3836 13855
rect 3016 13824 3836 13852
rect 3016 13812 3022 13824
rect 3824 13821 3836 13824
rect 3870 13852 3882 13855
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 3870 13824 4261 13852
rect 3870 13821 3882 13824
rect 3824 13815 3882 13821
rect 4249 13821 4261 13824
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 1394 13744 1400 13796
rect 1452 13784 1458 13796
rect 1854 13784 1860 13796
rect 1452 13756 1860 13784
rect 1452 13744 1458 13756
rect 1854 13744 1860 13756
rect 1912 13744 1918 13796
rect 2314 13784 2320 13796
rect 2056 13756 2320 13784
rect 2056 13728 2084 13756
rect 2314 13744 2320 13756
rect 2372 13793 2378 13796
rect 2372 13787 2420 13793
rect 2372 13753 2374 13787
rect 2408 13784 2420 13787
rect 3237 13787 3295 13793
rect 3237 13784 3249 13787
rect 2408 13756 3249 13784
rect 2408 13753 2420 13756
rect 2372 13747 2420 13753
rect 3237 13753 3249 13756
rect 3283 13753 3295 13787
rect 4356 13784 4384 13892
rect 5074 13880 5080 13892
rect 5132 13920 5138 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5132 13892 5273 13920
rect 5132 13880 5138 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5905 13923 5963 13929
rect 5905 13920 5917 13923
rect 5500 13892 5917 13920
rect 5500 13880 5506 13892
rect 5905 13889 5917 13892
rect 5951 13920 5963 13923
rect 7190 13920 7196 13932
rect 5951 13892 7196 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 7190 13880 7196 13892
rect 7248 13880 7254 13932
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9766 13920 9772 13932
rect 9723 13892 9772 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 12986 13920 12992 13932
rect 12492 13892 12992 13920
rect 12492 13880 12498 13892
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15470 13920 15476 13932
rect 15059 13892 15476 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 23750 13880 23756 13932
rect 23808 13920 23814 13932
rect 24719 13923 24777 13929
rect 24719 13920 24731 13923
rect 23808 13892 24731 13920
rect 23808 13880 23814 13892
rect 24719 13889 24731 13892
rect 24765 13889 24777 13923
rect 24719 13883 24777 13889
rect 6822 13861 6828 13864
rect 6821 13852 6828 13861
rect 6783 13824 6828 13852
rect 6821 13815 6828 13824
rect 6822 13812 6828 13815
rect 6880 13812 6886 13864
rect 8570 13812 8576 13864
rect 8628 13861 8634 13864
rect 8628 13855 8666 13861
rect 8654 13852 8666 13855
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8654 13824 9045 13852
rect 8654 13821 8666 13824
rect 8628 13815 8666 13821
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 15378 13852 15384 13864
rect 9033 13815 9091 13821
rect 15120 13824 15384 13852
rect 8628 13812 8634 13815
rect 3237 13747 3295 13753
rect 4080 13756 4384 13784
rect 5353 13787 5411 13793
rect 2372 13744 2378 13747
rect 4080 13728 4108 13756
rect 5353 13753 5365 13787
rect 5399 13784 5411 13787
rect 5534 13784 5540 13796
rect 5399 13756 5540 13784
rect 5399 13753 5411 13756
rect 5353 13747 5411 13753
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2038 13716 2044 13728
rect 1995 13688 2044 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 4062 13676 4068 13728
rect 4120 13676 4126 13728
rect 5077 13719 5135 13725
rect 5077 13685 5089 13719
rect 5123 13716 5135 13719
rect 5368 13716 5396 13747
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 6270 13784 6276 13796
rect 6183 13756 6276 13784
rect 6270 13744 6276 13756
rect 6328 13784 6334 13796
rect 6641 13787 6699 13793
rect 6641 13784 6653 13787
rect 6328 13756 6653 13784
rect 6328 13744 6334 13756
rect 6641 13753 6653 13756
rect 6687 13784 6699 13787
rect 7187 13787 7245 13793
rect 7187 13784 7199 13787
rect 6687 13756 7199 13784
rect 6687 13753 6699 13756
rect 6641 13747 6699 13753
rect 7187 13753 7199 13756
rect 7233 13784 7245 13787
rect 9585 13787 9643 13793
rect 9585 13784 9597 13787
rect 7233 13756 9597 13784
rect 7233 13753 7245 13756
rect 7187 13747 7245 13753
rect 9585 13753 9597 13756
rect 9631 13784 9643 13787
rect 10039 13787 10097 13793
rect 10039 13784 10051 13787
rect 9631 13756 10051 13784
rect 9631 13753 9643 13756
rect 9585 13747 9643 13753
rect 10039 13753 10051 13756
rect 10085 13784 10097 13787
rect 10226 13784 10232 13796
rect 10085 13756 10232 13784
rect 10085 13753 10097 13756
rect 10039 13747 10097 13753
rect 10226 13744 10232 13756
rect 10284 13784 10290 13796
rect 12758 13787 12816 13793
rect 12758 13784 12770 13787
rect 10284 13756 11468 13784
rect 10284 13744 10290 13756
rect 11440 13728 11468 13756
rect 12176 13756 12770 13784
rect 11422 13716 11428 13728
rect 5123 13688 5396 13716
rect 11383 13688 11428 13716
rect 5123 13685 5135 13688
rect 5077 13679 5135 13685
rect 11422 13676 11428 13688
rect 11480 13716 11486 13728
rect 12176 13725 12204 13756
rect 12758 13753 12770 13756
rect 12804 13784 12816 13787
rect 13538 13784 13544 13796
rect 12804 13756 13544 13784
rect 12804 13753 12816 13756
rect 12758 13747 12816 13753
rect 13538 13744 13544 13756
rect 13596 13784 13602 13796
rect 13633 13787 13691 13793
rect 13633 13784 13645 13787
rect 13596 13756 13645 13784
rect 13596 13744 13602 13756
rect 13633 13753 13645 13756
rect 13679 13753 13691 13787
rect 13633 13747 13691 13753
rect 14185 13787 14243 13793
rect 14185 13753 14197 13787
rect 14231 13784 14243 13787
rect 15120 13784 15148 13824
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 16390 13852 16396 13864
rect 15988 13824 16396 13852
rect 15988 13812 15994 13824
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 17218 13812 17224 13864
rect 17276 13852 17282 13864
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17276 13824 17785 13852
rect 17276 13812 17282 13824
rect 17773 13821 17785 13824
rect 17819 13852 17831 13855
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 17819 13824 18153 13852
rect 17819 13821 17831 13824
rect 17773 13815 17831 13821
rect 18141 13821 18153 13824
rect 18187 13821 18199 13855
rect 18141 13815 18199 13821
rect 18690 13812 18696 13864
rect 18748 13852 18754 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 18748 13824 18797 13852
rect 18748 13812 18754 13824
rect 18785 13821 18797 13824
rect 18831 13852 18843 13855
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 18831 13824 19625 13852
rect 18831 13821 18843 13824
rect 18785 13815 18843 13821
rect 19613 13821 19625 13824
rect 19659 13852 19671 13855
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 19659 13824 20453 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20441 13821 20453 13824
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 20676 13855 20734 13861
rect 20676 13821 20688 13855
rect 20722 13821 20734 13855
rect 20676 13815 20734 13821
rect 20763 13855 20821 13861
rect 20763 13821 20775 13855
rect 20809 13852 20821 13855
rect 21174 13852 21180 13864
rect 20809 13824 21180 13852
rect 20809 13821 20821 13824
rect 20763 13815 20821 13821
rect 15794 13787 15852 13793
rect 15794 13784 15806 13787
rect 14231 13756 15148 13784
rect 15396 13756 15806 13784
rect 14231 13753 14243 13756
rect 14185 13747 14243 13753
rect 15396 13728 15424 13756
rect 15794 13753 15806 13756
rect 15840 13753 15852 13787
rect 15794 13747 15852 13753
rect 19978 13744 19984 13796
rect 20036 13784 20042 13796
rect 20686 13784 20714 13815
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 21704 13855 21762 13861
rect 21704 13821 21716 13855
rect 21750 13852 21762 13855
rect 22557 13855 22615 13861
rect 22557 13852 22569 13855
rect 21750 13824 22569 13852
rect 21750 13821 21762 13824
rect 21704 13815 21762 13821
rect 22557 13821 22569 13824
rect 22603 13852 22615 13855
rect 23106 13852 23112 13864
rect 22603 13824 23112 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 23106 13812 23112 13824
rect 23164 13812 23170 13864
rect 23934 13852 23940 13864
rect 23895 13824 23940 13852
rect 23934 13812 23940 13824
rect 23992 13812 23998 13864
rect 24632 13855 24690 13861
rect 24632 13821 24644 13855
rect 24678 13852 24690 13855
rect 24826 13852 24854 13960
rect 25041 13957 25053 13960
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 24678 13824 24854 13852
rect 24678 13821 24690 13824
rect 24632 13815 24690 13821
rect 20036 13756 20944 13784
rect 20036 13744 20042 13756
rect 20916 13728 20944 13756
rect 12161 13719 12219 13725
rect 12161 13716 12173 13719
rect 11480 13688 12173 13716
rect 11480 13676 11486 13688
rect 12161 13685 12173 13688
rect 12207 13685 12219 13719
rect 12161 13679 12219 13685
rect 15378 13676 15384 13728
rect 15436 13676 15442 13728
rect 20898 13676 20904 13728
rect 20956 13716 20962 13728
rect 21085 13719 21143 13725
rect 21085 13716 21097 13719
rect 20956 13688 21097 13716
rect 20956 13676 20962 13688
rect 21085 13685 21097 13688
rect 21131 13685 21143 13719
rect 21085 13679 21143 13685
rect 21775 13719 21833 13725
rect 21775 13685 21787 13719
rect 21821 13716 21833 13719
rect 22554 13716 22560 13728
rect 21821 13688 22560 13716
rect 21821 13685 21833 13688
rect 21775 13679 21833 13685
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 25590 13716 25596 13728
rect 25551 13688 25596 13716
rect 25590 13676 25596 13688
rect 25648 13676 25654 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2832 13484 3065 13512
rect 2832 13472 2838 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3053 13475 3111 13481
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 4212 13484 4537 13512
rect 4212 13472 4218 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 4525 13475 4583 13481
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 5258 13512 5264 13524
rect 5123 13484 5264 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 5592 13484 6377 13512
rect 5592 13472 5598 13484
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 6638 13512 6644 13524
rect 6599 13484 6644 13512
rect 6365 13475 6423 13481
rect 6638 13472 6644 13484
rect 6696 13512 6702 13524
rect 7285 13515 7343 13521
rect 7285 13512 7297 13515
rect 6696 13484 7297 13512
rect 6696 13472 6702 13484
rect 7285 13481 7297 13484
rect 7331 13481 7343 13515
rect 7285 13475 7343 13481
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 9582 13512 9588 13524
rect 9539 13484 9588 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16908 13484 16957 13512
rect 16908 13472 16914 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 17310 13512 17316 13524
rect 17271 13484 17316 13512
rect 16945 13475 17003 13481
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 18601 13515 18659 13521
rect 18601 13481 18613 13515
rect 18647 13512 18659 13515
rect 18690 13512 18696 13524
rect 18647 13484 18696 13512
rect 18647 13481 18659 13484
rect 18601 13475 18659 13481
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 19199 13515 19257 13521
rect 19199 13512 19211 13515
rect 18932 13484 19211 13512
rect 18932 13472 18938 13484
rect 19199 13481 19211 13484
rect 19245 13481 19257 13515
rect 19199 13475 19257 13481
rect 2038 13404 2044 13456
rect 2096 13444 2102 13456
rect 2454 13447 2512 13453
rect 2454 13444 2466 13447
rect 2096 13416 2466 13444
rect 2096 13404 2102 13416
rect 2454 13413 2466 13416
rect 2500 13413 2512 13447
rect 2454 13407 2512 13413
rect 5442 13404 5448 13456
rect 5500 13404 5506 13456
rect 5807 13447 5865 13453
rect 5807 13413 5819 13447
rect 5853 13444 5865 13447
rect 6270 13444 6276 13456
rect 5853 13416 6276 13444
rect 5853 13413 5865 13416
rect 5807 13407 5865 13413
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 8294 13444 8300 13456
rect 7484 13416 8300 13444
rect 3878 13336 3884 13388
rect 3936 13376 3942 13388
rect 4132 13379 4190 13385
rect 4132 13376 4144 13379
rect 3936 13348 4144 13376
rect 3936 13336 3942 13348
rect 4132 13345 4144 13348
rect 4178 13376 4190 13379
rect 4706 13376 4712 13388
rect 4178 13348 4712 13376
rect 4178 13345 4190 13348
rect 4132 13339 4190 13345
rect 4706 13336 4712 13348
rect 4764 13376 4770 13388
rect 5460 13376 5488 13404
rect 7484 13385 7512 13416
rect 8294 13404 8300 13416
rect 8352 13404 8358 13456
rect 9674 13404 9680 13456
rect 9732 13444 9738 13456
rect 10042 13444 10048 13456
rect 9732 13416 10048 13444
rect 9732 13404 9738 13416
rect 10042 13404 10048 13416
rect 10100 13404 10106 13456
rect 10226 13444 10232 13456
rect 10187 13416 10232 13444
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 10321 13447 10379 13453
rect 10321 13413 10333 13447
rect 10367 13444 10379 13447
rect 10686 13444 10692 13456
rect 10367 13416 10692 13444
rect 10367 13413 10379 13416
rect 10321 13407 10379 13413
rect 10686 13404 10692 13416
rect 10744 13444 10750 13456
rect 10870 13444 10876 13456
rect 10744 13416 10876 13444
rect 10744 13404 10750 13416
rect 10870 13404 10876 13416
rect 10928 13404 10934 13456
rect 13814 13444 13820 13456
rect 13775 13416 13820 13444
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 15470 13444 15476 13456
rect 14384 13416 15476 13444
rect 4764 13348 5488 13376
rect 7469 13379 7527 13385
rect 4764 13336 4770 13348
rect 7469 13345 7481 13379
rect 7515 13345 7527 13379
rect 7650 13376 7656 13388
rect 7611 13348 7656 13376
rect 7469 13339 7527 13345
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 12526 13376 12532 13388
rect 12487 13348 12532 13376
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 2682 13308 2688 13320
rect 2179 13280 2688 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 5534 13308 5540 13320
rect 5491 13280 5540 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13308 10931 13311
rect 11054 13308 11060 13320
rect 10919 13280 11060 13308
rect 10919 13277 10931 13280
rect 10873 13271 10931 13277
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 13262 13308 13268 13320
rect 12851 13280 13268 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13722 13308 13728 13320
rect 13683 13280 13728 13308
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14001 13311 14059 13317
rect 14001 13308 14013 13311
rect 13964 13280 14013 13308
rect 13964 13268 13970 13280
rect 14001 13277 14013 13280
rect 14047 13277 14059 13311
rect 14001 13271 14059 13277
rect 4203 13243 4261 13249
rect 4203 13209 4215 13243
rect 4249 13240 4261 13243
rect 4614 13240 4620 13252
rect 4249 13212 4620 13240
rect 4249 13209 4261 13212
rect 4203 13203 4261 13209
rect 4614 13200 4620 13212
rect 4672 13200 4678 13252
rect 14384 13240 14412 13416
rect 15470 13404 15476 13416
rect 15528 13444 15534 13456
rect 16117 13447 16175 13453
rect 16117 13444 16129 13447
rect 15528 13416 16129 13444
rect 15528 13404 15534 13416
rect 16117 13413 16129 13416
rect 16163 13444 16175 13447
rect 16758 13444 16764 13456
rect 16163 13416 16764 13444
rect 16163 13413 16175 13416
rect 16117 13407 16175 13413
rect 16758 13404 16764 13416
rect 16816 13404 16822 13456
rect 17678 13444 17684 13456
rect 17639 13416 17684 13444
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 19150 13385 19156 13388
rect 19128 13379 19156 13385
rect 19128 13345 19140 13379
rect 19128 13339 19156 13345
rect 19150 13336 19156 13339
rect 19208 13336 19214 13388
rect 20990 13385 20996 13388
rect 20968 13379 20996 13385
rect 20968 13345 20980 13379
rect 20968 13339 20996 13345
rect 20990 13336 20996 13339
rect 21048 13336 21054 13388
rect 22624 13379 22682 13385
rect 22624 13345 22636 13379
rect 22670 13376 22682 13379
rect 23382 13376 23388 13388
rect 22670 13348 23388 13376
rect 22670 13345 22682 13348
rect 22624 13339 22682 13345
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 23566 13336 23572 13388
rect 23624 13385 23630 13388
rect 23624 13379 23662 13385
rect 23650 13345 23662 13379
rect 23624 13339 23662 13345
rect 23624 13336 23630 13339
rect 24026 13336 24032 13388
rect 24084 13376 24090 13388
rect 24616 13379 24674 13385
rect 24616 13376 24628 13379
rect 24084 13348 24628 13376
rect 24084 13336 24090 13348
rect 24616 13345 24628 13348
rect 24662 13376 24674 13379
rect 25130 13376 25136 13388
rect 24662 13348 25136 13376
rect 24662 13345 24674 13348
rect 24616 13339 24674 13345
rect 25130 13336 25136 13348
rect 25188 13336 25194 13388
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17368 13280 17601 13308
rect 17368 13268 17374 13280
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 18230 13308 18236 13320
rect 18191 13280 18236 13308
rect 17589 13271 17647 13277
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 11072 13212 14412 13240
rect 11072 13184 11100 13212
rect 23474 13200 23480 13252
rect 23532 13240 23538 13252
rect 24719 13243 24777 13249
rect 24719 13240 24731 13243
rect 23532 13212 24731 13240
rect 23532 13200 23538 13212
rect 24719 13209 24731 13212
rect 24765 13209 24777 13243
rect 24719 13203 24777 13209
rect 1765 13175 1823 13181
rect 1765 13141 1777 13175
rect 1811 13172 1823 13175
rect 1854 13172 1860 13184
rect 1811 13144 1860 13172
rect 1811 13141 1823 13144
rect 1765 13135 1823 13141
rect 1854 13132 1860 13144
rect 1912 13172 1918 13184
rect 2222 13172 2228 13184
rect 1912 13144 2228 13172
rect 1912 13132 1918 13144
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 4982 13132 4988 13184
rect 5040 13172 5046 13184
rect 5442 13172 5448 13184
rect 5040 13144 5448 13172
rect 5040 13132 5046 13144
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 7098 13172 7104 13184
rect 6880 13144 7104 13172
rect 6880 13132 6886 13144
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 9861 13175 9919 13181
rect 9861 13172 9873 13175
rect 9824 13144 9873 13172
rect 9824 13132 9830 13144
rect 9861 13141 9873 13144
rect 9907 13141 9919 13175
rect 9861 13135 9919 13141
rect 11054 13132 11060 13184
rect 11112 13132 11118 13184
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 21082 13181 21088 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 15436 13144 15485 13172
rect 15436 13132 15442 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 21039 13175 21088 13181
rect 21039 13141 21051 13175
rect 21085 13141 21088 13175
rect 21039 13135 21088 13141
rect 21082 13132 21088 13135
rect 21140 13132 21146 13184
rect 22695 13175 22753 13181
rect 22695 13141 22707 13175
rect 22741 13172 22753 13175
rect 22830 13172 22836 13184
rect 22741 13144 22836 13172
rect 22741 13141 22753 13144
rect 22695 13135 22753 13141
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 23707 13175 23765 13181
rect 23707 13141 23719 13175
rect 23753 13172 23765 13175
rect 24210 13172 24216 13184
rect 23753 13144 24216 13172
rect 23753 13141 23765 13144
rect 23707 13135 23765 13141
rect 24210 13132 24216 13144
rect 24268 13132 24274 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3237 12971 3295 12977
rect 3237 12968 3249 12971
rect 2832 12940 3249 12968
rect 2832 12928 2838 12940
rect 3237 12937 3249 12940
rect 3283 12937 3295 12971
rect 3237 12931 3295 12937
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 4706 12968 4712 12980
rect 4571 12940 4712 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 1854 12764 1860 12776
rect 1815 12736 1860 12764
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 2222 12764 2228 12776
rect 2183 12736 2228 12764
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2409 12767 2467 12773
rect 2409 12733 2421 12767
rect 2455 12764 2467 12767
rect 2682 12764 2688 12776
rect 2455 12736 2688 12764
rect 2455 12733 2467 12736
rect 2409 12727 2467 12733
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 3252 12696 3280 12931
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 6089 12971 6147 12977
rect 6089 12937 6101 12971
rect 6135 12968 6147 12971
rect 6270 12968 6276 12980
rect 6135 12940 6276 12968
rect 6135 12937 6147 12940
rect 6089 12931 6147 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 7653 12971 7711 12977
rect 7653 12937 7665 12971
rect 7699 12968 7711 12971
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7699 12940 7941 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 7929 12937 7941 12940
rect 7975 12968 7987 12971
rect 8294 12968 8300 12980
rect 7975 12940 8300 12968
rect 7975 12937 7987 12940
rect 7929 12931 7987 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8895 12971 8953 12977
rect 8895 12937 8907 12971
rect 8941 12968 8953 12971
rect 10134 12968 10140 12980
rect 8941 12940 10140 12968
rect 8941 12937 8953 12940
rect 8895 12931 8953 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 13538 12928 13544 12980
rect 13596 12968 13602 12980
rect 13725 12971 13783 12977
rect 13725 12968 13737 12971
rect 13596 12940 13737 12968
rect 13596 12928 13602 12940
rect 13725 12937 13737 12940
rect 13771 12968 13783 12971
rect 13814 12968 13820 12980
rect 13771 12940 13820 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 15289 12971 15347 12977
rect 15289 12937 15301 12971
rect 15335 12968 15347 12971
rect 16022 12968 16028 12980
rect 15335 12940 16028 12968
rect 15335 12937 15347 12940
rect 15289 12931 15347 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16758 12968 16764 12980
rect 16719 12940 16764 12968
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 17552 12940 17601 12968
rect 17552 12928 17558 12940
rect 17589 12937 17601 12940
rect 17635 12968 17647 12971
rect 17678 12968 17684 12980
rect 17635 12940 17684 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 20165 12971 20223 12977
rect 20165 12937 20177 12971
rect 20211 12968 20223 12971
rect 20622 12968 20628 12980
rect 20211 12940 20628 12968
rect 20211 12937 20223 12940
rect 20165 12931 20223 12937
rect 4062 12900 4068 12912
rect 4023 12872 4068 12900
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 10870 12900 10876 12912
rect 10831 12872 10876 12900
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 18046 12860 18052 12912
rect 18104 12860 18110 12912
rect 3510 12832 3516 12844
rect 3471 12804 3516 12832
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12832 5135 12835
rect 5258 12832 5264 12844
rect 5123 12804 5264 12832
rect 5123 12801 5135 12804
rect 5077 12795 5135 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 7156 12804 7297 12832
rect 7156 12792 7162 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 8018 12832 8024 12844
rect 7800 12804 8024 12832
rect 7800 12792 7806 12804
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 11471 12835 11529 12841
rect 11471 12801 11483 12835
rect 11517 12832 11529 12835
rect 12342 12832 12348 12844
rect 11517 12804 12348 12832
rect 11517 12801 11529 12804
rect 11471 12795 11529 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 14550 12832 14556 12844
rect 14511 12804 14556 12832
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16022 12832 16028 12844
rect 15887 12804 16028 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16298 12832 16304 12844
rect 16259 12804 16304 12832
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 18064 12832 18092 12860
rect 18509 12835 18567 12841
rect 18509 12832 18521 12835
rect 18064 12804 18521 12832
rect 18509 12801 18521 12804
rect 18555 12801 18567 12835
rect 18509 12795 18567 12801
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 7006 12764 7012 12776
rect 6687 12736 7012 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12764 7435 12767
rect 7650 12764 7656 12776
rect 7423 12736 7656 12764
rect 7423 12733 7435 12736
rect 7377 12727 7435 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 8754 12724 8760 12776
rect 8812 12773 8818 12776
rect 8812 12767 8850 12773
rect 8838 12764 8850 12767
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8838 12736 9229 12764
rect 8838 12733 8850 12736
rect 8812 12727 8850 12733
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 8812 12724 8818 12727
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11368 12767 11426 12773
rect 11368 12764 11380 12767
rect 11204 12736 11380 12764
rect 11204 12724 11210 12736
rect 11368 12733 11380 12736
rect 11414 12733 11426 12767
rect 11368 12727 11426 12733
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12764 12498 12776
rect 12529 12767 12587 12773
rect 12529 12764 12541 12767
rect 12492 12736 12541 12764
rect 12492 12724 12498 12736
rect 12529 12733 12541 12736
rect 12575 12733 12587 12767
rect 17221 12767 17279 12773
rect 12529 12727 12587 12733
rect 13096 12736 13952 12764
rect 3605 12699 3663 12705
rect 3605 12696 3617 12699
rect 3252 12668 3617 12696
rect 3605 12665 3617 12668
rect 3651 12665 3663 12699
rect 3605 12659 3663 12665
rect 5169 12699 5227 12705
rect 5169 12665 5181 12699
rect 5215 12665 5227 12699
rect 5718 12696 5724 12708
rect 5679 12668 5724 12696
rect 5169 12659 5227 12665
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2096 12600 2697 12628
rect 2096 12588 2102 12600
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 2685 12591 2743 12597
rect 4798 12588 4804 12640
rect 4856 12628 4862 12640
rect 4893 12631 4951 12637
rect 4893 12628 4905 12631
rect 4856 12600 4905 12628
rect 4856 12588 4862 12600
rect 4893 12597 4905 12600
rect 4939 12628 4951 12631
rect 5184 12628 5212 12659
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 9861 12699 9919 12705
rect 9861 12696 9873 12699
rect 8588 12668 9873 12696
rect 8588 12640 8616 12668
rect 9861 12665 9873 12668
rect 9907 12665 9919 12699
rect 9861 12659 9919 12665
rect 9953 12699 10011 12705
rect 9953 12665 9965 12699
rect 9999 12665 10011 12699
rect 9953 12659 10011 12665
rect 10505 12699 10563 12705
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 10686 12696 10692 12708
rect 10551 12668 10692 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 4939 12600 5212 12628
rect 4939 12597 4951 12600
rect 4893 12591 4951 12597
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 7156 12600 7665 12628
rect 7156 12588 7162 12600
rect 7653 12597 7665 12600
rect 7699 12597 7711 12631
rect 8570 12628 8576 12640
rect 8531 12600 8576 12628
rect 7653 12591 7711 12597
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12628 9735 12631
rect 9968 12628 9996 12659
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 11885 12699 11943 12705
rect 11885 12665 11897 12699
rect 11931 12696 11943 12699
rect 11931 12668 12296 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 11054 12628 11060 12640
rect 9723 12600 11060 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 12268 12628 12296 12668
rect 12342 12656 12348 12708
rect 12400 12696 12406 12708
rect 13096 12696 13124 12736
rect 12400 12668 13124 12696
rect 13173 12699 13231 12705
rect 12400 12656 12406 12668
rect 13173 12665 13185 12699
rect 13219 12696 13231 12699
rect 13630 12696 13636 12708
rect 13219 12668 13636 12696
rect 13219 12665 13231 12668
rect 13173 12659 13231 12665
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 13924 12696 13952 12736
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 17586 12764 17592 12776
rect 17267 12736 17592 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17586 12724 17592 12736
rect 17644 12764 17650 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17644 12736 18061 12764
rect 17644 12724 17650 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 18138 12724 18144 12776
rect 18196 12764 18202 12776
rect 18325 12767 18383 12773
rect 18196 12736 18241 12764
rect 18196 12724 18202 12736
rect 18325 12733 18337 12767
rect 18371 12764 18383 12767
rect 18690 12764 18696 12776
rect 18371 12736 18696 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 14274 12696 14280 12708
rect 13924 12668 14280 12696
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 14366 12656 14372 12708
rect 14424 12696 14430 12708
rect 15933 12699 15991 12705
rect 14424 12668 14469 12696
rect 14424 12656 14430 12668
rect 15933 12665 15945 12699
rect 15979 12665 15991 12699
rect 15933 12659 15991 12665
rect 12526 12628 12532 12640
rect 12268 12600 12532 12628
rect 12526 12588 12532 12600
rect 12584 12628 12590 12640
rect 12710 12628 12716 12640
rect 12584 12600 12716 12628
rect 12584 12588 12590 12600
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 14093 12631 14151 12637
rect 14093 12597 14105 12631
rect 14139 12628 14151 12631
rect 14384 12628 14412 12656
rect 14139 12600 14412 12628
rect 14139 12597 14151 12600
rect 14093 12591 14151 12597
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 15565 12631 15623 12637
rect 15565 12628 15577 12631
rect 15344 12600 15577 12628
rect 15344 12588 15350 12600
rect 15565 12597 15577 12600
rect 15611 12628 15623 12631
rect 15948 12628 15976 12659
rect 15611 12600 15976 12628
rect 15611 12597 15623 12600
rect 15565 12591 15623 12597
rect 18046 12588 18052 12640
rect 18104 12628 18110 12640
rect 18340 12628 18368 12727
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 19680 12767 19738 12773
rect 19680 12733 19692 12767
rect 19726 12764 19738 12767
rect 20180 12764 20208 12931
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 21637 12971 21695 12977
rect 21637 12968 21649 12971
rect 21048 12940 21649 12968
rect 21048 12928 21054 12940
rect 21637 12937 21649 12940
rect 21683 12937 21695 12971
rect 23382 12968 23388 12980
rect 23343 12940 23388 12968
rect 21637 12931 21695 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23624 12940 23857 12968
rect 23624 12928 23630 12940
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 24210 12928 24216 12980
rect 24268 12968 24274 12980
rect 24397 12971 24455 12977
rect 24397 12968 24409 12971
rect 24268 12940 24409 12968
rect 24268 12928 24274 12940
rect 24397 12937 24409 12940
rect 24443 12937 24455 12971
rect 25130 12968 25136 12980
rect 25091 12940 25136 12968
rect 24397 12931 24455 12937
rect 19726 12736 20208 12764
rect 19726 12733 19738 12736
rect 19680 12727 19738 12733
rect 20806 12724 20812 12776
rect 20864 12773 20870 12776
rect 22646 12773 22652 12776
rect 20864 12767 20902 12773
rect 20890 12764 20902 12767
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 20890 12736 21281 12764
rect 20890 12733 20902 12736
rect 20864 12727 20902 12733
rect 21269 12733 21281 12736
rect 21315 12733 21327 12767
rect 22624 12767 22652 12773
rect 22624 12764 22636 12767
rect 22559 12736 22636 12764
rect 21269 12727 21327 12733
rect 22624 12733 22636 12736
rect 22704 12764 22710 12776
rect 24412 12764 24440 12931
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 22704 12736 23152 12764
rect 24412 12736 24593 12764
rect 22624 12727 22652 12733
rect 20864 12724 20870 12727
rect 22646 12724 22652 12727
rect 22704 12724 22710 12736
rect 23124 12705 23152 12736
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 23109 12699 23167 12705
rect 23109 12665 23121 12699
rect 23155 12696 23167 12699
rect 25038 12696 25044 12708
rect 23155 12668 25044 12696
rect 23155 12665 23167 12668
rect 23109 12659 23167 12665
rect 25038 12656 25044 12668
rect 25096 12656 25102 12708
rect 18104 12600 18368 12628
rect 18104 12588 18110 12600
rect 18414 12588 18420 12640
rect 18472 12628 18478 12640
rect 18690 12628 18696 12640
rect 18472 12600 18696 12628
rect 18472 12588 18478 12600
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 19150 12628 19156 12640
rect 19111 12600 19156 12628
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20990 12637 20996 12640
rect 19751 12631 19809 12637
rect 19751 12628 19763 12631
rect 19392 12600 19763 12628
rect 19392 12588 19398 12600
rect 19751 12597 19763 12600
rect 19797 12597 19809 12631
rect 19751 12591 19809 12597
rect 20947 12631 20996 12637
rect 20947 12597 20959 12631
rect 20993 12597 20996 12631
rect 20947 12591 20996 12597
rect 20990 12588 20996 12591
rect 21048 12588 21054 12640
rect 22695 12631 22753 12637
rect 22695 12597 22707 12631
rect 22741 12628 22753 12631
rect 23382 12628 23388 12640
rect 22741 12600 23388 12628
rect 22741 12597 22753 12600
rect 22695 12591 22753 12597
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 24765 12631 24823 12637
rect 24765 12597 24777 12631
rect 24811 12628 24823 12631
rect 25130 12628 25136 12640
rect 24811 12600 25136 12628
rect 24811 12597 24823 12600
rect 24765 12591 24823 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3053 12427 3111 12433
rect 3053 12424 3065 12427
rect 2832 12396 3065 12424
rect 2832 12384 2838 12396
rect 3053 12393 3065 12396
rect 3099 12393 3111 12427
rect 3510 12424 3516 12436
rect 3471 12396 3516 12424
rect 3053 12387 3111 12393
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 5350 12424 5356 12436
rect 5040 12396 5356 12424
rect 5040 12384 5046 12396
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 5534 12424 5540 12436
rect 5447 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12424 5598 12436
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 5592 12396 5733 12424
rect 5592 12384 5598 12396
rect 5721 12393 5733 12396
rect 5767 12393 5779 12427
rect 5721 12387 5779 12393
rect 7834 12384 7840 12436
rect 7892 12384 7898 12436
rect 9490 12424 9496 12436
rect 9451 12396 9496 12424
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 9766 12384 9772 12436
rect 9824 12384 9830 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 10597 12427 10655 12433
rect 9916 12396 10548 12424
rect 9916 12384 9922 12396
rect 1578 12316 1584 12368
rect 1636 12356 1642 12368
rect 2133 12359 2191 12365
rect 2133 12356 2145 12359
rect 1636 12328 2145 12356
rect 1636 12316 1642 12328
rect 2133 12325 2145 12328
rect 2179 12325 2191 12359
rect 2133 12319 2191 12325
rect 2225 12359 2283 12365
rect 2225 12325 2237 12359
rect 2271 12356 2283 12359
rect 2314 12356 2320 12368
rect 2271 12328 2320 12356
rect 2271 12325 2283 12328
rect 2225 12319 2283 12325
rect 2314 12316 2320 12328
rect 2372 12316 2378 12368
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 4249 12359 4307 12365
rect 4249 12356 4261 12359
rect 4212 12328 4261 12356
rect 4212 12316 4218 12328
rect 4249 12325 4261 12328
rect 4295 12325 4307 12359
rect 7650 12356 7656 12368
rect 4249 12319 4307 12325
rect 7208 12328 7656 12356
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12257 5963 12291
rect 6086 12288 6092 12300
rect 6047 12260 6092 12288
rect 5905 12251 5963 12257
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 2958 12220 2964 12232
rect 2823 12192 2964 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 4028 12192 4169 12220
rect 4028 12180 4034 12192
rect 4157 12189 4169 12192
rect 4203 12220 4215 12223
rect 4246 12220 4252 12232
rect 4203 12192 4252 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 5442 12220 5448 12232
rect 4847 12192 5448 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 5442 12180 5448 12192
rect 5500 12220 5506 12232
rect 5718 12220 5724 12232
rect 5500 12192 5724 12220
rect 5500 12180 5506 12192
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 5920 12220 5948 12251
rect 6086 12248 6092 12260
rect 6144 12288 6150 12300
rect 7208 12297 7236 12328
rect 7650 12316 7656 12328
rect 7708 12316 7714 12368
rect 6825 12291 6883 12297
rect 6825 12288 6837 12291
rect 6144 12260 6837 12288
rect 6144 12248 6150 12260
rect 6825 12257 6837 12260
rect 6871 12288 6883 12291
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 6871 12260 7205 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7742 12288 7748 12300
rect 7703 12260 7748 12288
rect 7193 12251 7251 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 5994 12220 6000 12232
rect 5920 12192 6000 12220
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 7852 12220 7880 12384
rect 9784 12356 9812 12384
rect 10039 12359 10097 12365
rect 10039 12356 10051 12359
rect 9784 12328 10051 12356
rect 10039 12325 10051 12328
rect 10085 12356 10097 12359
rect 10520 12356 10548 12396
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 11054 12424 11060 12436
rect 10643 12396 11060 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 13722 12424 13728 12436
rect 13683 12396 13728 12424
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 14332 12396 14657 12424
rect 14332 12384 14338 12396
rect 14645 12393 14657 12396
rect 14691 12393 14703 12427
rect 14645 12387 14703 12393
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 18601 12427 18659 12433
rect 18601 12424 18613 12427
rect 18196 12396 18613 12424
rect 18196 12384 18202 12396
rect 18601 12393 18613 12396
rect 18647 12393 18659 12427
rect 18601 12387 18659 12393
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 22462 12424 22468 12436
rect 22336 12396 22468 12424
rect 22336 12384 22342 12396
rect 22462 12384 22468 12396
rect 22520 12384 22526 12436
rect 10778 12356 10784 12368
rect 10085 12328 10456 12356
rect 10520 12328 10784 12356
rect 10085 12325 10097 12328
rect 10039 12319 10097 12325
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12288 8079 12291
rect 8478 12288 8484 12300
rect 8067 12260 8484 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8478 12248 8484 12260
rect 8536 12288 8542 12300
rect 9122 12288 9128 12300
rect 8536 12260 9128 12288
rect 8536 12248 8542 12260
rect 9122 12248 9128 12260
rect 9180 12248 9186 12300
rect 10428 12288 10456 12328
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 12437 12359 12495 12365
rect 12437 12325 12449 12359
rect 12483 12356 12495 12359
rect 12526 12356 12532 12368
rect 12483 12328 12532 12356
rect 12483 12325 12495 12328
rect 12437 12319 12495 12325
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 12989 12359 13047 12365
rect 12989 12325 13001 12359
rect 13035 12356 13047 12359
rect 14366 12356 14372 12368
rect 13035 12328 14372 12356
rect 13035 12325 13047 12328
rect 12989 12319 13047 12325
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 16206 12356 16212 12368
rect 16167 12328 16212 12356
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 17770 12356 17776 12368
rect 17683 12328 17776 12356
rect 17770 12316 17776 12328
rect 17828 12356 17834 12368
rect 18414 12356 18420 12368
rect 17828 12328 18420 12356
rect 17828 12316 17834 12328
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 11422 12288 11428 12300
rect 10428 12260 11428 12288
rect 11422 12248 11428 12260
rect 11480 12288 11486 12300
rect 12158 12288 12164 12300
rect 11480 12260 12164 12288
rect 11480 12248 11486 12260
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 14274 12288 14280 12300
rect 14231 12260 14280 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 19242 12288 19248 12300
rect 19203 12260 19248 12288
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 22278 12297 22284 12300
rect 20936 12291 20994 12297
rect 20936 12288 20948 12291
rect 20864 12260 20948 12288
rect 20864 12248 20870 12260
rect 20936 12257 20948 12260
rect 20982 12257 20994 12291
rect 20936 12251 20994 12257
rect 22256 12291 22284 12297
rect 22256 12257 22268 12291
rect 22256 12251 22284 12257
rect 22278 12248 22284 12251
rect 22336 12248 22342 12300
rect 23728 12291 23786 12297
rect 23728 12257 23740 12291
rect 23774 12288 23786 12291
rect 24118 12288 24124 12300
rect 23774 12260 24124 12288
rect 23774 12257 23786 12260
rect 23728 12251 23786 12257
rect 24118 12248 24124 12260
rect 24176 12248 24182 12300
rect 24762 12297 24768 12300
rect 24740 12291 24768 12297
rect 24740 12257 24752 12291
rect 24740 12251 24768 12257
rect 24762 12248 24768 12251
rect 24820 12248 24826 12300
rect 7708 12192 7880 12220
rect 7708 12180 7714 12192
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 8113 12223 8171 12229
rect 8113 12220 8125 12223
rect 7984 12192 8125 12220
rect 7984 12180 7990 12192
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 9364 12192 9689 12220
rect 9364 12180 9370 12192
rect 9651 12189 9689 12192
rect 9723 12220 9735 12223
rect 9723 12192 9784 12220
rect 9723 12189 9735 12192
rect 9651 12183 9735 12189
rect 1394 12112 1400 12164
rect 1452 12152 1458 12164
rect 8662 12152 8668 12164
rect 1452 12124 8668 12152
rect 1452 12112 1458 12124
rect 8662 12112 8668 12124
rect 8720 12112 8726 12164
rect 9651 12152 9679 12183
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10192 12192 10885 12220
rect 10192 12180 10198 12192
rect 10873 12189 10885 12192
rect 10919 12189 10931 12223
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 10873 12183 10931 12189
rect 12084 12192 12357 12220
rect 10594 12152 10600 12164
rect 9651 12124 10600 12152
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 1765 12087 1823 12093
rect 1765 12053 1777 12087
rect 1811 12084 1823 12087
rect 1854 12084 1860 12096
rect 1811 12056 1860 12084
rect 1811 12053 1823 12056
rect 1765 12047 1823 12053
rect 1854 12044 1860 12056
rect 1912 12084 1918 12096
rect 2130 12084 2136 12096
rect 1912 12056 2136 12084
rect 1912 12044 1918 12056
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 12084 12093 12112 12192
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 16117 12223 16175 12229
rect 16117 12189 16129 12223
rect 16163 12220 16175 12223
rect 16298 12220 16304 12232
rect 16163 12192 16304 12220
rect 16163 12189 16175 12192
rect 16117 12183 16175 12189
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 16758 12220 16764 12232
rect 16719 12192 16764 12220
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17678 12220 17684 12232
rect 17639 12192 17684 12220
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17954 12220 17960 12232
rect 17915 12192 17960 12220
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 14369 12155 14427 12161
rect 14369 12121 14381 12155
rect 14415 12152 14427 12155
rect 14826 12152 14832 12164
rect 14415 12124 14832 12152
rect 14415 12121 14427 12124
rect 14369 12115 14427 12121
rect 14826 12112 14832 12124
rect 14884 12112 14890 12164
rect 22094 12112 22100 12164
rect 22152 12152 22158 12164
rect 22327 12155 22385 12161
rect 22327 12152 22339 12155
rect 22152 12124 22339 12152
rect 22152 12112 22158 12124
rect 22327 12121 22339 12124
rect 22373 12121 22385 12155
rect 22327 12115 22385 12121
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 10744 12056 12081 12084
rect 10744 12044 10750 12056
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12069 12047 12127 12053
rect 15841 12087 15899 12093
rect 15841 12053 15853 12087
rect 15887 12084 15899 12087
rect 16022 12084 16028 12096
rect 15887 12056 16028 12084
rect 15887 12053 15899 12056
rect 15841 12047 15899 12053
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 17497 12087 17555 12093
rect 17497 12053 17509 12087
rect 17543 12084 17555 12087
rect 18138 12084 18144 12096
rect 17543 12056 18144 12084
rect 17543 12053 17555 12056
rect 17497 12047 17555 12053
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 19426 12084 19432 12096
rect 19387 12056 19432 12084
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 20714 12044 20720 12096
rect 20772 12084 20778 12096
rect 21039 12087 21097 12093
rect 21039 12084 21051 12087
rect 20772 12056 21051 12084
rect 20772 12044 20778 12056
rect 21039 12053 21051 12056
rect 21085 12053 21097 12087
rect 21039 12047 21097 12053
rect 22922 12044 22928 12096
rect 22980 12084 22986 12096
rect 23799 12087 23857 12093
rect 23799 12084 23811 12087
rect 22980 12056 23811 12084
rect 22980 12044 22986 12056
rect 23799 12053 23811 12056
rect 23845 12053 23857 12087
rect 23799 12047 23857 12053
rect 24811 12087 24869 12093
rect 24811 12053 24823 12087
rect 24857 12084 24869 12087
rect 24946 12084 24952 12096
rect 24857 12056 24952 12084
rect 24857 12053 24869 12056
rect 24811 12047 24869 12053
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 2041 11883 2099 11889
rect 2041 11849 2053 11883
rect 2087 11880 2099 11883
rect 2314 11880 2320 11892
rect 2087 11852 2320 11880
rect 2087 11849 2099 11852
rect 2041 11843 2099 11849
rect 2314 11840 2320 11852
rect 2372 11880 2378 11892
rect 2774 11880 2780 11892
rect 2372 11852 2780 11880
rect 2372 11840 2378 11852
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 5261 11883 5319 11889
rect 5261 11849 5273 11883
rect 5307 11880 5319 11883
rect 6086 11880 6092 11892
rect 5307 11852 6092 11880
rect 5307 11849 5319 11852
rect 5261 11843 5319 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 6914 11840 6920 11892
rect 6972 11880 6978 11892
rect 7374 11880 7380 11892
rect 6972 11852 7380 11880
rect 6972 11840 6978 11852
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 10594 11880 10600 11892
rect 10555 11852 10600 11880
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 15933 11883 15991 11889
rect 15933 11849 15945 11883
rect 15979 11880 15991 11883
rect 16206 11880 16212 11892
rect 15979 11852 16212 11880
rect 15979 11849 15991 11852
rect 15933 11843 15991 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16669 11883 16727 11889
rect 16669 11849 16681 11883
rect 16715 11880 16727 11883
rect 17678 11880 17684 11892
rect 16715 11852 17684 11880
rect 16715 11849 16727 11852
rect 16669 11843 16727 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 19058 11880 19064 11892
rect 19019 11852 19064 11880
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 22278 11880 22284 11892
rect 22239 11852 22284 11880
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 25133 11883 25191 11889
rect 25133 11880 25145 11883
rect 24820 11852 25145 11880
rect 24820 11840 24826 11852
rect 25133 11849 25145 11852
rect 25179 11849 25191 11883
rect 25133 11843 25191 11849
rect 3145 11815 3203 11821
rect 3145 11812 3157 11815
rect 2240 11784 3157 11812
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1578 11744 1584 11756
rect 1360 11716 1584 11744
rect 1360 11704 1366 11716
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 1670 11704 1676 11756
rect 1728 11744 1734 11756
rect 2240 11753 2268 11784
rect 3145 11781 3157 11784
rect 3191 11781 3203 11815
rect 3145 11775 3203 11781
rect 3510 11772 3516 11824
rect 3568 11812 3574 11824
rect 3694 11812 3700 11824
rect 3568 11784 3700 11812
rect 3568 11772 3574 11784
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 5629 11815 5687 11821
rect 5629 11781 5641 11815
rect 5675 11812 5687 11815
rect 5905 11815 5963 11821
rect 5905 11812 5917 11815
rect 5675 11784 5917 11812
rect 5675 11781 5687 11784
rect 5629 11775 5687 11781
rect 5905 11781 5917 11784
rect 5951 11812 5963 11815
rect 5994 11812 6000 11824
rect 5951 11784 6000 11812
rect 5951 11781 5963 11784
rect 5905 11775 5963 11781
rect 5994 11772 6000 11784
rect 6052 11812 6058 11824
rect 6730 11812 6736 11824
rect 6052 11784 6736 11812
rect 6052 11772 6058 11784
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 8297 11815 8355 11821
rect 8297 11781 8309 11815
rect 8343 11812 8355 11815
rect 8478 11812 8484 11824
rect 8343 11784 8484 11812
rect 8343 11781 8355 11784
rect 8297 11775 8355 11781
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 10318 11812 10324 11824
rect 10279 11784 10324 11812
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 11425 11815 11483 11821
rect 11425 11781 11437 11815
rect 11471 11812 11483 11815
rect 12342 11812 12348 11824
rect 11471 11784 12348 11812
rect 11471 11781 11483 11784
rect 11425 11775 11483 11781
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 1728 11716 2237 11744
rect 1728 11704 1734 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 2406 11704 2412 11756
rect 2464 11744 2470 11756
rect 3786 11744 3792 11756
rect 2464 11716 3792 11744
rect 2464 11704 2470 11716
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7282 11744 7288 11756
rect 6963 11716 7288 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9490 11744 9496 11756
rect 9447 11716 9496 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12676 11716 12725 11744
rect 12676 11704 12682 11716
rect 12713 11713 12725 11716
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15010 11744 15016 11756
rect 14700 11716 15016 11744
rect 14700 11704 14706 11716
rect 15010 11704 15016 11716
rect 15068 11704 15074 11756
rect 18138 11744 18144 11756
rect 18099 11716 18144 11744
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 18230 11704 18236 11756
rect 18288 11744 18294 11756
rect 18417 11747 18475 11753
rect 18417 11744 18429 11747
rect 18288 11716 18429 11744
rect 18288 11704 18294 11716
rect 18417 11713 18429 11716
rect 18463 11713 18475 11747
rect 19076 11744 19104 11840
rect 24489 11815 24547 11821
rect 24489 11812 24501 11815
rect 23722 11784 24501 11812
rect 19705 11747 19763 11753
rect 19705 11744 19717 11747
rect 19076 11716 19717 11744
rect 18417 11707 18475 11713
rect 19705 11713 19717 11716
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 5997 11679 6055 11685
rect 5997 11676 6009 11679
rect 5767 11648 6009 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 5997 11645 6009 11648
rect 6043 11645 6055 11679
rect 5997 11639 6055 11645
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 8424 11679 8482 11685
rect 8424 11676 8436 11679
rect 7892 11648 8436 11676
rect 7892 11636 7898 11648
rect 8404 11645 8436 11648
rect 8470 11645 8482 11679
rect 8404 11639 8482 11645
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11676 11299 11679
rect 14274 11676 14280 11688
rect 11287 11648 11744 11676
rect 14187 11648 14280 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 2222 11568 2228 11620
rect 2280 11608 2286 11620
rect 2317 11611 2375 11617
rect 2317 11608 2329 11611
rect 2280 11580 2329 11608
rect 2280 11568 2286 11580
rect 2317 11577 2329 11580
rect 2363 11577 2375 11611
rect 2317 11571 2375 11577
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 2958 11608 2964 11620
rect 2915 11580 2964 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 2958 11568 2964 11580
rect 3016 11568 3022 11620
rect 3881 11611 3939 11617
rect 3881 11577 3893 11611
rect 3927 11577 3939 11611
rect 3881 11571 3939 11577
rect 4433 11611 4491 11617
rect 4433 11577 4445 11611
rect 4479 11608 4491 11611
rect 5810 11608 5816 11620
rect 4479 11580 5816 11608
rect 4479 11577 4491 11580
rect 4433 11571 4491 11577
rect 3602 11540 3608 11552
rect 3515 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11540 3666 11552
rect 3896 11540 3924 11571
rect 5810 11568 5816 11580
rect 5868 11608 5874 11620
rect 5868 11580 6500 11608
rect 5868 11568 5874 11580
rect 4154 11540 4160 11552
rect 3660 11512 4160 11540
rect 3660 11500 3666 11512
rect 4154 11500 4160 11512
rect 4212 11540 4218 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 4212 11512 4721 11540
rect 4212 11500 4218 11512
rect 4709 11509 4721 11512
rect 4755 11509 4767 11543
rect 4709 11503 4767 11509
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6273 11543 6331 11549
rect 6273 11540 6285 11543
rect 6043 11512 6285 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6273 11509 6285 11512
rect 6319 11540 6331 11543
rect 6362 11540 6368 11552
rect 6319 11512 6368 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 6472 11540 6500 11580
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 6914 11608 6920 11620
rect 6604 11580 6920 11608
rect 6604 11568 6610 11580
rect 6914 11568 6920 11580
rect 6972 11608 6978 11620
rect 7009 11611 7067 11617
rect 7009 11608 7021 11611
rect 6972 11580 7021 11608
rect 6972 11568 6978 11580
rect 7009 11577 7021 11580
rect 7055 11577 7067 11611
rect 7009 11571 7067 11577
rect 7561 11611 7619 11617
rect 7561 11577 7573 11611
rect 7607 11577 7619 11611
rect 7561 11571 7619 11577
rect 7576 11540 7604 11571
rect 7834 11540 7840 11552
rect 6472 11512 7604 11540
rect 7795 11512 7840 11540
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8404 11540 8432 11639
rect 8527 11611 8585 11617
rect 8527 11577 8539 11611
rect 8573 11608 8585 11611
rect 9582 11608 9588 11620
rect 8573 11580 9588 11608
rect 8573 11577 8585 11580
rect 8527 11571 8585 11577
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 9722 11611 9780 11617
rect 9722 11577 9734 11611
rect 9768 11577 9780 11611
rect 9722 11571 9780 11577
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 8404 11512 8953 11540
rect 8941 11509 8953 11512
rect 8987 11540 8999 11543
rect 9030 11540 9036 11552
rect 8987 11512 9036 11540
rect 8987 11509 8999 11512
rect 8941 11503 8999 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9309 11543 9367 11549
rect 9309 11509 9321 11543
rect 9355 11540 9367 11543
rect 9490 11540 9496 11552
rect 9355 11512 9496 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9490 11500 9496 11512
rect 9548 11540 9554 11552
rect 9737 11540 9765 11571
rect 11716 11552 11744 11648
rect 14274 11636 14280 11648
rect 14332 11676 14338 11688
rect 14826 11676 14832 11688
rect 14332 11648 14832 11676
rect 14332 11636 14338 11648
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 16758 11676 16764 11688
rect 16719 11648 16764 11676
rect 16758 11636 16764 11648
rect 16816 11676 16822 11688
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 16816 11648 17233 11676
rect 16816 11636 16822 11648
rect 17221 11645 17233 11648
rect 17267 11645 17279 11679
rect 21266 11676 21272 11688
rect 21227 11648 21272 11676
rect 17221 11639 17279 11645
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 23474 11636 23480 11688
rect 23532 11676 23538 11688
rect 23722 11685 23750 11784
rect 24489 11781 24501 11784
rect 24535 11781 24547 11815
rect 24489 11775 24547 11781
rect 23934 11704 23940 11756
rect 23992 11704 23998 11756
rect 23707 11679 23765 11685
rect 23707 11676 23719 11679
rect 23532 11648 23719 11676
rect 23532 11636 23538 11648
rect 23707 11645 23719 11648
rect 23753 11645 23765 11679
rect 23707 11639 23765 11645
rect 15378 11617 15384 11620
rect 13034 11611 13092 11617
rect 13034 11608 13046 11611
rect 12268 11580 13046 11608
rect 12268 11552 12296 11580
rect 13034 11577 13046 11580
rect 13080 11608 13092 11611
rect 14921 11611 14979 11617
rect 14921 11608 14933 11611
rect 13080 11580 14933 11608
rect 13080 11577 13092 11580
rect 13034 11571 13092 11577
rect 14921 11577 14933 11580
rect 14967 11608 14979 11611
rect 15334 11611 15384 11617
rect 15334 11608 15346 11611
rect 14967 11580 15346 11608
rect 14967 11577 14979 11580
rect 14921 11571 14979 11577
rect 15334 11577 15346 11580
rect 15380 11577 15384 11611
rect 15334 11571 15384 11577
rect 15378 11568 15384 11571
rect 15436 11608 15442 11620
rect 15838 11608 15844 11620
rect 15436 11580 15844 11608
rect 15436 11568 15442 11580
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 17126 11568 17132 11620
rect 17184 11608 17190 11620
rect 17865 11611 17923 11617
rect 17865 11608 17877 11611
rect 17184 11580 17877 11608
rect 17184 11568 17190 11580
rect 17865 11577 17877 11580
rect 17911 11608 17923 11611
rect 18233 11611 18291 11617
rect 18233 11608 18245 11611
rect 17911 11580 18245 11608
rect 17911 11577 17923 11580
rect 17865 11571 17923 11577
rect 18233 11577 18245 11580
rect 18279 11577 18291 11611
rect 18233 11571 18291 11577
rect 19426 11568 19432 11620
rect 19484 11608 19490 11620
rect 19797 11611 19855 11617
rect 19797 11608 19809 11611
rect 19484 11580 19809 11608
rect 19484 11568 19490 11580
rect 19797 11577 19809 11580
rect 19843 11577 19855 11611
rect 20346 11608 20352 11620
rect 20307 11580 20352 11608
rect 19797 11571 19855 11577
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 11698 11540 11704 11552
rect 9548 11512 9765 11540
rect 11659 11512 11704 11540
rect 9548 11500 9554 11512
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12250 11540 12256 11552
rect 12211 11512 12256 11540
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 13633 11543 13691 11549
rect 13633 11540 13645 11543
rect 13320 11512 13645 11540
rect 13320 11500 13326 11512
rect 13633 11509 13645 11512
rect 13679 11509 13691 11543
rect 13633 11503 13691 11509
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16390 11540 16396 11552
rect 16264 11512 16396 11540
rect 16264 11500 16270 11512
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16942 11540 16948 11552
rect 16903 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 20901 11543 20959 11549
rect 20901 11540 20913 11543
rect 20864 11512 20913 11540
rect 20864 11500 20870 11512
rect 20901 11509 20913 11512
rect 20947 11509 20959 11543
rect 21634 11540 21640 11552
rect 21595 11512 21640 11540
rect 20901 11503 20959 11509
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 23658 11500 23664 11552
rect 23716 11540 23722 11552
rect 23799 11543 23857 11549
rect 23799 11540 23811 11543
rect 23716 11512 23811 11540
rect 23716 11500 23722 11512
rect 23799 11509 23811 11512
rect 23845 11509 23857 11543
rect 23952 11540 23980 11704
rect 24118 11676 24124 11688
rect 24079 11648 24124 11676
rect 24118 11636 24124 11648
rect 24176 11636 24182 11688
rect 24302 11636 24308 11688
rect 24360 11676 24366 11688
rect 24740 11679 24798 11685
rect 24740 11676 24752 11679
rect 24360 11648 24752 11676
rect 24360 11636 24366 11648
rect 24740 11645 24752 11648
rect 24786 11676 24798 11679
rect 25501 11679 25559 11685
rect 25501 11676 25513 11679
rect 24786 11648 25513 11676
rect 24786 11645 24798 11648
rect 24740 11639 24798 11645
rect 25501 11645 25513 11648
rect 25547 11645 25559 11679
rect 25501 11639 25559 11645
rect 24118 11540 24124 11552
rect 23952 11512 24124 11540
rect 23799 11503 23857 11509
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24394 11500 24400 11552
rect 24452 11540 24458 11552
rect 24811 11543 24869 11549
rect 24811 11540 24823 11543
rect 24452 11512 24823 11540
rect 24452 11500 24458 11512
rect 24811 11509 24823 11512
rect 24857 11509 24869 11543
rect 24811 11503 24869 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1535 11339 1593 11345
rect 1535 11305 1547 11339
rect 1581 11336 1593 11339
rect 1946 11336 1952 11348
rect 1581 11308 1952 11336
rect 1581 11305 1593 11308
rect 1535 11299 1593 11305
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2222 11336 2228 11348
rect 2183 11308 2228 11336
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4246 11336 4252 11348
rect 4207 11308 4252 11336
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5368 11308 5733 11336
rect 5368 11280 5396 11308
rect 5721 11305 5733 11308
rect 5767 11336 5779 11339
rect 5810 11336 5816 11348
rect 5767 11308 5816 11336
rect 5767 11305 5779 11308
rect 5721 11299 5779 11305
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7340 11308 7389 11336
rect 7340 11296 7346 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 9490 11336 9496 11348
rect 9451 11308 9496 11336
rect 7377 11299 7435 11305
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 12526 11336 12532 11348
rect 12487 11308 12532 11336
rect 12526 11296 12532 11308
rect 12584 11336 12590 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 12584 11308 12817 11336
rect 12584 11296 12590 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 15010 11336 15016 11348
rect 14971 11308 15016 11336
rect 12805 11299 12863 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 16298 11336 16304 11348
rect 16259 11308 16304 11336
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 18141 11339 18199 11345
rect 18141 11305 18153 11339
rect 18187 11305 18199 11339
rect 18414 11336 18420 11348
rect 18375 11308 18420 11336
rect 18141 11299 18199 11305
rect 2498 11268 2504 11280
rect 2459 11240 2504 11268
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 2593 11271 2651 11277
rect 2593 11237 2605 11271
rect 2639 11268 2651 11271
rect 3142 11268 3148 11280
rect 2639 11240 3148 11268
rect 2639 11237 2651 11240
rect 2593 11231 2651 11237
rect 3142 11228 3148 11240
rect 3200 11268 3206 11280
rect 3602 11268 3608 11280
rect 3200 11240 3608 11268
rect 3200 11228 3206 11240
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 4798 11268 4804 11280
rect 4212 11240 4804 11268
rect 4212 11228 4218 11240
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 5350 11268 5356 11280
rect 5263 11240 5356 11268
rect 5350 11228 5356 11240
rect 5408 11228 5414 11280
rect 6546 11277 6552 11280
rect 6543 11268 6552 11277
rect 6507 11240 6552 11268
rect 6543 11231 6552 11240
rect 6546 11228 6552 11231
rect 6604 11228 6610 11280
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 8168 11240 8217 11268
rect 8168 11228 8174 11240
rect 8205 11237 8217 11240
rect 8251 11268 8263 11271
rect 8386 11268 8392 11280
rect 8251 11240 8392 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 9508 11268 9536 11296
rect 9998 11271 10056 11277
rect 9998 11268 10010 11271
rect 9508 11240 10010 11268
rect 9998 11237 10010 11240
rect 10044 11237 10056 11271
rect 9998 11231 10056 11237
rect 11971 11271 12029 11277
rect 11971 11237 11983 11271
rect 12017 11268 12029 11271
rect 12250 11268 12256 11280
rect 12017 11240 12256 11268
rect 12017 11237 12029 11240
rect 11971 11231 12029 11237
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12676 11240 13185 11268
rect 12676 11228 12682 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 13262 11228 13268 11280
rect 13320 11268 13326 11280
rect 13817 11271 13875 11277
rect 13817 11268 13829 11271
rect 13320 11240 13829 11268
rect 13320 11228 13326 11240
rect 13817 11237 13829 11240
rect 13863 11237 13875 11271
rect 14366 11268 14372 11280
rect 14327 11240 14372 11268
rect 13817 11231 13875 11237
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 15470 11268 15476 11280
rect 15431 11240 15476 11268
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 17542 11271 17600 11277
rect 17542 11268 17554 11271
rect 17460 11240 17554 11268
rect 17460 11228 17466 11240
rect 17542 11237 17554 11240
rect 17588 11237 17600 11271
rect 18156 11268 18184 11299
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 19981 11339 20039 11345
rect 19981 11336 19993 11339
rect 19260 11308 19993 11336
rect 19260 11280 19288 11308
rect 19981 11305 19993 11308
rect 20027 11305 20039 11339
rect 21266 11336 21272 11348
rect 21227 11308 21272 11336
rect 19981 11299 20039 11305
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 18877 11271 18935 11277
rect 18877 11268 18889 11271
rect 18156 11240 18889 11268
rect 17542 11231 17600 11237
rect 18877 11237 18889 11240
rect 18923 11268 18935 11271
rect 19153 11271 19211 11277
rect 19153 11268 19165 11271
rect 18923 11240 19165 11268
rect 18923 11237 18935 11240
rect 18877 11231 18935 11237
rect 19153 11237 19165 11240
rect 19199 11268 19211 11271
rect 19242 11268 19248 11280
rect 19199 11240 19248 11268
rect 19199 11237 19211 11240
rect 19153 11231 19211 11237
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 19705 11271 19763 11277
rect 19705 11237 19717 11271
rect 19751 11268 19763 11271
rect 20346 11268 20352 11280
rect 19751 11240 20352 11268
rect 19751 11237 19763 11240
rect 19705 11231 19763 11237
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 21634 11228 21640 11280
rect 21692 11268 21698 11280
rect 21729 11271 21787 11277
rect 21729 11268 21741 11271
rect 21692 11240 21741 11268
rect 21692 11228 21698 11240
rect 21729 11237 21741 11240
rect 21775 11237 21787 11271
rect 21729 11231 21787 11237
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11200 1522 11203
rect 1670 11200 1676 11212
rect 1510 11172 1676 11200
rect 1510 11169 1522 11172
rect 1464 11163 1522 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6972 11172 7113 11200
rect 6972 11160 6978 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9456 11172 9689 11200
rect 9456 11160 9462 11172
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 11790 11200 11796 11212
rect 11655 11172 11796 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 23604 11203 23662 11209
rect 23604 11200 23616 11203
rect 23492 11172 23616 11200
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 4212 11104 4721 11132
rect 4212 11092 4218 11104
rect 4709 11101 4721 11104
rect 4755 11132 4767 11135
rect 4890 11132 4896 11144
rect 4755 11104 4896 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11132 6239 11135
rect 7929 11135 7987 11141
rect 6227 11104 6261 11132
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7975 11104 8125 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8113 11101 8125 11104
rect 8159 11132 8171 11135
rect 8202 11132 8208 11144
rect 8159 11104 8208 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 2958 11024 2964 11076
rect 3016 11064 3022 11076
rect 3053 11067 3111 11073
rect 3053 11064 3065 11067
rect 3016 11036 3065 11064
rect 3016 11024 3022 11036
rect 3053 11033 3065 11036
rect 3099 11064 3111 11067
rect 6089 11067 6147 11073
rect 3099 11036 4108 11064
rect 3099 11033 3111 11036
rect 3053 11027 3111 11033
rect 4080 10996 4108 11036
rect 6089 11033 6101 11067
rect 6135 11064 6147 11067
rect 6196 11064 6224 11095
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9766 11132 9772 11144
rect 8803 11104 9772 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 13722 11132 13728 11144
rect 13683 11104 13728 11132
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 15378 11132 15384 11144
rect 15339 11104 15384 11132
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 6135 11036 6868 11064
rect 6135 11033 6147 11036
rect 6089 11027 6147 11033
rect 4246 10996 4252 11008
rect 4080 10968 4252 10996
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 6840 10996 6868 11036
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 8478 11064 8484 11076
rect 7340 11036 8484 11064
rect 7340 11024 7346 11036
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 15672 11064 15700 11095
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 16632 11104 17049 11132
rect 16632 11092 16638 11104
rect 17037 11101 17049 11104
rect 17083 11132 17095 11135
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 17083 11104 17233 11132
rect 17083 11101 17095 11104
rect 17037 11095 17095 11101
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 19061 11135 19119 11141
rect 19061 11132 19073 11135
rect 18288 11104 19073 11132
rect 18288 11092 18294 11104
rect 19061 11101 19073 11104
rect 19107 11132 19119 11135
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 19107 11104 20361 11132
rect 19107 11101 19119 11104
rect 19061 11095 19119 11101
rect 20349 11101 20361 11104
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11132 21695 11135
rect 22094 11132 22100 11144
rect 21683 11104 22100 11132
rect 21683 11101 21695 11104
rect 21637 11095 21695 11101
rect 22094 11092 22100 11104
rect 22152 11092 22158 11144
rect 15120 11036 15700 11064
rect 22189 11067 22247 11073
rect 6914 10996 6920 11008
rect 6840 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 10597 10999 10655 11005
rect 10597 10965 10609 10999
rect 10643 10996 10655 10999
rect 11054 10996 11060 11008
rect 10643 10968 11060 10996
rect 10643 10965 10655 10968
rect 10597 10959 10655 10965
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 15120 10996 15148 11036
rect 22189 11033 22201 11067
rect 22235 11033 22247 11067
rect 23492 11064 23520 11172
rect 23604 11169 23616 11172
rect 23650 11169 23662 11203
rect 23604 11163 23662 11169
rect 24210 11160 24216 11212
rect 24268 11200 24274 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24268 11172 24593 11200
rect 24268 11160 24274 11172
rect 24581 11169 24593 11172
rect 24627 11200 24639 11203
rect 24670 11200 24676 11212
rect 24627 11172 24676 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 23934 11092 23940 11144
rect 23992 11132 23998 11144
rect 24394 11132 24400 11144
rect 23992 11104 24400 11132
rect 23992 11092 23998 11104
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 22189 11027 22247 11033
rect 23400 11036 23520 11064
rect 23707 11067 23765 11073
rect 13872 10968 15148 10996
rect 13872 10956 13878 10968
rect 21818 10956 21824 11008
rect 21876 10996 21882 11008
rect 22204 10996 22232 11027
rect 21876 10968 22232 10996
rect 21876 10956 21882 10968
rect 23014 10956 23020 11008
rect 23072 10996 23078 11008
rect 23400 10996 23428 11036
rect 23707 11033 23719 11067
rect 23753 11064 23765 11067
rect 24854 11064 24860 11076
rect 23753 11036 24860 11064
rect 23753 11033 23765 11036
rect 23707 11027 23765 11033
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 24762 10996 24768 11008
rect 23072 10968 23428 10996
rect 24723 10968 24768 10996
rect 23072 10956 23078 10968
rect 24762 10956 24768 10968
rect 24820 10956 24826 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 3142 10792 3148 10804
rect 3099 10764 3148 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9677 10795 9735 10801
rect 9677 10792 9689 10795
rect 9548 10764 9689 10792
rect 9548 10752 9554 10764
rect 9677 10761 9689 10764
rect 9723 10761 9735 10795
rect 9677 10755 9735 10761
rect 10686 10752 10692 10804
rect 10744 10752 10750 10804
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 11977 10795 12035 10801
rect 11977 10792 11989 10795
rect 11848 10764 11989 10792
rect 11848 10752 11854 10764
rect 11977 10761 11989 10764
rect 12023 10761 12035 10795
rect 13262 10792 13268 10804
rect 13223 10764 13268 10792
rect 11977 10755 12035 10761
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15470 10792 15476 10804
rect 15427 10764 15476 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15896 10764 16037 10792
rect 15896 10752 15902 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 17126 10792 17132 10804
rect 17087 10764 17132 10792
rect 16025 10755 16083 10761
rect 2498 10684 2504 10736
rect 2556 10724 2562 10736
rect 3329 10727 3387 10733
rect 3329 10724 3341 10727
rect 2556 10696 3341 10724
rect 2556 10684 2562 10696
rect 3329 10693 3341 10696
rect 3375 10693 3387 10727
rect 3329 10687 3387 10693
rect 4525 10727 4583 10733
rect 4525 10693 4537 10727
rect 4571 10724 4583 10727
rect 5166 10724 5172 10736
rect 4571 10696 5172 10724
rect 4571 10693 4583 10696
rect 4525 10687 4583 10693
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 3881 10591 3939 10597
rect 2179 10560 2728 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2038 10520 2044 10532
rect 1951 10492 2044 10520
rect 2038 10480 2044 10492
rect 2096 10520 2102 10532
rect 2498 10529 2504 10532
rect 2454 10523 2504 10529
rect 2454 10520 2466 10523
rect 2096 10492 2466 10520
rect 2096 10480 2102 10492
rect 2454 10489 2466 10492
rect 2500 10489 2504 10523
rect 2454 10483 2504 10489
rect 2498 10480 2504 10483
rect 2556 10480 2562 10532
rect 2700 10452 2728 10560
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 4540 10588 4568 10687
rect 5166 10684 5172 10696
rect 5224 10724 5230 10736
rect 7742 10724 7748 10736
rect 5224 10696 7748 10724
rect 5224 10684 5230 10696
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 9766 10684 9772 10736
rect 9824 10724 9830 10736
rect 10597 10727 10655 10733
rect 10597 10724 10609 10727
rect 9824 10696 10609 10724
rect 9824 10684 9830 10696
rect 10597 10693 10609 10696
rect 10643 10724 10655 10727
rect 10704 10724 10732 10752
rect 10643 10696 10732 10724
rect 10643 10693 10655 10696
rect 10597 10687 10655 10693
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5350 10656 5356 10668
rect 5307 10628 5356 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 5994 10656 6000 10668
rect 5951 10628 6000 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 5994 10616 6000 10628
rect 6052 10656 6058 10668
rect 6178 10656 6184 10668
rect 6052 10628 6184 10656
rect 6052 10616 6058 10628
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 8202 10656 8208 10668
rect 7392 10628 8208 10656
rect 3927 10560 4568 10588
rect 6641 10591 6699 10597
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7098 10588 7104 10600
rect 6687 10560 7104 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 7392 10597 7420 10628
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 9732 10628 10057 10656
rect 9732 10616 9738 10628
rect 10045 10625 10057 10628
rect 10091 10656 10103 10659
rect 10134 10656 10140 10668
rect 10091 10628 10140 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14093 10659 14151 10665
rect 14093 10656 14105 10659
rect 13872 10628 14105 10656
rect 13872 10616 13878 10628
rect 14093 10625 14105 10628
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 15013 10659 15071 10665
rect 15013 10625 15025 10659
rect 15059 10656 15071 10659
rect 15378 10656 15384 10668
rect 15059 10628 15384 10656
rect 15059 10625 15071 10628
rect 15013 10619 15071 10625
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 16040 10656 16068 10755
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 20990 10792 20996 10804
rect 20951 10764 20996 10792
rect 20990 10752 20996 10764
rect 21048 10792 21054 10804
rect 21453 10795 21511 10801
rect 21048 10764 21404 10792
rect 21048 10752 21054 10764
rect 20717 10727 20775 10733
rect 20717 10693 20729 10727
rect 20763 10724 20775 10727
rect 21266 10724 21272 10736
rect 20763 10696 21272 10724
rect 20763 10693 20775 10696
rect 20717 10687 20775 10693
rect 21266 10684 21272 10696
rect 21324 10684 21330 10736
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 16040 10628 16344 10656
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 7892 10560 8309 10588
rect 7892 10548 7898 10560
rect 8297 10557 8309 10560
rect 8343 10588 8355 10591
rect 8662 10588 8668 10600
rect 8343 10560 8668 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 8849 10551 8907 10557
rect 15764 10560 16221 10588
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 5408 10492 5453 10520
rect 5408 10480 5414 10492
rect 7650 10480 7656 10532
rect 7708 10520 7714 10532
rect 8864 10520 8892 10551
rect 7708 10492 8892 10520
rect 10137 10523 10195 10529
rect 7708 10480 7714 10492
rect 7852 10464 7880 10492
rect 10137 10489 10149 10523
rect 10183 10489 10195 10523
rect 10137 10483 10195 10489
rect 12713 10523 12771 10529
rect 12713 10489 12725 10523
rect 12759 10520 12771 10523
rect 13541 10523 13599 10529
rect 13541 10520 13553 10523
rect 12759 10492 13553 10520
rect 12759 10489 12771 10492
rect 12713 10483 12771 10489
rect 13541 10489 13553 10492
rect 13587 10520 13599 10523
rect 13817 10523 13875 10529
rect 13817 10520 13829 10523
rect 13587 10492 13829 10520
rect 13587 10489 13599 10492
rect 13541 10483 13599 10489
rect 13817 10489 13829 10492
rect 13863 10489 13875 10523
rect 13817 10483 13875 10489
rect 3602 10452 3608 10464
rect 2700 10424 3608 10452
rect 3602 10412 3608 10424
rect 3660 10452 3666 10464
rect 3697 10455 3755 10461
rect 3697 10452 3709 10455
rect 3660 10424 3709 10452
rect 3660 10412 3666 10424
rect 3697 10421 3709 10424
rect 3743 10421 3755 10455
rect 3697 10415 3755 10421
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 3844 10424 4077 10452
rect 3844 10412 3850 10424
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 6178 10452 6184 10464
rect 5224 10424 6184 10452
rect 5224 10412 5230 10424
rect 6178 10412 6184 10424
rect 6236 10452 6242 10464
rect 6546 10452 6552 10464
rect 6236 10424 6552 10452
rect 6236 10412 6242 10424
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6914 10452 6920 10464
rect 6875 10424 6920 10452
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7834 10452 7840 10464
rect 7795 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 8481 10455 8539 10461
rect 8481 10452 8493 10455
rect 8352 10424 8493 10452
rect 8352 10412 8358 10424
rect 8481 10421 8493 10424
rect 8527 10421 8539 10455
rect 10152 10452 10180 10483
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 15102 10520 15108 10532
rect 13964 10492 15108 10520
rect 13964 10480 13970 10492
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 15764 10464 15792 10560
rect 16209 10557 16221 10560
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16316 10520 16344 10628
rect 17788 10628 18153 10656
rect 16530 10523 16588 10529
rect 16530 10520 16542 10523
rect 16316 10492 16542 10520
rect 16530 10489 16542 10492
rect 16576 10520 16588 10523
rect 17402 10520 17408 10532
rect 16576 10492 17408 10520
rect 16576 10489 16588 10492
rect 16530 10483 16588 10489
rect 17402 10480 17408 10492
rect 17460 10480 17466 10532
rect 11054 10452 11060 10464
rect 10152 10424 11060 10452
rect 8481 10415 8539 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10452 11759 10455
rect 12250 10452 12256 10464
rect 11747 10424 12256 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 15746 10452 15752 10464
rect 15707 10424 15752 10452
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17788 10461 17816 10628
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 21376 10656 21404 10764
rect 21453 10761 21465 10795
rect 21499 10792 21511 10795
rect 21634 10792 21640 10804
rect 21499 10764 21640 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 21634 10752 21640 10764
rect 21692 10752 21698 10804
rect 22094 10752 22100 10804
rect 22152 10792 22158 10804
rect 22557 10795 22615 10801
rect 22557 10792 22569 10795
rect 22152 10764 22569 10792
rect 22152 10752 22158 10764
rect 22557 10761 22569 10764
rect 22603 10761 22615 10795
rect 23014 10792 23020 10804
rect 22975 10764 23020 10792
rect 22557 10755 22615 10761
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 21637 10659 21695 10665
rect 21637 10656 21649 10659
rect 21376 10628 21649 10656
rect 18141 10619 18199 10625
rect 21637 10625 21649 10628
rect 21683 10625 21695 10659
rect 21637 10619 21695 10625
rect 21818 10616 21824 10668
rect 21876 10656 21882 10668
rect 21913 10659 21971 10665
rect 21913 10656 21925 10659
rect 21876 10628 21925 10656
rect 21876 10616 21882 10628
rect 21913 10625 21925 10628
rect 21959 10625 21971 10659
rect 21913 10619 21971 10625
rect 24670 10616 24676 10668
rect 24728 10656 24734 10668
rect 25130 10656 25136 10668
rect 24728 10628 25136 10656
rect 24728 10616 24734 10628
rect 25130 10616 25136 10628
rect 25188 10616 25194 10668
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18322 10588 18328 10600
rect 18283 10560 18328 10588
rect 18049 10551 18107 10557
rect 18064 10520 18092 10551
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 19797 10591 19855 10597
rect 19797 10588 19809 10591
rect 19536 10560 19809 10588
rect 18230 10520 18236 10532
rect 18064 10492 18236 10520
rect 18230 10480 18236 10492
rect 18288 10480 18294 10532
rect 19536 10464 19564 10560
rect 19797 10557 19809 10560
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 23477 10591 23535 10597
rect 23477 10557 23489 10591
rect 23523 10588 23535 10591
rect 23753 10591 23811 10597
rect 23753 10588 23765 10591
rect 23523 10560 23765 10588
rect 23523 10557 23535 10560
rect 23477 10551 23535 10557
rect 23753 10557 23765 10560
rect 23799 10588 23811 10591
rect 23842 10588 23848 10600
rect 23799 10560 23848 10588
rect 23799 10557 23811 10560
rect 23753 10551 23811 10557
rect 23842 10548 23848 10560
rect 23900 10548 23906 10600
rect 24854 10548 24860 10600
rect 24912 10588 24918 10600
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 24912 10560 25237 10588
rect 24912 10548 24918 10560
rect 25225 10557 25237 10560
rect 25271 10588 25283 10591
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25271 10560 25789 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 20159 10523 20217 10529
rect 20159 10489 20171 10523
rect 20205 10489 20217 10523
rect 20159 10483 20217 10489
rect 21729 10523 21787 10529
rect 21729 10489 21741 10523
rect 21775 10489 21787 10523
rect 21729 10483 21787 10489
rect 24397 10523 24455 10529
rect 24397 10489 24409 10523
rect 24443 10520 24455 10523
rect 25038 10520 25044 10532
rect 24443 10492 25044 10520
rect 24443 10489 24455 10492
rect 24397 10483 24455 10489
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 17000 10424 17785 10452
rect 17000 10412 17006 10424
rect 17773 10421 17785 10424
rect 17819 10421 17831 10455
rect 18506 10452 18512 10464
rect 18467 10424 18512 10452
rect 17773 10415 17831 10421
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 19337 10455 19395 10461
rect 19337 10421 19349 10455
rect 19383 10452 19395 10455
rect 19518 10452 19524 10464
rect 19383 10424 19524 10452
rect 19383 10421 19395 10424
rect 19337 10415 19395 10421
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19705 10455 19763 10461
rect 19705 10421 19717 10455
rect 19751 10452 19763 10455
rect 20180 10452 20208 10483
rect 20346 10452 20352 10464
rect 19751 10424 20352 10452
rect 19751 10421 19763 10424
rect 19705 10415 19763 10421
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21744 10452 21772 10483
rect 25038 10480 25044 10492
rect 25096 10480 25102 10532
rect 21324 10424 21772 10452
rect 21324 10412 21330 10424
rect 23106 10412 23112 10464
rect 23164 10452 23170 10464
rect 23474 10452 23480 10464
rect 23164 10424 23480 10452
rect 23164 10412 23170 10424
rect 23474 10412 23480 10424
rect 23532 10412 23538 10464
rect 25406 10452 25412 10464
rect 25367 10424 25412 10452
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 2832 10220 2881 10248
rect 2832 10208 2838 10220
rect 2869 10217 2881 10220
rect 2915 10217 2927 10251
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 2869 10211 2927 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3881 10251 3939 10257
rect 3881 10217 3893 10251
rect 3927 10248 3939 10251
rect 4062 10248 4068 10260
rect 3927 10220 4068 10248
rect 3927 10217 3939 10220
rect 3881 10211 3939 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5537 10251 5595 10257
rect 5537 10248 5549 10251
rect 5500 10220 5549 10248
rect 5500 10208 5506 10220
rect 5537 10217 5549 10220
rect 5583 10217 5595 10251
rect 7650 10248 7656 10260
rect 7611 10220 7656 10248
rect 5537 10211 5595 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8444 10220 8585 10248
rect 8444 10208 8450 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 9398 10248 9404 10260
rect 9359 10220 9404 10248
rect 8573 10211 8631 10217
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10192 10220 10701 10248
rect 10192 10208 10198 10220
rect 10689 10217 10701 10220
rect 10735 10217 10747 10251
rect 11514 10248 11520 10260
rect 11475 10220 11520 10248
rect 10689 10211 10747 10217
rect 11514 10208 11520 10220
rect 11572 10248 11578 10260
rect 13354 10248 13360 10260
rect 11572 10220 13216 10248
rect 13315 10220 13360 10248
rect 11572 10208 11578 10220
rect 2311 10183 2369 10189
rect 2311 10149 2323 10183
rect 2357 10180 2369 10183
rect 2498 10180 2504 10192
rect 2357 10152 2504 10180
rect 2357 10149 2369 10152
rect 2311 10143 2369 10149
rect 2498 10140 2504 10152
rect 2556 10140 2562 10192
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4249 10183 4307 10189
rect 4249 10180 4261 10183
rect 4028 10152 4261 10180
rect 4028 10140 4034 10152
rect 4249 10149 4261 10152
rect 4295 10149 4307 10183
rect 4249 10143 4307 10149
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 5994 10180 6000 10192
rect 4847 10152 6000 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 6178 10189 6184 10192
rect 6175 10180 6184 10189
rect 6139 10152 6184 10180
rect 6175 10143 6184 10152
rect 6178 10140 6184 10143
rect 6236 10140 6242 10192
rect 7101 10183 7159 10189
rect 7101 10149 7113 10183
rect 7147 10180 7159 10183
rect 9861 10183 9919 10189
rect 7147 10152 8156 10180
rect 7147 10149 7159 10152
rect 7101 10143 7159 10149
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10112 5319 10115
rect 5350 10112 5356 10124
rect 5307 10084 5356 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 5350 10072 5356 10084
rect 5408 10112 5414 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 5408 10084 6745 10112
rect 5408 10072 5414 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 7742 10112 7748 10124
rect 7703 10084 7748 10112
rect 6733 10075 6791 10081
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 8128 10121 8156 10152
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 10410 10180 10416 10192
rect 9907 10152 10416 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 12529 10183 12587 10189
rect 12529 10149 12541 10183
rect 12575 10180 12587 10183
rect 13188 10180 13216 10220
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 13872 10220 14381 10248
rect 13872 10208 13878 10220
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 15378 10248 15384 10260
rect 15339 10220 15384 10248
rect 14369 10211 14427 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18656 10220 18797 10248
rect 18656 10208 18662 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 18785 10211 18843 10217
rect 21266 10208 21272 10260
rect 21324 10248 21330 10260
rect 21545 10251 21603 10257
rect 21545 10248 21557 10251
rect 21324 10220 21557 10248
rect 21324 10208 21330 10220
rect 21545 10217 21557 10220
rect 21591 10217 21603 10251
rect 21545 10211 21603 10217
rect 21634 10208 21640 10260
rect 21692 10248 21698 10260
rect 22554 10248 22560 10260
rect 21692 10220 22560 10248
rect 21692 10208 21698 10220
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 23382 10208 23388 10260
rect 23440 10248 23446 10260
rect 23750 10248 23756 10260
rect 23440 10220 23756 10248
rect 23440 10208 23446 10220
rect 23750 10208 23756 10220
rect 23808 10248 23814 10260
rect 24305 10251 24363 10257
rect 24305 10248 24317 10251
rect 23808 10220 24317 10248
rect 23808 10208 23814 10220
rect 24305 10217 24317 10220
rect 24351 10217 24363 10251
rect 24305 10211 24363 10217
rect 12575 10152 13124 10180
rect 13188 10152 15332 10180
rect 12575 10149 12587 10152
rect 12529 10143 12587 10149
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10112 8171 10115
rect 8202 10112 8208 10124
rect 8159 10084 8208 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 12066 10112 12072 10124
rect 11379 10084 12072 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 13096 10112 13124 10152
rect 15304 10124 15332 10152
rect 19886 10140 19892 10192
rect 19944 10180 19950 10192
rect 20162 10180 20168 10192
rect 19944 10152 20168 10180
rect 19944 10140 19950 10152
rect 20162 10140 20168 10152
rect 20220 10140 20226 10192
rect 20530 10140 20536 10192
rect 20588 10140 20594 10192
rect 21910 10180 21916 10192
rect 21871 10152 21916 10180
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 23474 10180 23480 10192
rect 23435 10152 23480 10180
rect 23474 10140 23480 10152
rect 23532 10140 23538 10192
rect 24946 10180 24952 10192
rect 24907 10152 24952 10180
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 25038 10140 25044 10192
rect 25096 10180 25102 10192
rect 25096 10152 25141 10180
rect 25096 10140 25102 10152
rect 13170 10112 13176 10124
rect 13096 10084 13176 10112
rect 13170 10072 13176 10084
rect 13228 10072 13234 10124
rect 13814 10112 13820 10124
rect 13775 10084 13820 10112
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 13976 10115 14034 10121
rect 13976 10081 13988 10115
rect 14022 10112 14034 10115
rect 14090 10112 14096 10124
rect 14022 10084 14096 10112
rect 14022 10081 14034 10084
rect 13976 10075 14034 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 15286 10112 15292 10124
rect 15199 10084 15292 10112
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15620 10084 15761 10112
rect 15620 10072 15626 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 16945 10115 17003 10121
rect 16945 10081 16957 10115
rect 16991 10112 17003 10115
rect 17126 10112 17132 10124
rect 16991 10084 17132 10112
rect 16991 10081 17003 10084
rect 16945 10075 17003 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10081 19855 10115
rect 19978 10112 19984 10124
rect 19939 10084 19984 10112
rect 19797 10075 19855 10081
rect 1946 10044 1952 10056
rect 1907 10016 1952 10044
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4246 10044 4252 10056
rect 4203 10016 4252 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 6178 10044 6184 10056
rect 5859 10016 6184 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 9766 10044 9772 10056
rect 9679 10016 9772 10044
rect 9766 10004 9772 10016
rect 9824 10044 9830 10056
rect 10870 10044 10876 10056
rect 9824 10016 10876 10044
rect 9824 10004 9830 10016
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 11931 10016 12449 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 12437 10013 12449 10016
rect 12483 10044 12495 10047
rect 13446 10044 13452 10056
rect 12483 10016 13452 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 19812 10044 19840 10075
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20548 10056 20576 10140
rect 20162 10044 20168 10056
rect 19812 10016 20168 10044
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 20530 10004 20536 10056
rect 20588 10004 20594 10056
rect 21358 10004 21364 10056
rect 21416 10044 21422 10056
rect 21818 10044 21824 10056
rect 21416 10016 21824 10044
rect 21416 10004 21422 10016
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 23382 10004 23388 10056
rect 23440 10044 23446 10056
rect 23661 10047 23719 10053
rect 23440 10016 23485 10044
rect 23440 10004 23446 10016
rect 23661 10013 23673 10047
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 10318 9976 10324 9988
rect 10279 9948 10324 9976
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 11330 9976 11336 9988
rect 10744 9948 11336 9976
rect 10744 9936 10750 9948
rect 11330 9936 11336 9948
rect 11388 9936 11394 9988
rect 12986 9976 12992 9988
rect 12947 9948 12992 9976
rect 12986 9936 12992 9948
rect 13044 9936 13050 9988
rect 18230 9936 18236 9988
rect 18288 9976 18294 9988
rect 18509 9979 18567 9985
rect 18509 9976 18521 9979
rect 18288 9948 18521 9976
rect 18288 9936 18294 9948
rect 18509 9945 18521 9948
rect 18555 9976 18567 9979
rect 18966 9976 18972 9988
rect 18555 9948 18972 9976
rect 18555 9945 18567 9948
rect 18509 9939 18567 9945
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 22373 9979 22431 9985
rect 22373 9945 22385 9979
rect 22419 9976 22431 9979
rect 23290 9976 23296 9988
rect 22419 9948 23296 9976
rect 22419 9945 22431 9948
rect 22373 9939 22431 9945
rect 23290 9936 23296 9948
rect 23348 9976 23354 9988
rect 23676 9976 23704 10007
rect 25130 10004 25136 10056
rect 25188 10044 25194 10056
rect 25225 10047 25283 10053
rect 25225 10044 25237 10047
rect 25188 10016 25237 10044
rect 25188 10004 25194 10016
rect 25225 10013 25237 10016
rect 25271 10013 25283 10047
rect 25225 10007 25283 10013
rect 23348 9948 23704 9976
rect 23348 9936 23354 9948
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 4154 9908 4160 9920
rect 3660 9880 4160 9908
rect 3660 9868 3666 9880
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 12158 9908 12164 9920
rect 12119 9880 12164 9908
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14047 9911 14105 9917
rect 14047 9908 14059 9911
rect 13872 9880 14059 9908
rect 13872 9868 13878 9880
rect 14047 9877 14059 9880
rect 14093 9877 14105 9911
rect 16390 9908 16396 9920
rect 16351 9880 16396 9908
rect 14047 9871 14105 9877
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 17678 9908 17684 9920
rect 17276 9880 17684 9908
rect 17276 9868 17282 9880
rect 17678 9868 17684 9880
rect 17736 9908 17742 9920
rect 18049 9911 18107 9917
rect 18049 9908 18061 9911
rect 17736 9880 18061 9908
rect 17736 9868 17742 9880
rect 18049 9877 18061 9880
rect 18095 9908 18107 9911
rect 18322 9908 18328 9920
rect 18095 9880 18328 9908
rect 18095 9877 18107 9880
rect 18049 9871 18107 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 20438 9908 20444 9920
rect 20399 9880 20444 9908
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 7742 9704 7748 9716
rect 7340 9676 7748 9704
rect 7340 9664 7346 9676
rect 7742 9664 7748 9676
rect 7800 9664 7806 9716
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 8168 9676 8217 9704
rect 8168 9664 8174 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8205 9667 8263 9673
rect 13909 9707 13967 9713
rect 13909 9673 13921 9707
rect 13955 9704 13967 9707
rect 14090 9704 14096 9716
rect 13955 9676 14096 9704
rect 13955 9673 13967 9676
rect 13909 9667 13967 9673
rect 14090 9664 14096 9676
rect 14148 9664 14154 9716
rect 15286 9704 15292 9716
rect 15247 9676 15292 9704
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 18322 9664 18328 9716
rect 18380 9704 18386 9716
rect 18690 9704 18696 9716
rect 18380 9676 18696 9704
rect 18380 9664 18386 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 21818 9664 21824 9716
rect 21876 9704 21882 9716
rect 23290 9704 23296 9716
rect 21876 9676 23296 9704
rect 21876 9664 21882 9676
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3789 9639 3847 9645
rect 3789 9636 3801 9639
rect 3099 9608 3801 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3789 9605 3801 9608
rect 3835 9636 3847 9639
rect 3970 9636 3976 9648
rect 3835 9608 3976 9636
rect 3835 9605 3847 9608
rect 3789 9599 3847 9605
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 4706 9636 4712 9648
rect 4571 9608 4712 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9568 2191 9571
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 2179 9540 3433 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 3421 9537 3433 9540
rect 3467 9568 3479 9571
rect 3510 9568 3516 9580
rect 3467 9540 3516 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4540 9500 4568 9599
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 7098 9636 7104 9648
rect 6880 9608 7104 9636
rect 6880 9596 6886 9608
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9568 5319 9571
rect 5442 9568 5448 9580
rect 5307 9540 5448 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 5994 9568 6000 9580
rect 5951 9540 6000 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 7006 9528 7012 9580
rect 7064 9528 7070 9580
rect 3927 9472 4568 9500
rect 6641 9503 6699 9509
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 7024 9500 7052 9528
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 6687 9472 7113 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 7101 9469 7113 9472
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 2498 9441 2504 9444
rect 1673 9435 1731 9441
rect 1673 9401 1685 9435
rect 1719 9432 1731 9435
rect 2041 9435 2099 9441
rect 2041 9432 2053 9435
rect 1719 9404 2053 9432
rect 1719 9401 1731 9404
rect 1673 9395 1731 9401
rect 2041 9401 2053 9404
rect 2087 9432 2099 9435
rect 2495 9432 2504 9441
rect 2087 9404 2504 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 2495 9395 2504 9404
rect 2498 9392 2504 9395
rect 2556 9392 2562 9444
rect 5353 9435 5411 9441
rect 5353 9401 5365 9435
rect 5399 9401 5411 9435
rect 7116 9432 7144 9463
rect 7282 9460 7288 9512
rect 7340 9500 7346 9512
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 7340 9472 7389 9500
rect 7340 9460 7346 9472
rect 7377 9469 7389 9472
rect 7423 9500 7435 9503
rect 8128 9500 8156 9664
rect 9214 9636 9220 9648
rect 9175 9608 9220 9636
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 10318 9636 10324 9648
rect 10279 9608 10324 9636
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 10870 9596 10876 9648
rect 10928 9636 10934 9648
rect 11379 9639 11437 9645
rect 11379 9636 11391 9639
rect 10928 9608 11391 9636
rect 10928 9596 10934 9608
rect 11379 9605 11391 9608
rect 11425 9605 11437 9639
rect 11790 9636 11796 9648
rect 11751 9608 11796 9636
rect 11379 9599 11437 9605
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13081 9639 13139 9645
rect 13081 9636 13093 9639
rect 13044 9608 13093 9636
rect 13044 9596 13050 9608
rect 13081 9605 13093 9608
rect 13127 9605 13139 9639
rect 13081 9599 13139 9605
rect 15657 9639 15715 9645
rect 15657 9605 15669 9639
rect 15703 9636 15715 9639
rect 16390 9636 16396 9648
rect 15703 9608 16396 9636
rect 15703 9605 15715 9608
rect 15657 9599 15715 9605
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 19242 9636 19248 9648
rect 17788 9608 19248 9636
rect 7423 9472 8156 9500
rect 8732 9503 8790 9509
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 8732 9469 8744 9503
rect 8778 9500 8790 9503
rect 9232 9500 9260 9596
rect 8778 9472 9260 9500
rect 8778 9469 8790 9472
rect 8732 9463 8790 9469
rect 10410 9460 10416 9512
rect 10468 9500 10474 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 10468 9472 10793 9500
rect 10468 9460 10474 9472
rect 10781 9469 10793 9472
rect 10827 9500 10839 9503
rect 11054 9500 11060 9512
rect 10827 9472 11060 9500
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11308 9503 11366 9509
rect 11308 9469 11320 9503
rect 11354 9500 11366 9503
rect 11808 9500 11836 9596
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 13354 9568 13360 9580
rect 12575 9540 13360 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 13538 9568 13544 9580
rect 13451 9540 13544 9568
rect 13538 9528 13544 9540
rect 13596 9568 13602 9580
rect 13596 9540 14504 9568
rect 13596 9528 13602 9540
rect 14476 9512 14504 9540
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 14884 9540 16037 9568
rect 14884 9528 14890 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17788 9577 17816 9608
rect 18432 9580 18460 9608
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19334 9596 19340 9648
rect 19392 9596 19398 9648
rect 19518 9636 19524 9648
rect 19479 9608 19524 9636
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 20162 9596 20168 9648
rect 20220 9636 20226 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 20220 9608 21373 9636
rect 20220 9596 20226 9608
rect 21361 9605 21373 9608
rect 21407 9636 21419 9639
rect 21729 9639 21787 9645
rect 21729 9636 21741 9639
rect 21407 9608 21741 9636
rect 21407 9605 21419 9608
rect 21361 9599 21419 9605
rect 21729 9605 21741 9608
rect 21775 9636 21787 9639
rect 21910 9636 21916 9648
rect 21775 9608 21916 9636
rect 21775 9605 21787 9608
rect 21729 9599 21787 9605
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 17773 9571 17831 9577
rect 17773 9568 17785 9571
rect 16908 9540 17785 9568
rect 16908 9528 16914 9540
rect 17773 9537 17785 9540
rect 17819 9537 17831 9571
rect 17773 9531 17831 9537
rect 18414 9528 18420 9580
rect 18472 9528 18478 9580
rect 19352 9568 19380 9596
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 19352 9540 19901 9568
rect 19889 9537 19901 9540
rect 19935 9537 19947 9571
rect 20346 9568 20352 9580
rect 20259 9540 20352 9568
rect 19889 9531 19947 9537
rect 20346 9528 20352 9540
rect 20404 9568 20410 9580
rect 20806 9568 20812 9580
rect 20404 9540 20812 9568
rect 20404 9528 20410 9540
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 22572 9568 22600 9676
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 23474 9704 23480 9716
rect 23400 9676 23480 9704
rect 23198 9596 23204 9648
rect 23256 9636 23262 9648
rect 23400 9645 23428 9676
rect 23474 9664 23480 9676
rect 23532 9664 23538 9716
rect 24118 9664 24124 9716
rect 24176 9664 24182 9716
rect 24949 9707 25007 9713
rect 24949 9673 24961 9707
rect 24995 9704 25007 9707
rect 25038 9704 25044 9716
rect 24995 9676 25044 9704
rect 24995 9673 25007 9676
rect 24949 9667 25007 9673
rect 25038 9664 25044 9676
rect 25096 9664 25102 9716
rect 23385 9639 23443 9645
rect 23256 9608 23336 9636
rect 23256 9596 23262 9608
rect 22572 9540 23244 9568
rect 23216 9512 23244 9540
rect 11354 9472 11836 9500
rect 14277 9503 14335 9509
rect 11354 9469 11366 9472
rect 11308 9463 11366 9469
rect 14277 9469 14289 9503
rect 14323 9469 14335 9503
rect 14458 9500 14464 9512
rect 14419 9472 14464 9500
rect 14277 9463 14335 9469
rect 8294 9432 8300 9444
rect 7116 9404 8300 9432
rect 5353 9395 5411 9401
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5368 9364 5396 9395
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 9582 9432 9588 9444
rect 9324 9404 9588 9432
rect 5810 9364 5816 9376
rect 5123 9336 5816 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 6052 9336 6193 9364
rect 6052 9324 6058 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6914 9364 6920 9376
rect 6875 9336 6920 9364
rect 6181 9327 6239 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7834 9364 7840 9376
rect 7795 9336 7840 9364
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8803 9367 8861 9373
rect 8803 9333 8815 9367
rect 8849 9364 8861 9367
rect 9324 9364 9352 9404
rect 9582 9392 9588 9404
rect 9640 9392 9646 9444
rect 9769 9435 9827 9441
rect 9769 9401 9781 9435
rect 9815 9401 9827 9435
rect 9769 9395 9827 9401
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9432 9919 9435
rect 10870 9432 10876 9444
rect 9907 9404 10876 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 9490 9364 9496 9376
rect 8849 9336 9352 9364
rect 9451 9336 9496 9364
rect 8849 9333 8861 9336
rect 8803 9327 8861 9333
rect 9490 9324 9496 9336
rect 9548 9364 9554 9376
rect 9784 9364 9812 9395
rect 10870 9392 10876 9404
rect 10928 9432 10934 9444
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 10928 9404 11161 9432
rect 10928 9392 10934 9404
rect 11149 9401 11161 9404
rect 11195 9432 11207 9435
rect 12158 9432 12164 9444
rect 11195 9404 12164 9432
rect 11195 9401 11207 9404
rect 11149 9395 11207 9401
rect 12158 9392 12164 9404
rect 12216 9432 12222 9444
rect 12621 9435 12679 9441
rect 12621 9432 12633 9435
rect 12216 9404 12633 9432
rect 12216 9392 12222 9404
rect 12621 9401 12633 9404
rect 12667 9401 12679 9435
rect 14292 9432 14320 9463
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15565 9503 15623 9509
rect 15565 9500 15577 9503
rect 15344 9472 15577 9500
rect 15344 9460 15350 9472
rect 15565 9469 15577 9472
rect 15611 9469 15623 9503
rect 15838 9500 15844 9512
rect 15799 9472 15844 9500
rect 15565 9463 15623 9469
rect 14366 9432 14372 9444
rect 14292 9404 14372 9432
rect 12621 9395 12679 9401
rect 14366 9392 14372 9404
rect 14424 9392 14430 9444
rect 15580 9432 15608 9463
rect 15838 9460 15844 9472
rect 15896 9500 15902 9512
rect 16577 9503 16635 9509
rect 16577 9500 16589 9503
rect 15896 9472 16589 9500
rect 15896 9460 15902 9472
rect 16577 9469 16589 9472
rect 16623 9500 16635 9503
rect 17126 9500 17132 9512
rect 16623 9472 17132 9500
rect 16623 9469 16635 9472
rect 16577 9463 16635 9469
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 18230 9500 18236 9512
rect 18191 9472 18236 9500
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18598 9500 18604 9512
rect 18559 9472 18604 9500
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 17037 9435 17095 9441
rect 17037 9432 17049 9435
rect 15580 9404 17049 9432
rect 17037 9401 17049 9404
rect 17083 9432 17095 9435
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 17083 9404 17417 9432
rect 17083 9401 17095 9404
rect 17037 9395 17095 9401
rect 17405 9401 17417 9404
rect 17451 9432 17463 9435
rect 18138 9432 18144 9444
rect 17451 9404 18144 9432
rect 17451 9401 17463 9404
rect 17405 9395 17463 9401
rect 18138 9392 18144 9404
rect 18196 9432 18202 9444
rect 18984 9432 19012 9463
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19337 9503 19395 9509
rect 19337 9500 19349 9503
rect 19300 9472 19349 9500
rect 19300 9460 19306 9472
rect 19337 9469 19349 9472
rect 19383 9469 19395 9503
rect 19337 9463 19395 9469
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 20438 9500 20444 9512
rect 19484 9472 20444 9500
rect 19484 9460 19490 9472
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 22511 9472 22545 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 20806 9441 20812 9444
rect 18196 9404 19012 9432
rect 18196 9392 18202 9404
rect 20803 9395 20812 9441
rect 20864 9432 20870 9444
rect 22373 9435 22431 9441
rect 20864 9404 20903 9432
rect 20806 9392 20812 9395
rect 20864 9392 20870 9404
rect 22373 9401 22385 9435
rect 22419 9432 22431 9435
rect 22480 9432 22508 9463
rect 23198 9460 23204 9512
rect 23256 9460 23262 9512
rect 23308 9432 23336 9608
rect 23385 9605 23397 9639
rect 23431 9605 23443 9639
rect 24136 9636 24164 9664
rect 24302 9636 24308 9648
rect 24136 9608 24308 9636
rect 23385 9599 23443 9605
rect 24302 9596 24308 9608
rect 24360 9596 24366 9648
rect 23750 9568 23756 9580
rect 23711 9540 23756 9568
rect 23750 9528 23756 9540
rect 23808 9528 23814 9580
rect 24118 9528 24124 9580
rect 24176 9568 24182 9580
rect 24397 9571 24455 9577
rect 24397 9568 24409 9571
rect 24176 9540 24409 9568
rect 24176 9528 24182 9540
rect 24397 9537 24409 9540
rect 24443 9568 24455 9571
rect 25130 9568 25136 9580
rect 24443 9540 25136 9568
rect 24443 9537 24455 9540
rect 24397 9531 24455 9537
rect 25130 9528 25136 9540
rect 25188 9528 25194 9580
rect 25222 9500 25228 9512
rect 25183 9472 25228 9500
rect 25222 9460 25228 9472
rect 25280 9500 25286 9512
rect 25777 9503 25835 9509
rect 25777 9500 25789 9503
rect 25280 9472 25789 9500
rect 25280 9460 25286 9472
rect 25777 9469 25789 9472
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 22419 9404 23336 9432
rect 22419 9401 22431 9404
rect 22373 9395 22431 9401
rect 23842 9392 23848 9444
rect 23900 9432 23906 9444
rect 23900 9404 23945 9432
rect 23900 9392 23906 9404
rect 24026 9392 24032 9444
rect 24084 9392 24090 9444
rect 12066 9364 12072 9376
rect 9548 9336 9812 9364
rect 12027 9336 12072 9364
rect 9548 9324 9554 9336
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 14090 9364 14096 9376
rect 14051 9336 14096 9364
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 15930 9364 15936 9376
rect 15252 9336 15936 9364
rect 15252 9324 15258 9336
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 22649 9367 22707 9373
rect 22649 9333 22661 9367
rect 22695 9364 22707 9367
rect 23290 9364 23296 9376
rect 22695 9336 23296 9364
rect 22695 9333 22707 9336
rect 22649 9327 22707 9333
rect 23290 9324 23296 9336
rect 23348 9324 23354 9376
rect 23750 9324 23756 9376
rect 23808 9364 23814 9376
rect 24044 9364 24072 9392
rect 23808 9336 24072 9364
rect 23808 9324 23814 9336
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 25409 9367 25467 9373
rect 25409 9364 25421 9367
rect 24912 9336 25421 9364
rect 24912 9324 24918 9336
rect 25409 9333 25421 9336
rect 25455 9333 25467 9367
rect 25409 9327 25467 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1857 9163 1915 9169
rect 1857 9129 1869 9163
rect 1903 9160 1915 9163
rect 1946 9160 1952 9172
rect 1903 9132 1952 9160
rect 1903 9129 1915 9132
rect 1857 9123 1915 9129
rect 1946 9120 1952 9132
rect 2004 9160 2010 9172
rect 2593 9163 2651 9169
rect 2593 9160 2605 9163
rect 2004 9132 2605 9160
rect 2004 9120 2010 9132
rect 2593 9129 2605 9132
rect 2639 9129 2651 9163
rect 4246 9160 4252 9172
rect 4207 9132 4252 9160
rect 2593 9123 2651 9129
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 5810 9160 5816 9172
rect 5771 9132 5816 9160
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 6178 9160 6184 9172
rect 6091 9132 6184 9160
rect 6178 9120 6184 9132
rect 6236 9160 6242 9172
rect 6914 9160 6920 9172
rect 6236 9132 6920 9160
rect 6236 9120 6242 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7282 9160 7288 9172
rect 7243 9132 7288 9160
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 9766 9160 9772 9172
rect 9539 9132 9772 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 11885 9163 11943 9169
rect 11885 9129 11897 9163
rect 11931 9160 11943 9163
rect 12526 9160 12532 9172
rect 11931 9132 12532 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 12526 9120 12532 9132
rect 12584 9160 12590 9172
rect 13722 9160 13728 9172
rect 12584 9132 13728 9160
rect 12584 9120 12590 9132
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 14240 9132 14381 9160
rect 14240 9120 14246 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 15746 9160 15752 9172
rect 15707 9132 15752 9160
rect 14369 9123 14427 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19797 9163 19855 9169
rect 19797 9160 19809 9163
rect 19392 9132 19809 9160
rect 19392 9120 19398 9132
rect 19797 9129 19809 9132
rect 19843 9129 19855 9163
rect 20162 9160 20168 9172
rect 20123 9132 20168 9160
rect 19797 9123 19855 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 21358 9160 21364 9172
rect 21319 9132 21364 9160
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 23198 9120 23204 9172
rect 23256 9160 23262 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 23256 9132 23305 9160
rect 23256 9120 23262 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 23293 9123 23351 9129
rect 23753 9163 23811 9169
rect 23753 9129 23765 9163
rect 23799 9160 23811 9163
rect 23842 9160 23848 9172
rect 23799 9132 23848 9160
rect 23799 9129 23811 9132
rect 23753 9123 23811 9129
rect 2130 9092 2136 9104
rect 1872 9064 2136 9092
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 1872 9033 1900 9064
rect 2130 9052 2136 9064
rect 2188 9052 2194 9104
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5166 9092 5172 9104
rect 5040 9064 5172 9092
rect 5040 9052 5046 9064
rect 5166 9052 5172 9064
rect 5224 9101 5230 9104
rect 5224 9095 5272 9101
rect 5224 9061 5226 9095
rect 5260 9092 5272 9095
rect 5994 9092 6000 9104
rect 5260 9064 6000 9092
rect 5260 9061 5272 9064
rect 5224 9055 5272 9061
rect 5224 9052 5230 9055
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 6822 9092 6828 9104
rect 6783 9064 6828 9092
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 1857 9027 1915 9033
rect 1857 9024 1869 9027
rect 1728 8996 1869 9024
rect 1728 8984 1734 8996
rect 1857 8993 1869 8996
rect 1903 8993 1915 9027
rect 2038 9024 2044 9036
rect 1999 8996 2044 9024
rect 1857 8987 1915 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 7300 9024 7328 9120
rect 8199 9095 8257 9101
rect 8199 9061 8211 9095
rect 8245 9092 8257 9095
rect 9306 9092 9312 9104
rect 8245 9064 9312 9092
rect 8245 9061 8257 9064
rect 8199 9055 8257 9061
rect 9306 9052 9312 9064
rect 9364 9092 9370 9104
rect 9674 9092 9680 9104
rect 9364 9064 9680 9092
rect 9364 9052 9370 9064
rect 9674 9052 9680 9064
rect 9732 9092 9738 9104
rect 9998 9095 10056 9101
rect 9998 9092 10010 9095
rect 9732 9064 10010 9092
rect 9732 9052 9738 9064
rect 9998 9061 10010 9064
rect 10044 9061 10056 9095
rect 9998 9055 10056 9061
rect 12250 9052 12256 9104
rect 12308 9101 12314 9104
rect 12308 9095 12356 9101
rect 12308 9061 12310 9095
rect 12344 9061 12356 9095
rect 12308 9055 12356 9061
rect 12308 9052 12314 9055
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 13170 9092 13176 9104
rect 12768 9064 13176 9092
rect 12768 9052 12774 9064
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 14458 9052 14464 9104
rect 14516 9092 14522 9104
rect 14737 9095 14795 9101
rect 14737 9092 14749 9095
rect 14516 9064 14749 9092
rect 14516 9052 14522 9064
rect 14737 9061 14749 9064
rect 14783 9092 14795 9095
rect 15654 9092 15660 9104
rect 14783 9064 15660 9092
rect 14783 9061 14795 9064
rect 14737 9055 14795 9061
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 16298 9092 16304 9104
rect 15764 9064 16304 9092
rect 11974 9024 11980 9036
rect 6236 8996 7328 9024
rect 11935 8996 11980 9024
rect 6236 8984 6242 8996
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 14185 9027 14243 9033
rect 14185 8993 14197 9027
rect 14231 9024 14243 9027
rect 14274 9024 14280 9036
rect 14231 8996 14280 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 15764 9024 15792 9064
rect 16298 9052 16304 9064
rect 16356 9092 16362 9104
rect 19352 9092 19380 9120
rect 16356 9064 16620 9092
rect 16356 9052 16362 9064
rect 16592 9036 16620 9064
rect 18248 9064 19380 9092
rect 18248 9036 18276 9064
rect 21726 9052 21732 9104
rect 21784 9101 21790 9104
rect 21784 9095 21832 9101
rect 21784 9061 21786 9095
rect 21820 9061 21832 9095
rect 21784 9055 21832 9061
rect 21784 9052 21790 9055
rect 15930 9024 15936 9036
rect 15151 8996 15792 9024
rect 15891 8996 15936 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16390 9024 16396 9036
rect 16351 8996 16396 9024
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 16574 9024 16580 9036
rect 16487 8996 16580 9024
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 16850 9024 16856 9036
rect 16811 8996 16856 9024
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 18230 9024 18236 9036
rect 18191 8996 18236 9024
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 18782 9024 18788 9036
rect 18743 8996 18788 9024
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 18966 9024 18972 9036
rect 18927 8996 18972 9024
rect 18966 8984 18972 8996
rect 19024 8984 19030 9036
rect 19334 9024 19340 9036
rect 19295 8996 19340 9024
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 22373 9027 22431 9033
rect 22373 8993 22385 9027
rect 22419 9024 22431 9027
rect 23768 9024 23796 9123
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 23934 9120 23940 9172
rect 23992 9160 23998 9172
rect 23992 9132 24256 9160
rect 23992 9120 23998 9132
rect 24118 9092 24124 9104
rect 24079 9064 24124 9092
rect 24118 9052 24124 9064
rect 24176 9052 24182 9104
rect 24228 9101 24256 9132
rect 24946 9120 24952 9172
rect 25004 9160 25010 9172
rect 25041 9163 25099 9169
rect 25041 9160 25053 9163
rect 25004 9132 25053 9160
rect 25004 9120 25010 9132
rect 25041 9129 25053 9132
rect 25087 9129 25099 9163
rect 25041 9123 25099 9129
rect 24213 9095 24271 9101
rect 24213 9061 24225 9095
rect 24259 9061 24271 9095
rect 24213 9055 24271 9061
rect 22419 8996 23796 9024
rect 22419 8993 22431 8996
rect 22373 8987 22431 8993
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 2130 8956 2136 8968
rect 1452 8928 2136 8956
rect 1452 8916 1458 8928
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 4890 8956 4896 8968
rect 4851 8928 4896 8956
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7791 8928 7849 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 7837 8925 7849 8928
rect 7883 8956 7895 8959
rect 8202 8956 8208 8968
rect 7883 8928 8208 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9674 8956 9680 8968
rect 9548 8928 9680 8956
rect 9548 8916 9554 8928
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11146 8956 11152 8968
rect 10744 8928 11152 8956
rect 10744 8916 10750 8928
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13964 8928 14105 8956
rect 13964 8916 13970 8928
rect 14093 8925 14105 8928
rect 14139 8956 14151 8959
rect 14366 8956 14372 8968
rect 14139 8928 14372 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14366 8916 14372 8928
rect 14424 8956 14430 8968
rect 15562 8956 15568 8968
rect 14424 8928 15568 8956
rect 14424 8916 14430 8928
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18800 8956 18828 8984
rect 18003 8928 18828 8956
rect 19521 8959 19579 8965
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 19521 8925 19533 8959
rect 19567 8956 19579 8959
rect 21453 8959 21511 8965
rect 21453 8956 21465 8959
rect 19567 8928 21465 8956
rect 19567 8925 19579 8928
rect 19521 8919 19579 8925
rect 21453 8925 21465 8928
rect 21499 8956 21511 8959
rect 21910 8956 21916 8968
rect 21499 8928 21916 8956
rect 21499 8925 21511 8928
rect 21453 8919 21511 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 24210 8916 24216 8968
rect 24268 8956 24274 8968
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 24268 8928 24409 8956
rect 24268 8916 24274 8928
rect 24397 8925 24409 8928
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 15194 8848 15200 8900
rect 15252 8848 15258 8900
rect 566 8780 572 8832
rect 624 8820 630 8832
rect 7006 8820 7012 8832
rect 624 8792 7012 8820
rect 624 8780 630 8792
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 9674 8820 9680 8832
rect 8803 8792 9680 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 10597 8823 10655 8829
rect 10597 8789 10609 8823
rect 10643 8820 10655 8823
rect 10686 8820 10692 8832
rect 10643 8792 10692 8820
rect 10643 8789 10655 8792
rect 10597 8783 10655 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 12894 8820 12900 8832
rect 12855 8792 12900 8820
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 15212 8820 15240 8848
rect 15378 8820 15384 8832
rect 15212 8792 15384 8820
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15562 8820 15568 8832
rect 15523 8792 15568 8820
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 17862 8820 17868 8832
rect 17635 8792 17868 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 21634 8780 21640 8832
rect 21692 8820 21698 8832
rect 24026 8820 24032 8832
rect 21692 8792 24032 8820
rect 21692 8780 21698 8792
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 2832 8588 3893 8616
rect 2832 8576 2838 8588
rect 3881 8585 3893 8588
rect 3927 8616 3939 8619
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3927 8588 3985 8616
rect 3927 8585 3939 8588
rect 3881 8579 3939 8585
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 3973 8579 4031 8585
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 4948 8588 5549 8616
rect 4948 8576 4954 8588
rect 5537 8585 5549 8588
rect 5583 8585 5595 8619
rect 5537 8579 5595 8585
rect 5552 8548 5580 8579
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6328 8588 6561 8616
rect 6328 8576 6334 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 6549 8579 6607 8585
rect 5718 8548 5724 8560
rect 5552 8520 5724 8548
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 5905 8551 5963 8557
rect 5905 8517 5917 8551
rect 5951 8548 5963 8551
rect 6362 8548 6368 8560
rect 5951 8520 6368 8548
rect 5951 8517 5963 8520
rect 5905 8511 5963 8517
rect 6362 8508 6368 8520
rect 6420 8508 6426 8560
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 3743 8452 4261 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 4249 8449 4261 8452
rect 4295 8480 4307 8483
rect 4338 8480 4344 8492
rect 4295 8452 4344 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 5442 8480 5448 8492
rect 4939 8452 5448 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 2222 8412 2228 8424
rect 1903 8384 2228 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2406 8412 2412 8424
rect 2367 8384 2412 8412
rect 2406 8372 2412 8384
rect 2464 8412 2470 8424
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2464 8384 2973 8412
rect 2464 8372 2470 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 6564 8412 6592 8579
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 9306 8616 9312 8628
rect 9267 8588 9312 8616
rect 9306 8576 9312 8588
rect 9364 8616 9370 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9364 8588 9597 8616
rect 9364 8576 9370 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 9600 8480 9628 8579
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 10652 8588 10701 8616
rect 10652 8576 10658 8588
rect 10689 8585 10701 8588
rect 10735 8616 10747 8619
rect 10870 8616 10876 8628
rect 10735 8588 10876 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 13633 8619 13691 8625
rect 13633 8585 13645 8619
rect 13679 8616 13691 8619
rect 14274 8616 14280 8628
rect 13679 8588 14280 8616
rect 13679 8585 13691 8588
rect 13633 8579 13691 8585
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 19392 8588 20637 8616
rect 19392 8576 19398 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23566 8616 23572 8628
rect 23523 8588 23572 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23566 8576 23572 8588
rect 23624 8576 23630 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25501 8619 25559 8625
rect 25501 8616 25513 8619
rect 25188 8588 25513 8616
rect 25188 8576 25194 8588
rect 25501 8585 25513 8588
rect 25547 8585 25559 8619
rect 25501 8579 25559 8585
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 14185 8551 14243 8557
rect 14185 8548 14197 8551
rect 13872 8520 14197 8548
rect 13872 8508 13878 8520
rect 14185 8517 14197 8520
rect 14231 8548 14243 8551
rect 14458 8548 14464 8560
rect 14231 8520 14464 8548
rect 14231 8517 14243 8520
rect 14185 8511 14243 8517
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 17126 8508 17132 8560
rect 17184 8548 17190 8560
rect 17497 8551 17555 8557
rect 17497 8548 17509 8551
rect 17184 8520 17509 8548
rect 17184 8508 17190 8520
rect 17497 8517 17509 8520
rect 17543 8548 17555 8551
rect 18782 8548 18788 8560
rect 17543 8520 18788 8548
rect 17543 8517 17555 8520
rect 17497 8511 17555 8517
rect 18782 8508 18788 8520
rect 18840 8548 18846 8560
rect 19889 8551 19947 8557
rect 19889 8548 19901 8551
rect 18840 8520 19901 8548
rect 18840 8508 18846 8520
rect 19889 8517 19901 8520
rect 19935 8517 19947 8551
rect 19889 8511 19947 8517
rect 23934 8508 23940 8560
rect 23992 8548 23998 8560
rect 25225 8551 25283 8557
rect 25225 8548 25237 8551
rect 23992 8520 25237 8548
rect 23992 8508 23998 8520
rect 25225 8517 25237 8520
rect 25271 8517 25283 8551
rect 25225 8511 25283 8517
rect 9766 8480 9772 8492
rect 8358 8452 9628 8480
rect 9727 8452 9772 8480
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 5767 8384 6316 8412
rect 6564 8384 6837 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 6288 8356 6316 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7984 8384 8033 8412
rect 7984 8372 7990 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4341 8347 4399 8353
rect 4341 8344 4353 8347
rect 3927 8316 4353 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4341 8313 4353 8316
rect 4387 8313 4399 8347
rect 6270 8344 6276 8356
rect 6231 8316 6276 8344
rect 4341 8307 4399 8313
rect 6270 8304 6276 8316
rect 6328 8304 6334 8356
rect 8358 8353 8386 8452
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9398 8412 9404 8424
rect 8987 8384 9404 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 8343 8347 8401 8353
rect 8343 8313 8355 8347
rect 8389 8344 8401 8347
rect 9600 8344 9628 8452
rect 9766 8440 9772 8452
rect 9824 8480 9830 8492
rect 10965 8483 11023 8489
rect 10965 8480 10977 8483
rect 9824 8452 10977 8480
rect 9824 8440 9830 8452
rect 10965 8449 10977 8452
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11563 8452 11989 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 11977 8449 11989 8452
rect 12023 8480 12035 8483
rect 12250 8480 12256 8492
rect 12023 8452 12256 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12986 8480 12992 8492
rect 12947 8452 12992 8480
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14056 8452 14565 8480
rect 14056 8440 14062 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 16850 8480 16856 8492
rect 14553 8443 14611 8449
rect 15120 8452 16856 8480
rect 11054 8412 11060 8424
rect 9784 8384 11060 8412
rect 9784 8356 9812 8384
rect 11054 8372 11060 8384
rect 11112 8412 11118 8424
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11112 8384 11621 8412
rect 11112 8372 11118 8384
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 14366 8412 14372 8424
rect 14327 8384 14372 8412
rect 14093 8375 14151 8381
rect 8389 8316 8422 8344
rect 9600 8316 9720 8344
rect 8389 8313 8401 8316
rect 8343 8307 8401 8313
rect 2222 8276 2228 8288
rect 2183 8248 2228 8276
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5169 8279 5227 8285
rect 5169 8276 5181 8279
rect 5040 8248 5181 8276
rect 5040 8236 5046 8248
rect 5169 8245 5181 8248
rect 5215 8276 5227 8279
rect 7469 8279 7527 8285
rect 7469 8276 7481 8279
rect 5215 8248 7481 8276
rect 5215 8245 5227 8248
rect 5169 8239 5227 8245
rect 7469 8245 7481 8248
rect 7515 8276 7527 8279
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7515 8248 7849 8276
rect 7515 8245 7527 8248
rect 7469 8239 7527 8245
rect 7837 8245 7849 8248
rect 7883 8276 7895 8279
rect 8357 8276 8385 8307
rect 7883 8248 8385 8276
rect 9692 8276 9720 8316
rect 9766 8304 9772 8356
rect 9824 8304 9830 8356
rect 10090 8347 10148 8353
rect 10090 8344 10102 8347
rect 9876 8316 10102 8344
rect 9876 8276 9904 8316
rect 10090 8313 10102 8316
rect 10136 8344 10148 8347
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 10136 8316 11529 8344
rect 10136 8313 10148 8316
rect 10090 8307 10148 8313
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11624 8344 11652 8375
rect 12621 8347 12679 8353
rect 12621 8344 12633 8347
rect 11624 8316 12633 8344
rect 11517 8307 11575 8313
rect 12621 8313 12633 8316
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 14001 8347 14059 8353
rect 14001 8313 14013 8347
rect 14047 8344 14059 8347
rect 14108 8344 14136 8375
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14826 8372 14832 8424
rect 14884 8412 14890 8424
rect 15120 8421 15148 8452
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 19659 8452 21465 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 21453 8449 21465 8452
rect 21499 8480 21511 8483
rect 22649 8483 22707 8489
rect 22649 8480 22661 8483
rect 21499 8452 22661 8480
rect 21499 8449 21511 8452
rect 21453 8443 21511 8449
rect 22649 8449 22661 8452
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24489 8483 24547 8489
rect 24489 8480 24501 8483
rect 24268 8452 24501 8480
rect 24268 8440 24274 8452
rect 24489 8449 24501 8452
rect 24535 8449 24547 8483
rect 24489 8443 24547 8449
rect 15105 8415 15163 8421
rect 15105 8412 15117 8415
rect 14884 8384 15117 8412
rect 14884 8372 14890 8384
rect 15105 8381 15117 8384
rect 15151 8381 15163 8415
rect 15930 8412 15936 8424
rect 15891 8384 15936 8412
rect 15105 8375 15163 8381
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16390 8412 16396 8424
rect 16351 8384 16396 8412
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 16574 8412 16580 8424
rect 16535 8384 16580 8412
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 16945 8415 17003 8421
rect 16945 8381 16957 8415
rect 16991 8412 17003 8415
rect 18230 8412 18236 8424
rect 16991 8384 17816 8412
rect 18191 8384 18236 8412
rect 16991 8381 17003 8384
rect 16945 8375 17003 8381
rect 15286 8344 15292 8356
rect 14047 8316 15292 8344
rect 14047 8313 14059 8316
rect 14001 8307 14059 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15565 8347 15623 8353
rect 15565 8344 15577 8347
rect 15396 8316 15577 8344
rect 9692 8248 9904 8276
rect 7883 8245 7895 8248
rect 7837 8239 7895 8245
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 15396 8276 15424 8316
rect 15565 8313 15577 8316
rect 15611 8344 15623 8347
rect 16960 8344 16988 8375
rect 17788 8353 17816 8384
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 18782 8412 18788 8424
rect 18743 8384 18788 8412
rect 18782 8372 18788 8384
rect 18840 8372 18846 8424
rect 18966 8412 18972 8424
rect 18879 8384 18972 8412
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19518 8412 19524 8424
rect 19431 8384 19524 8412
rect 19518 8372 19524 8384
rect 19576 8412 19582 8424
rect 19978 8412 19984 8424
rect 19576 8384 19984 8412
rect 19576 8372 19582 8384
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8381 20499 8415
rect 20441 8375 20499 8381
rect 22373 8415 22431 8421
rect 22373 8381 22385 8415
rect 22419 8412 22431 8415
rect 23934 8412 23940 8424
rect 22419 8384 23940 8412
rect 22419 8381 22431 8384
rect 22373 8375 22431 8381
rect 15611 8316 16988 8344
rect 17773 8347 17831 8353
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 17773 8313 17785 8347
rect 17819 8313 17831 8347
rect 17773 8307 17831 8313
rect 12216 8248 15424 8276
rect 15933 8279 15991 8285
rect 12216 8236 12222 8248
rect 15933 8245 15945 8279
rect 15979 8276 15991 8279
rect 16482 8276 16488 8288
rect 15979 8248 16488 8276
rect 15979 8245 15991 8248
rect 15933 8239 15991 8245
rect 16482 8236 16488 8248
rect 16540 8236 16546 8288
rect 17788 8276 17816 8307
rect 17862 8304 17868 8356
rect 17920 8344 17926 8356
rect 18984 8344 19012 8372
rect 20254 8344 20260 8356
rect 17920 8316 19012 8344
rect 20215 8316 20260 8344
rect 17920 8304 17926 8316
rect 20254 8304 20260 8316
rect 20312 8344 20318 8356
rect 20456 8344 20484 8375
rect 23934 8372 23940 8384
rect 23992 8372 23998 8424
rect 21726 8344 21732 8356
rect 20312 8316 20484 8344
rect 21684 8316 21732 8344
rect 20312 8304 20318 8316
rect 21726 8304 21732 8316
rect 21784 8353 21790 8356
rect 21784 8347 21832 8353
rect 21784 8313 21786 8347
rect 21820 8313 21832 8347
rect 21784 8307 21832 8313
rect 21784 8304 21817 8307
rect 23566 8304 23572 8356
rect 23624 8344 23630 8356
rect 24213 8347 24271 8353
rect 24213 8344 24225 8347
rect 23624 8316 24225 8344
rect 23624 8304 23630 8316
rect 24213 8313 24225 8316
rect 24259 8313 24271 8347
rect 24213 8307 24271 8313
rect 24305 8347 24363 8353
rect 24305 8313 24317 8347
rect 24351 8313 24363 8347
rect 24305 8307 24363 8313
rect 18046 8276 18052 8288
rect 17788 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 20806 8236 20812 8288
rect 20864 8276 20870 8288
rect 20901 8279 20959 8285
rect 20901 8276 20913 8279
rect 20864 8248 20913 8276
rect 20864 8236 20870 8248
rect 20901 8245 20913 8248
rect 20947 8276 20959 8279
rect 21269 8279 21327 8285
rect 21269 8276 21281 8279
rect 20947 8248 21281 8276
rect 20947 8245 20959 8248
rect 20901 8239 20959 8245
rect 21269 8245 21281 8248
rect 21315 8276 21327 8279
rect 21789 8276 21817 8304
rect 24026 8276 24032 8288
rect 21315 8248 21817 8276
rect 23987 8248 24032 8276
rect 21315 8245 21327 8248
rect 21269 8239 21327 8245
rect 24026 8236 24032 8248
rect 24084 8276 24090 8288
rect 24320 8276 24348 8307
rect 24084 8248 24348 8276
rect 24084 8236 24090 8248
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1670 8072 1676 8084
rect 1452 8044 1676 8072
rect 1452 8032 1458 8044
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 4154 8072 4160 8084
rect 4115 8044 4160 8072
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 5718 8072 5724 8084
rect 5679 8044 5724 8072
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 7282 8072 7288 8084
rect 7243 8044 7288 8072
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 9490 8072 9496 8084
rect 9451 8044 9496 8072
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 9674 8032 9680 8084
rect 9732 8032 9738 8084
rect 11974 8072 11980 8084
rect 11935 8044 11980 8072
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 12437 8075 12495 8081
rect 12437 8072 12449 8075
rect 12400 8044 12449 8072
rect 12400 8032 12406 8044
rect 12437 8041 12449 8044
rect 12483 8072 12495 8075
rect 12526 8072 12532 8084
rect 12483 8044 12532 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 14001 8075 14059 8081
rect 14001 8072 14013 8075
rect 13688 8044 14013 8072
rect 13688 8032 13694 8044
rect 14001 8041 14013 8044
rect 14047 8072 14059 8075
rect 14090 8072 14096 8084
rect 14047 8044 14096 8072
rect 14047 8041 14059 8044
rect 14001 8035 14059 8041
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 16390 8072 16396 8084
rect 16303 8044 16396 8072
rect 16390 8032 16396 8044
rect 16448 8072 16454 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 16448 8044 17049 8072
rect 16448 8032 16454 8044
rect 17037 8041 17049 8044
rect 17083 8072 17095 8075
rect 17126 8072 17132 8084
rect 17083 8044 17132 8072
rect 17083 8041 17095 8044
rect 17037 8035 17095 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 19426 8072 19432 8084
rect 19387 8044 19432 8072
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 21910 8072 21916 8084
rect 21871 8044 21916 8072
rect 21910 8032 21916 8044
rect 21968 8032 21974 8084
rect 2314 7964 2320 8016
rect 2372 8004 2378 8016
rect 2498 8004 2504 8016
rect 2372 7976 2504 8004
rect 2372 7964 2378 7976
rect 2498 7964 2504 7976
rect 2556 8013 2562 8016
rect 2556 8007 2604 8013
rect 2556 7973 2558 8007
rect 2592 7973 2604 8007
rect 2556 7967 2604 7973
rect 2556 7964 2562 7967
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 7098 8004 7104 8016
rect 6880 7976 7104 8004
rect 6880 7964 6886 7976
rect 7098 7964 7104 7976
rect 7156 8004 7162 8016
rect 9692 8004 9720 8032
rect 9769 8007 9827 8013
rect 9769 8004 9781 8007
rect 7156 7976 7696 8004
rect 9692 7976 9781 8004
rect 7156 7964 7162 7976
rect 2222 7936 2228 7948
rect 2183 7908 2228 7936
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 4154 7936 4160 7948
rect 4115 7908 4160 7936
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 5905 7939 5963 7945
rect 5905 7905 5917 7939
rect 5951 7936 5963 7939
rect 5994 7936 6000 7948
rect 5951 7908 6000 7936
rect 5951 7905 5963 7908
rect 5905 7899 5963 7905
rect 2038 7868 2044 7880
rect 1951 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7868 2102 7880
rect 4540 7868 4568 7899
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6178 7936 6184 7948
rect 6139 7908 6184 7936
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 7668 7945 7696 7976
rect 9769 7973 9781 7976
rect 9815 7973 9827 8007
rect 9769 7967 9827 7973
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 10226 8004 10232 8016
rect 9907 7976 10232 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 10226 7964 10232 7976
rect 10284 8004 10290 8016
rect 12710 8004 12716 8016
rect 10284 7976 12716 8004
rect 10284 7964 10290 7976
rect 12710 7964 12716 7976
rect 12768 7964 12774 8016
rect 12805 8007 12863 8013
rect 12805 7973 12817 8007
rect 12851 8004 12863 8007
rect 12894 8004 12900 8016
rect 12851 7976 12900 8004
rect 12851 7973 12863 7976
rect 12805 7967 12863 7973
rect 12894 7964 12900 7976
rect 12952 8004 12958 8016
rect 13170 8004 13176 8016
rect 12952 7976 13176 8004
rect 12952 7964 12958 7976
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 14366 7964 14372 8016
rect 14424 8004 14430 8016
rect 14737 8007 14795 8013
rect 14737 8004 14749 8007
rect 14424 7976 14749 8004
rect 14424 7964 14430 7976
rect 14737 7973 14749 7976
rect 14783 8004 14795 8007
rect 15105 8007 15163 8013
rect 15105 8004 15117 8007
rect 14783 7976 15117 8004
rect 14783 7973 14795 7976
rect 14737 7967 14795 7973
rect 15105 7973 15117 7976
rect 15151 8004 15163 8007
rect 15151 7976 15608 8004
rect 15151 7973 15163 7976
rect 15105 7967 15163 7973
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 7469 7899 7527 7905
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 7699 7908 8401 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 8389 7905 8401 7908
rect 8435 7936 8447 7939
rect 8846 7936 8852 7948
rect 8435 7908 8852 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 6196 7868 6224 7896
rect 2096 7840 6224 7868
rect 7484 7868 7512 7899
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 11422 7936 11428 7948
rect 11383 7908 11428 7936
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7936 14243 7939
rect 14458 7936 14464 7948
rect 14231 7908 14464 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15580 7945 15608 7976
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 16669 8007 16727 8013
rect 16669 8004 16681 8007
rect 16632 7976 16681 8004
rect 16632 7964 16638 7976
rect 16669 7973 16681 7976
rect 16715 7973 16727 8007
rect 16669 7967 16727 7973
rect 20990 7964 20996 8016
rect 21048 8004 21054 8016
rect 21085 8007 21143 8013
rect 21085 8004 21097 8007
rect 21048 7976 21097 8004
rect 21048 7964 21054 7976
rect 21085 7973 21097 7976
rect 21131 7973 21143 8007
rect 21085 7967 21143 7973
rect 22554 7964 22560 8016
rect 22612 8004 22618 8016
rect 22649 8007 22707 8013
rect 22649 8004 22661 8007
rect 22612 7976 22661 8004
rect 22612 7964 22618 7976
rect 22649 7973 22661 7976
rect 22695 7973 22707 8007
rect 24026 8004 24032 8016
rect 23987 7976 24032 8004
rect 22649 7967 22707 7973
rect 24026 7964 24032 7976
rect 24084 7964 24090 8016
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 15930 7936 15936 7948
rect 15611 7908 15936 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 15930 7896 15936 7908
rect 15988 7896 15994 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16816 7908 16865 7936
rect 16816 7896 16822 7908
rect 16853 7905 16865 7908
rect 16899 7936 16911 7939
rect 16942 7936 16948 7948
rect 16899 7908 16948 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7936 17463 7939
rect 18230 7936 18236 7948
rect 17451 7908 18236 7936
rect 17451 7905 17463 7908
rect 17405 7899 17463 7905
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 18656 7908 18705 7936
rect 18656 7896 18662 7908
rect 18693 7905 18705 7908
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 19061 7939 19119 7945
rect 19061 7905 19073 7939
rect 19107 7905 19119 7939
rect 19518 7936 19524 7948
rect 19479 7908 19524 7936
rect 19061 7899 19119 7905
rect 8110 7868 8116 7880
rect 7484 7840 8116 7868
rect 2096 7828 2102 7840
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 10134 7868 10140 7880
rect 10095 7840 10140 7868
rect 10134 7828 10140 7840
rect 10192 7868 10198 7880
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 10192 7840 10701 7868
rect 10192 7828 10198 7840
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12400 7840 12725 7868
rect 12400 7828 12406 7840
rect 12713 7837 12725 7840
rect 12759 7868 12771 7871
rect 12986 7868 12992 7880
rect 12759 7840 12992 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 15746 7868 15752 7880
rect 15707 7840 15752 7868
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 19076 7868 19104 7899
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22152 7908 22232 7936
rect 22152 7896 22158 7908
rect 18196 7840 19104 7868
rect 20993 7871 21051 7877
rect 18196 7828 18202 7840
rect 20993 7837 21005 7871
rect 21039 7868 21051 7871
rect 21082 7868 21088 7880
rect 21039 7840 21088 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 21082 7828 21088 7840
rect 21140 7828 21146 7880
rect 22204 7868 22232 7908
rect 23934 7896 23940 7948
rect 23992 7936 23998 7948
rect 24121 7939 24179 7945
rect 24121 7936 24133 7939
rect 23992 7908 24133 7936
rect 23992 7896 23998 7908
rect 24121 7905 24133 7908
rect 24167 7905 24179 7939
rect 24121 7899 24179 7905
rect 22557 7871 22615 7877
rect 22557 7868 22569 7871
rect 22204 7840 22569 7868
rect 22557 7837 22569 7840
rect 22603 7868 22615 7871
rect 23290 7868 23296 7880
rect 22603 7840 23296 7868
rect 22603 7837 22615 7840
rect 22557 7831 22615 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 6822 7800 6828 7812
rect 2464 7772 6828 7800
rect 2464 7760 2470 7772
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 11609 7803 11667 7809
rect 11609 7769 11621 7803
rect 11655 7800 11667 7803
rect 12158 7800 12164 7812
rect 11655 7772 12164 7800
rect 11655 7769 11667 7772
rect 11609 7763 11667 7769
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 15381 7803 15439 7809
rect 15381 7769 15393 7803
rect 15427 7800 15439 7803
rect 15654 7800 15660 7812
rect 15427 7772 15660 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 16850 7760 16856 7812
rect 16908 7800 16914 7812
rect 18049 7803 18107 7809
rect 18049 7800 18061 7803
rect 16908 7772 18061 7800
rect 16908 7760 16914 7772
rect 18049 7769 18061 7772
rect 18095 7769 18107 7803
rect 18049 7763 18107 7769
rect 21545 7803 21603 7809
rect 21545 7769 21557 7803
rect 21591 7800 21603 7803
rect 22002 7800 22008 7812
rect 21591 7772 22008 7800
rect 21591 7769 21603 7772
rect 21545 7763 21603 7769
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 23109 7803 23167 7809
rect 23109 7769 23121 7803
rect 23155 7800 23167 7803
rect 23198 7800 23204 7812
rect 23155 7772 23204 7800
rect 23155 7769 23167 7772
rect 23109 7763 23167 7769
rect 23198 7760 23204 7772
rect 23256 7800 23262 7812
rect 24026 7800 24032 7812
rect 23256 7772 24032 7800
rect 23256 7760 23262 7772
rect 24026 7760 24032 7772
rect 24084 7760 24090 7812
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3145 7735 3203 7741
rect 3145 7732 3157 7735
rect 3108 7704 3157 7732
rect 3108 7692 3114 7704
rect 3145 7701 3157 7704
rect 3191 7701 3203 7735
rect 3145 7695 3203 7701
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5534 7732 5540 7744
rect 4856 7704 5540 7732
rect 4856 7692 4862 7704
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 7984 7704 8861 7732
rect 7984 7692 7990 7704
rect 8849 7701 8861 7704
rect 8895 7732 8907 7735
rect 9766 7732 9772 7744
rect 8895 7704 9772 7732
rect 8895 7701 8907 7704
rect 8849 7695 8907 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10410 7692 10416 7744
rect 10468 7732 10474 7744
rect 10686 7732 10692 7744
rect 10468 7704 10692 7732
rect 10468 7692 10474 7704
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 13722 7732 13728 7744
rect 13683 7704 13728 7732
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14369 7735 14427 7741
rect 14369 7701 14381 7735
rect 14415 7732 14427 7735
rect 15838 7732 15844 7744
rect 14415 7704 15844 7732
rect 14415 7701 14427 7704
rect 14369 7695 14427 7701
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 17773 7735 17831 7741
rect 17773 7701 17785 7735
rect 17819 7732 17831 7735
rect 17862 7732 17868 7744
rect 17819 7704 17868 7732
rect 17819 7701 17831 7704
rect 17773 7695 17831 7701
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 20162 7732 20168 7744
rect 20123 7704 20168 7732
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 23750 7692 23756 7744
rect 23808 7732 23814 7744
rect 24118 7732 24124 7744
rect 23808 7704 24124 7732
rect 23808 7692 23814 7704
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 4709 7531 4767 7537
rect 4709 7528 4721 7531
rect 2372 7500 4721 7528
rect 2372 7488 2378 7500
rect 4709 7497 4721 7500
rect 4755 7528 4767 7531
rect 4982 7528 4988 7540
rect 4755 7500 4988 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 6052 7500 6193 7528
rect 6052 7488 6058 7500
rect 6181 7497 6193 7500
rect 6227 7528 6239 7531
rect 6730 7528 6736 7540
rect 6227 7500 6736 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6730 7488 6736 7500
rect 6788 7528 6794 7540
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 6788 7500 7941 7528
rect 6788 7488 6794 7500
rect 7929 7497 7941 7500
rect 7975 7528 7987 7531
rect 8110 7528 8116 7540
rect 7975 7500 8116 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8294 7528 8300 7540
rect 8255 7500 8300 7528
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 9769 7531 9827 7537
rect 9769 7528 9781 7531
rect 9456 7500 9781 7528
rect 9456 7488 9462 7500
rect 9769 7497 9781 7500
rect 9815 7528 9827 7531
rect 10226 7528 10232 7540
rect 9815 7500 10232 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 11422 7528 11428 7540
rect 11383 7500 11428 7528
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12434 7528 12440 7540
rect 12308 7500 12440 7528
rect 12308 7488 12314 7500
rect 12434 7488 12440 7500
rect 12492 7528 12498 7540
rect 12492 7500 12572 7528
rect 12492 7488 12498 7500
rect 2041 7463 2099 7469
rect 2041 7429 2053 7463
rect 2087 7460 2099 7463
rect 2682 7460 2688 7472
rect 2087 7432 2688 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 2056 7324 2084 7423
rect 2682 7420 2688 7432
rect 2740 7420 2746 7472
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 4212 7432 6561 7460
rect 4212 7420 4218 7432
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 10870 7460 10876 7472
rect 10831 7432 10876 7460
rect 6549 7423 6607 7429
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7392 3666 7404
rect 4062 7392 4068 7404
rect 3660 7364 4068 7392
rect 3660 7352 3666 7364
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 1443 7296 2084 7324
rect 6564 7324 6592 7423
rect 10870 7420 10876 7432
rect 10928 7420 10934 7472
rect 12544 7469 12572 7500
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 13262 7528 13268 7540
rect 12860 7500 13268 7528
rect 12860 7488 12866 7500
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 13541 7531 13599 7537
rect 13541 7497 13553 7531
rect 13587 7528 13599 7531
rect 13630 7528 13636 7540
rect 13587 7500 13636 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 15930 7528 15936 7540
rect 15887 7500 15936 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 15930 7488 15936 7500
rect 15988 7528 15994 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 15988 7500 16129 7528
rect 15988 7488 15994 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 18104 7500 18337 7528
rect 18104 7488 18110 7500
rect 18325 7497 18337 7500
rect 18371 7528 18383 7531
rect 19518 7528 19524 7540
rect 18371 7500 19524 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 23992 7500 24685 7528
rect 23992 7488 23998 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 24673 7491 24731 7497
rect 12529 7463 12587 7469
rect 12529 7429 12541 7463
rect 12575 7429 12587 7463
rect 14090 7460 14096 7472
rect 14051 7432 14096 7460
rect 12529 7423 12587 7429
rect 14090 7420 14096 7432
rect 14148 7420 14154 7472
rect 14826 7460 14832 7472
rect 14476 7432 14832 7460
rect 7742 7392 7748 7404
rect 6840 7364 7748 7392
rect 6840 7333 6868 7364
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 10134 7352 10140 7404
rect 10192 7392 10198 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 10192 7364 10333 7392
rect 10192 7352 10198 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 14476 7392 14504 7432
rect 14826 7420 14832 7432
rect 14884 7420 14890 7472
rect 20990 7420 20996 7472
rect 21048 7460 21054 7472
rect 21085 7463 21143 7469
rect 21085 7460 21097 7463
rect 21048 7432 21097 7460
rect 21048 7420 21054 7432
rect 21085 7429 21097 7432
rect 21131 7429 21143 7463
rect 21085 7423 21143 7429
rect 22002 7420 22008 7472
rect 22060 7460 22066 7472
rect 22060 7432 22324 7460
rect 22060 7420 22066 7432
rect 14642 7392 14648 7404
rect 10321 7355 10379 7361
rect 12544 7364 14504 7392
rect 14603 7364 14648 7392
rect 12544 7336 12572 7364
rect 14016 7336 14044 7364
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15344 7364 15485 7392
rect 15344 7352 15350 7364
rect 15473 7361 15485 7364
rect 15519 7392 15531 7395
rect 17862 7392 17868 7404
rect 15519 7364 17868 7392
rect 15519 7361 15531 7364
rect 15473 7355 15531 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 21729 7395 21787 7401
rect 21729 7392 21741 7395
rect 19383 7364 21741 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 21729 7361 21741 7364
rect 21775 7392 21787 7395
rect 22094 7392 22100 7404
rect 21775 7364 22100 7392
rect 21775 7361 21787 7364
rect 21729 7355 21787 7361
rect 22094 7352 22100 7364
rect 22152 7352 22158 7404
rect 22296 7401 22324 7432
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 23474 7352 23480 7404
rect 23532 7392 23538 7404
rect 23750 7392 23756 7404
rect 23532 7364 23756 7392
rect 23532 7352 23538 7364
rect 23750 7352 23756 7364
rect 23808 7352 23814 7404
rect 24026 7392 24032 7404
rect 23987 7364 24032 7392
rect 24026 7352 24032 7364
rect 24084 7352 24090 7404
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6564 7296 6837 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 7156 7296 7297 7324
rect 7156 7284 7162 7296
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 8352 7296 8401 7324
rect 8352 7284 8358 7296
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8846 7324 8852 7336
rect 8807 7296 8852 7324
rect 8389 7287 8447 7293
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12526 7324 12532 7336
rect 12483 7296 12532 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 13998 7324 14004 7336
rect 13911 7296 14004 7324
rect 12713 7287 12771 7293
rect 2958 7256 2964 7268
rect 2919 7228 2964 7256
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3108 7228 3153 7256
rect 3108 7216 3114 7228
rect 4982 7216 4988 7268
rect 5040 7256 5046 7268
rect 5214 7259 5272 7265
rect 5214 7256 5226 7259
rect 5040 7228 5226 7256
rect 5040 7216 5046 7228
rect 5214 7225 5226 7228
rect 5260 7256 5272 7259
rect 5350 7256 5356 7268
rect 5260 7228 5356 7256
rect 5260 7225 5272 7228
rect 5214 7219 5272 7225
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 10137 7259 10195 7265
rect 10137 7225 10149 7259
rect 10183 7256 10195 7259
rect 10410 7256 10416 7268
rect 10183 7228 10416 7256
rect 10183 7225 10195 7228
rect 10137 7219 10195 7225
rect 10410 7216 10416 7228
rect 10468 7216 10474 7268
rect 11885 7259 11943 7265
rect 11885 7225 11897 7259
rect 11931 7256 11943 7259
rect 12728 7256 12756 7287
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 16574 7324 16580 7336
rect 16535 7296 16580 7324
rect 14277 7287 14335 7293
rect 14292 7256 14320 7287
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 19150 7324 19156 7336
rect 19111 7296 19156 7324
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 20162 7324 20168 7336
rect 19484 7296 20168 7324
rect 19484 7284 19490 7296
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 25222 7324 25228 7336
rect 25183 7296 25228 7324
rect 25222 7284 25228 7296
rect 25280 7324 25286 7336
rect 25777 7327 25835 7333
rect 25777 7324 25789 7327
rect 25280 7296 25789 7324
rect 25280 7284 25286 7296
rect 25777 7293 25789 7296
rect 25823 7293 25835 7327
rect 25777 7287 25835 7293
rect 17126 7256 17132 7268
rect 11931 7228 12756 7256
rect 13832 7228 14320 7256
rect 17087 7228 17132 7256
rect 11931 7225 11943 7228
rect 11885 7219 11943 7225
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2314 7188 2320 7200
rect 2096 7160 2320 7188
rect 2096 7148 2102 7160
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 3068 7188 3096 7216
rect 12452 7200 12480 7228
rect 13832 7200 13860 7228
rect 17126 7216 17132 7228
rect 17184 7216 17190 7268
rect 20486 7259 20544 7265
rect 20486 7256 20498 7259
rect 20272 7228 20498 7256
rect 20272 7200 20300 7228
rect 20486 7225 20498 7228
rect 20532 7256 20544 7259
rect 20806 7256 20812 7268
rect 20532 7228 20812 7256
rect 20532 7225 20544 7228
rect 20486 7219 20544 7225
rect 20806 7216 20812 7228
rect 20864 7216 20870 7268
rect 20898 7216 20904 7268
rect 20956 7256 20962 7268
rect 21361 7259 21419 7265
rect 21361 7256 21373 7259
rect 20956 7228 21373 7256
rect 20956 7216 20962 7228
rect 21361 7225 21373 7228
rect 21407 7225 21419 7259
rect 21361 7219 21419 7225
rect 21542 7216 21548 7268
rect 21600 7256 21606 7268
rect 22002 7256 22008 7268
rect 21600 7228 22008 7256
rect 21600 7216 21606 7228
rect 22002 7216 22008 7228
rect 22060 7216 22066 7268
rect 22094 7216 22100 7268
rect 22152 7256 22158 7268
rect 23474 7256 23480 7268
rect 22152 7228 22197 7256
rect 23435 7228 23480 7256
rect 22152 7216 22158 7228
rect 23474 7216 23480 7228
rect 23532 7216 23538 7268
rect 23845 7259 23903 7265
rect 23845 7225 23857 7259
rect 23891 7225 23903 7259
rect 23845 7219 23903 7225
rect 4154 7188 4160 7200
rect 2823 7160 3096 7188
rect 4115 7160 4160 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5592 7160 5825 7188
rect 5592 7148 5598 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 6914 7188 6920 7200
rect 6875 7160 6920 7188
rect 5813 7151 5871 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 8478 7188 8484 7200
rect 8439 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 12250 7188 12256 7200
rect 12211 7160 12256 7188
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 12434 7148 12440 7200
rect 12492 7148 12498 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13814 7188 13820 7200
rect 13775 7160 13820 7188
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 15105 7191 15163 7197
rect 15105 7188 15117 7191
rect 14516 7160 15117 7188
rect 14516 7148 14522 7160
rect 15105 7157 15117 7160
rect 15151 7188 15163 7191
rect 15194 7188 15200 7200
rect 15151 7160 15200 7188
rect 15151 7157 15163 7160
rect 15105 7151 15163 7157
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 16816 7160 17417 7188
rect 16816 7148 16822 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17405 7151 17463 7157
rect 17865 7191 17923 7197
rect 17865 7157 17877 7191
rect 17911 7188 17923 7191
rect 18138 7188 18144 7200
rect 17911 7160 18144 7188
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 18138 7148 18144 7160
rect 18196 7148 18202 7200
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 18656 7160 19625 7188
rect 18656 7148 18662 7160
rect 19613 7157 19625 7160
rect 19659 7157 19671 7191
rect 19613 7151 19671 7157
rect 20073 7191 20131 7197
rect 20073 7157 20085 7191
rect 20119 7188 20131 7191
rect 20254 7188 20260 7200
rect 20119 7160 20260 7188
rect 20119 7157 20131 7160
rect 20073 7151 20131 7157
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 20990 7148 20996 7200
rect 21048 7188 21054 7200
rect 22554 7188 22560 7200
rect 21048 7160 22560 7188
rect 21048 7148 21054 7160
rect 22554 7148 22560 7160
rect 22612 7188 22618 7200
rect 22925 7191 22983 7197
rect 22925 7188 22937 7191
rect 22612 7160 22937 7188
rect 22612 7148 22618 7160
rect 22925 7157 22937 7160
rect 22971 7157 22983 7191
rect 23492 7188 23520 7216
rect 23860 7188 23888 7219
rect 25406 7188 25412 7200
rect 23492 7160 23888 7188
rect 25367 7160 25412 7188
rect 22925 7151 22983 7157
rect 25406 7148 25412 7160
rect 25464 7148 25470 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2041 6987 2099 6993
rect 2041 6953 2053 6987
rect 2087 6984 2099 6987
rect 2222 6984 2228 6996
rect 2087 6956 2228 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 3881 6987 3939 6993
rect 3881 6953 3893 6987
rect 3927 6984 3939 6987
rect 3927 6956 4844 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 2314 6916 2320 6928
rect 2275 6888 2320 6916
rect 2314 6876 2320 6888
rect 2372 6876 2378 6928
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4249 6919 4307 6925
rect 4249 6916 4261 6919
rect 4212 6888 4261 6916
rect 4212 6876 4218 6888
rect 4249 6885 4261 6888
rect 4295 6885 4307 6919
rect 4816 6916 4844 6956
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 5077 6987 5135 6993
rect 5077 6984 5089 6987
rect 4948 6956 5089 6984
rect 4948 6944 4954 6956
rect 5077 6953 5089 6956
rect 5123 6953 5135 6987
rect 5077 6947 5135 6953
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 6178 6984 6184 6996
rect 5675 6956 6184 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5644 6916 5672 6947
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 6880 6956 6929 6984
rect 6880 6944 6886 6956
rect 6917 6953 6929 6956
rect 6963 6984 6975 6987
rect 7098 6984 7104 6996
rect 6963 6956 7104 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7098 6944 7104 6956
rect 7156 6984 7162 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 7156 6956 7297 6984
rect 7156 6944 7162 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 9766 6984 9772 6996
rect 9727 6956 9772 6984
rect 7285 6947 7343 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 13170 6984 13176 6996
rect 13131 6956 13176 6984
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 13998 6984 14004 6996
rect 13959 6956 14004 6984
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 16942 6984 16948 6996
rect 15028 6956 16436 6984
rect 16903 6956 16948 6984
rect 4816 6888 5672 6916
rect 6042 6919 6100 6925
rect 4249 6879 4307 6885
rect 6042 6885 6054 6919
rect 6088 6885 6100 6919
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 6042 6879 6100 6885
rect 7392 6888 7665 6916
rect 5718 6848 5724 6860
rect 5679 6820 5724 6848
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 1912 6752 2237 6780
rect 1912 6740 1918 6752
rect 2225 6749 2237 6752
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 2958 6780 2964 6792
rect 2915 6752 2964 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 2958 6740 2964 6752
rect 3016 6780 3022 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 3016 6752 3157 6780
rect 3016 6740 3022 6752
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 3510 6672 3516 6724
rect 3568 6712 3574 6724
rect 4172 6712 4200 6743
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 4396 6752 4445 6780
rect 4396 6740 4402 6752
rect 4433 6749 4445 6752
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 6057 6780 6085 6879
rect 7392 6860 7420 6888
rect 7653 6885 7665 6888
rect 7699 6885 7711 6919
rect 7653 6879 7711 6885
rect 13725 6919 13783 6925
rect 13725 6885 13737 6919
rect 13771 6916 13783 6919
rect 15028 6916 15056 6956
rect 15286 6916 15292 6928
rect 13771 6888 15056 6916
rect 15120 6888 15292 6916
rect 13771 6885 13783 6888
rect 13725 6879 13783 6885
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6848 6699 6851
rect 7374 6848 7380 6860
rect 6687 6820 7380 6848
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9582 6848 9588 6860
rect 9539 6820 9588 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 9953 6851 10011 6857
rect 9953 6817 9965 6851
rect 9999 6848 10011 6851
rect 10042 6848 10048 6860
rect 9999 6820 10048 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6817 10195 6851
rect 12158 6848 12164 6860
rect 12119 6820 12164 6848
rect 10137 6811 10195 6817
rect 5408 6752 6085 6780
rect 5408 6740 5414 6752
rect 7282 6740 7288 6792
rect 7340 6780 7346 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7340 6752 7573 6780
rect 7340 6740 7346 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7561 6743 7619 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 10152 6780 10180 6811
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 14182 6848 14188 6860
rect 12492 6820 12537 6848
rect 14143 6820 14188 6848
rect 12492 6808 12498 6820
rect 14182 6808 14188 6820
rect 14240 6848 14246 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 14240 6820 14657 6848
rect 14240 6808 14246 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 15120 6848 15148 6888
rect 15286 6876 15292 6888
rect 15344 6876 15350 6928
rect 16408 6916 16436 6956
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17405 6987 17463 6993
rect 17405 6953 17417 6987
rect 17451 6984 17463 6987
rect 18322 6984 18328 6996
rect 17451 6956 18328 6984
rect 17451 6953 17463 6956
rect 17405 6947 17463 6953
rect 17420 6916 17448 6947
rect 18322 6944 18328 6956
rect 18380 6984 18386 6996
rect 20717 6987 20775 6993
rect 18380 6956 19104 6984
rect 18380 6944 18386 6956
rect 16408 6888 17448 6916
rect 15838 6848 15844 6860
rect 14645 6811 14703 6817
rect 15028 6820 15148 6848
rect 15799 6820 15844 6848
rect 9364 6752 10180 6780
rect 11701 6783 11759 6789
rect 9364 6740 9370 6752
rect 11701 6749 11713 6783
rect 11747 6780 11759 6783
rect 12342 6780 12348 6792
rect 11747 6752 12348 6780
rect 11747 6749 11759 6752
rect 11701 6743 11759 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12618 6780 12624 6792
rect 12579 6752 12624 6780
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 5258 6712 5264 6724
rect 3568 6684 5264 6712
rect 3568 6672 3574 6684
rect 5258 6672 5264 6684
rect 5316 6672 5322 6724
rect 12250 6712 12256 6724
rect 10888 6684 12256 6712
rect 10888 6656 10916 6684
rect 12250 6672 12256 6684
rect 12308 6712 12314 6724
rect 12526 6712 12532 6724
rect 12308 6684 12532 6712
rect 12308 6672 12314 6684
rect 12526 6672 12532 6684
rect 12584 6672 12590 6724
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6712 14427 6715
rect 15028 6712 15056 6820
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6817 16083 6851
rect 16025 6811 16083 6817
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6780 15163 6783
rect 15654 6780 15660 6792
rect 15151 6752 15660 6780
rect 15151 6749 15163 6752
rect 15105 6743 15163 6749
rect 15654 6740 15660 6752
rect 15712 6780 15718 6792
rect 16040 6780 16068 6811
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 16577 6851 16635 6857
rect 16577 6848 16589 6851
rect 16448 6820 16589 6848
rect 16448 6808 16454 6820
rect 16577 6817 16589 6820
rect 16623 6848 16635 6851
rect 16666 6848 16672 6860
rect 16623 6820 16672 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 16868 6857 16896 6888
rect 16853 6851 16911 6857
rect 16853 6817 16865 6851
rect 16899 6817 16911 6851
rect 16853 6811 16911 6817
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 18230 6848 18236 6860
rect 18187 6820 18236 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 18598 6848 18604 6860
rect 18559 6820 18604 6848
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18693 6851 18751 6857
rect 18693 6817 18705 6851
rect 18739 6817 18751 6851
rect 18693 6811 18751 6817
rect 15712 6752 16068 6780
rect 15712 6740 15718 6752
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 18708 6780 18736 6811
rect 18966 6808 18972 6860
rect 19024 6848 19030 6860
rect 19076 6857 19104 6956
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 21082 6984 21088 6996
rect 20763 6956 21088 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 21082 6944 21088 6956
rect 21140 6944 21146 6996
rect 21634 6984 21640 6996
rect 21595 6956 21640 6984
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22002 6984 22008 6996
rect 21963 6956 22008 6984
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 23290 6984 23296 6996
rect 23251 6956 23296 6984
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 23750 6984 23756 6996
rect 23711 6956 23756 6984
rect 23750 6944 23756 6956
rect 23808 6944 23814 6996
rect 19061 6851 19119 6857
rect 19061 6848 19073 6851
rect 19024 6820 19073 6848
rect 19024 6808 19030 6820
rect 19061 6817 19073 6820
rect 19107 6817 19119 6851
rect 19061 6811 19119 6817
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 19981 6851 20039 6857
rect 19981 6848 19993 6851
rect 19392 6820 19993 6848
rect 19392 6808 19398 6820
rect 19981 6817 19993 6820
rect 20027 6848 20039 6851
rect 20898 6848 20904 6860
rect 20027 6820 20904 6848
rect 20027 6817 20039 6820
rect 19981 6811 20039 6817
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 21652 6848 21680 6944
rect 22462 6925 22468 6928
rect 22459 6916 22468 6925
rect 22423 6888 22468 6916
rect 22459 6879 22468 6888
rect 22462 6876 22468 6879
rect 22520 6876 22526 6928
rect 24121 6919 24179 6925
rect 24121 6885 24133 6919
rect 24167 6916 24179 6919
rect 24210 6916 24216 6928
rect 24167 6888 24216 6916
rect 24167 6885 24179 6888
rect 24121 6879 24179 6885
rect 24210 6876 24216 6888
rect 24268 6876 24274 6928
rect 21039 6820 21680 6848
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 21726 6808 21732 6860
rect 21784 6848 21790 6860
rect 22097 6851 22155 6857
rect 22097 6848 22109 6851
rect 21784 6820 22109 6848
rect 21784 6808 21790 6820
rect 22097 6817 22109 6820
rect 22143 6817 22155 6851
rect 22097 6811 22155 6817
rect 18874 6780 18880 6792
rect 17644 6752 18880 6780
rect 17644 6740 17650 6752
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6780 24087 6783
rect 24118 6780 24124 6792
rect 24075 6752 24124 6780
rect 24075 6749 24087 6752
rect 24029 6743 24087 6749
rect 24118 6740 24124 6752
rect 24176 6740 24182 6792
rect 24673 6783 24731 6789
rect 24673 6749 24685 6783
rect 24719 6780 24731 6783
rect 25038 6780 25044 6792
rect 24719 6752 25044 6780
rect 24719 6749 24731 6752
rect 24673 6743 24731 6749
rect 25038 6740 25044 6752
rect 25096 6740 25102 6792
rect 19242 6712 19248 6724
rect 14415 6684 15056 6712
rect 19203 6684 19248 6712
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 19242 6672 19248 6684
rect 19300 6672 19306 6724
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1544 6616 1593 6644
rect 1544 6604 1550 6616
rect 1581 6613 1593 6616
rect 1627 6644 1639 6647
rect 1946 6644 1952 6656
rect 1627 6616 1952 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 6638 6644 6644 6656
rect 4764 6616 6644 6644
rect 4764 6604 4770 6616
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 10870 6644 10876 6656
rect 10831 6616 10876 6644
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6644 12127 6647
rect 12434 6644 12440 6656
rect 12115 6616 12440 6644
rect 12115 6613 12127 6616
rect 12069 6607 12127 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 17402 6604 17408 6656
rect 17460 6644 17466 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17460 6616 17693 6644
rect 17460 6604 17466 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17681 6607 17739 6613
rect 18230 6604 18236 6656
rect 18288 6644 18294 6656
rect 19426 6644 19432 6656
rect 18288 6616 19432 6644
rect 18288 6604 18294 6616
rect 19426 6604 19432 6616
rect 19484 6644 19490 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 19484 6616 19625 6644
rect 19484 6604 19490 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 21174 6644 21180 6656
rect 21135 6616 21180 6644
rect 19613 6607 19671 6613
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 23017 6647 23075 6653
rect 23017 6613 23029 6647
rect 23063 6644 23075 6647
rect 24210 6644 24216 6656
rect 23063 6616 24216 6644
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 24210 6604 24216 6616
rect 24268 6604 24274 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4246 6440 4252 6452
rect 4207 6412 4252 6440
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 6914 6440 6920 6452
rect 4816 6412 6920 6440
rect 3605 6375 3663 6381
rect 3605 6341 3617 6375
rect 3651 6372 3663 6375
rect 4816 6372 4844 6412
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7432 6412 7849 6440
rect 7432 6400 7438 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 10042 6440 10048 6452
rect 9955 6412 10048 6440
rect 7837 6403 7895 6409
rect 10042 6400 10048 6412
rect 10100 6440 10106 6452
rect 10100 6412 11008 6440
rect 10100 6400 10106 6412
rect 3651 6344 4844 6372
rect 3651 6341 3663 6344
rect 3605 6335 3663 6341
rect 3620 6304 3648 6335
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 5408 6344 6193 6372
rect 5408 6332 5414 6344
rect 6181 6341 6193 6344
rect 6227 6372 6239 6375
rect 8662 6372 8668 6384
rect 6227 6344 8668 6372
rect 6227 6341 6239 6344
rect 6181 6335 6239 6341
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 10870 6372 10876 6384
rect 10831 6344 10876 6372
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 10980 6372 11008 6412
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 12216 6412 13461 6440
rect 12216 6400 12222 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13906 6440 13912 6452
rect 13867 6412 13912 6440
rect 13449 6403 13507 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17586 6440 17592 6452
rect 17543 6412 17592 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 13924 6372 13952 6400
rect 16206 6372 16212 6384
rect 10980 6344 13952 6372
rect 15580 6344 16212 6372
rect 5718 6304 5724 6316
rect 3160 6276 3648 6304
rect 5679 6276 5724 6304
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 3160 6236 3188 6276
rect 5718 6264 5724 6276
rect 5776 6304 5782 6316
rect 7834 6304 7840 6316
rect 5776 6276 7840 6304
rect 5776 6264 5782 6276
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 11238 6304 11244 6316
rect 11199 6276 11244 6304
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 11931 6276 12572 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12544 6248 12572 6276
rect 2363 6208 3188 6236
rect 3237 6239 3295 6245
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 3694 6236 3700 6248
rect 3283 6208 3700 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4706 6236 4712 6248
rect 4111 6208 4712 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6564 6208 6837 6236
rect 2038 6128 2044 6180
rect 2096 6168 2102 6180
rect 2133 6171 2191 6177
rect 2133 6168 2145 6171
rect 2096 6140 2145 6168
rect 2096 6128 2102 6140
rect 2133 6137 2145 6140
rect 2179 6168 2191 6171
rect 2638 6171 2696 6177
rect 2638 6168 2650 6171
rect 2179 6140 2650 6168
rect 2179 6137 2191 6140
rect 2133 6131 2191 6137
rect 2638 6137 2650 6140
rect 2684 6137 2696 6171
rect 5258 6168 5264 6180
rect 5219 6140 5264 6168
rect 2638 6131 2696 6137
rect 5258 6128 5264 6140
rect 5316 6128 5322 6180
rect 5353 6171 5411 6177
rect 5353 6137 5365 6171
rect 5399 6168 5411 6171
rect 5442 6168 5448 6180
rect 5399 6140 5448 6168
rect 5399 6137 5411 6140
rect 5353 6131 5411 6137
rect 1857 6103 1915 6109
rect 1857 6069 1869 6103
rect 1903 6100 1915 6103
rect 2314 6100 2320 6112
rect 1903 6072 2320 6100
rect 1903 6069 1915 6072
rect 1857 6063 1915 6069
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 3973 6103 4031 6109
rect 3973 6069 3985 6103
rect 4019 6100 4031 6103
rect 4154 6100 4160 6112
rect 4019 6072 4160 6100
rect 4019 6069 4031 6072
rect 3973 6063 4031 6069
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5368 6100 5396 6131
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 6564 6112 6592 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7156 6208 7297 6236
rect 7156 6196 7162 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 8754 6236 8760 6248
rect 8715 6208 8760 6236
rect 7285 6199 7343 6205
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6236 10839 6239
rect 11054 6236 11060 6248
rect 10827 6208 10861 6236
rect 10967 6208 11060 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 9119 6171 9177 6177
rect 9119 6137 9131 6171
rect 9165 6137 9177 6171
rect 9119 6131 9177 6137
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 10796 6168 10824 6199
rect 11054 6196 11060 6208
rect 11112 6236 11118 6248
rect 11112 6208 12296 6236
rect 11112 6196 11118 6208
rect 11698 6168 11704 6180
rect 10735 6140 11704 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 6546 6100 6552 6112
rect 5123 6072 5396 6100
rect 6507 6072 6552 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 6914 6100 6920 6112
rect 6875 6072 6920 6100
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 7340 6072 8217 6100
rect 7340 6060 7346 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8662 6100 8668 6112
rect 8623 6072 8668 6100
rect 8205 6063 8263 6069
rect 8662 6060 8668 6072
rect 8720 6100 8726 6112
rect 9140 6100 9168 6131
rect 11698 6128 11704 6140
rect 11756 6168 11762 6180
rect 11974 6168 11980 6180
rect 11756 6140 11980 6168
rect 11756 6128 11762 6140
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 12268 6168 12296 6208
rect 12342 6196 12348 6248
rect 12400 6236 12406 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12400 6208 12449 6236
rect 12400 6196 12406 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 12526 6196 12532 6248
rect 12584 6236 12590 6248
rect 12713 6239 12771 6245
rect 12584 6208 12629 6236
rect 12584 6196 12590 6208
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 13814 6236 13820 6248
rect 12759 6208 13820 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 12728 6168 12756 6199
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 13906 6196 13912 6248
rect 13964 6236 13970 6248
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13964 6208 14013 6236
rect 13964 6196 13970 6208
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14550 6236 14556 6248
rect 14511 6208 14556 6236
rect 14001 6199 14059 6205
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 15580 6245 15608 6344
rect 16206 6332 16212 6344
rect 16264 6372 16270 6384
rect 16669 6375 16727 6381
rect 16669 6372 16681 6375
rect 16264 6344 16681 6372
rect 16264 6332 16270 6344
rect 16669 6341 16681 6344
rect 16715 6372 16727 6375
rect 17512 6372 17540 6403
rect 17586 6400 17592 6412
rect 17644 6440 17650 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17644 6412 17785 6440
rect 17644 6400 17650 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 17773 6403 17831 6409
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 20956 6412 21281 6440
rect 20956 6400 20962 6412
rect 21269 6409 21281 6412
rect 21315 6409 21327 6443
rect 21726 6440 21732 6452
rect 21687 6412 21732 6440
rect 21269 6403 21327 6409
rect 21726 6400 21732 6412
rect 21784 6400 21790 6452
rect 22649 6443 22707 6449
rect 22649 6409 22661 6443
rect 22695 6440 22707 6443
rect 23382 6440 23388 6452
rect 22695 6412 23388 6440
rect 22695 6409 22707 6412
rect 22649 6403 22707 6409
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 24118 6440 24124 6452
rect 23523 6412 24124 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 24118 6400 24124 6412
rect 24176 6400 24182 6452
rect 25314 6440 25320 6452
rect 25275 6412 25320 6440
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 16715 6344 17540 6372
rect 16715 6341 16727 6344
rect 16669 6335 16727 6341
rect 16298 6304 16304 6316
rect 16259 6276 16304 6304
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 19797 6307 19855 6313
rect 19797 6304 19809 6307
rect 18616 6276 19809 6304
rect 18616 6248 18644 6276
rect 19797 6273 19809 6276
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 24397 6307 24455 6313
rect 24397 6273 24409 6307
rect 24443 6304 24455 6307
rect 25332 6304 25360 6400
rect 24443 6276 25360 6304
rect 24443 6273 24455 6276
rect 24397 6267 24455 6273
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 15657 6239 15715 6245
rect 15657 6205 15669 6239
rect 15703 6236 15715 6239
rect 15746 6236 15752 6248
rect 15703 6208 15752 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 17494 6236 17500 6248
rect 15887 6208 17500 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 12268 6140 12756 6168
rect 15105 6171 15163 6177
rect 12268 6112 12296 6140
rect 15105 6137 15117 6171
rect 15151 6168 15163 6171
rect 15286 6168 15292 6180
rect 15151 6140 15292 6168
rect 15151 6137 15163 6140
rect 15105 6131 15163 6137
rect 15286 6128 15292 6140
rect 15344 6168 15350 6180
rect 15856 6168 15884 6199
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 18230 6236 18236 6248
rect 18191 6208 18236 6236
rect 18230 6196 18236 6208
rect 18288 6196 18294 6248
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6236 18567 6239
rect 18598 6236 18604 6248
rect 18555 6208 18604 6236
rect 18555 6205 18567 6208
rect 18509 6199 18567 6205
rect 15344 6140 15884 6168
rect 15344 6128 15350 6140
rect 17402 6128 17408 6180
rect 17460 6168 17466 6180
rect 18524 6168 18552 6199
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 18874 6236 18880 6248
rect 18835 6208 18880 6236
rect 18874 6196 18880 6208
rect 18932 6196 18938 6248
rect 19058 6196 19064 6248
rect 19116 6236 19122 6248
rect 19337 6239 19395 6245
rect 19337 6236 19349 6239
rect 19116 6208 19349 6236
rect 19116 6196 19122 6208
rect 19337 6205 19349 6208
rect 19383 6205 19395 6239
rect 20346 6236 20352 6248
rect 20307 6208 20352 6236
rect 19337 6199 19395 6205
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 21266 6196 21272 6248
rect 21324 6236 21330 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 21324 6208 22477 6236
rect 21324 6196 21330 6208
rect 22465 6205 22477 6208
rect 22511 6236 22523 6239
rect 23017 6239 23075 6245
rect 23017 6236 23029 6239
rect 22511 6208 23029 6236
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 23017 6205 23029 6208
rect 23063 6205 23075 6239
rect 23017 6199 23075 6205
rect 17460 6140 18552 6168
rect 20711 6171 20769 6177
rect 17460 6128 17466 6140
rect 20711 6137 20723 6171
rect 20757 6168 20769 6171
rect 24489 6171 24547 6177
rect 20757 6140 20791 6168
rect 20757 6137 20769 6140
rect 20711 6131 20769 6137
rect 24489 6137 24501 6171
rect 24535 6137 24547 6171
rect 25038 6168 25044 6180
rect 24999 6140 25044 6168
rect 24489 6131 24547 6137
rect 8720 6072 9168 6100
rect 9677 6103 9735 6109
rect 8720 6060 8726 6072
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 9858 6100 9864 6112
rect 9723 6072 9864 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 12250 6100 12256 6112
rect 12211 6072 12256 6100
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12894 6100 12900 6112
rect 12855 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 14090 6100 14096 6112
rect 14051 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 15473 6103 15531 6109
rect 15473 6069 15485 6103
rect 15519 6100 15531 6103
rect 15746 6100 15752 6112
rect 15519 6072 15752 6100
rect 15519 6069 15531 6072
rect 15473 6063 15531 6069
rect 15746 6060 15752 6072
rect 15804 6100 15810 6112
rect 16758 6100 16764 6112
rect 15804 6072 16764 6100
rect 15804 6060 15810 6072
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 17037 6103 17095 6109
rect 17037 6069 17049 6103
rect 17083 6100 17095 6103
rect 17678 6100 17684 6112
rect 17083 6072 17684 6100
rect 17083 6069 17095 6072
rect 17037 6063 17095 6069
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 19242 6100 19248 6112
rect 19203 6072 19248 6100
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 20254 6100 20260 6112
rect 20167 6072 20260 6100
rect 20254 6060 20260 6072
rect 20312 6100 20318 6112
rect 20726 6100 20754 6131
rect 20898 6100 20904 6112
rect 20312 6072 20904 6100
rect 20312 6060 20318 6072
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 22189 6103 22247 6109
rect 22189 6069 22201 6103
rect 22235 6100 22247 6103
rect 22370 6100 22376 6112
rect 22235 6072 22376 6100
rect 22235 6069 22247 6072
rect 22189 6063 22247 6069
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 24026 6060 24032 6112
rect 24084 6100 24090 6112
rect 24121 6103 24179 6109
rect 24121 6100 24133 6103
rect 24084 6072 24133 6100
rect 24084 6060 24090 6072
rect 24121 6069 24133 6072
rect 24167 6100 24179 6103
rect 24504 6100 24532 6131
rect 25038 6128 25044 6140
rect 25096 6128 25102 6180
rect 24167 6072 24532 6100
rect 24167 6069 24179 6072
rect 24121 6063 24179 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1854 5896 1860 5908
rect 1815 5868 1860 5896
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 4154 5896 4160 5908
rect 2915 5868 4160 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 2038 5788 2044 5840
rect 2096 5828 2102 5840
rect 2270 5831 2328 5837
rect 2270 5828 2282 5831
rect 2096 5800 2282 5828
rect 2096 5788 2102 5800
rect 2270 5797 2282 5800
rect 2316 5797 2328 5831
rect 2270 5791 2328 5797
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1762 5760 1768 5772
rect 1636 5732 1768 5760
rect 1636 5720 1642 5732
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 1946 5692 1952 5704
rect 1907 5664 1952 5692
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 2884 5692 2912 5859
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 5813 5899 5871 5905
rect 5813 5865 5825 5899
rect 5859 5896 5871 5899
rect 5994 5896 6000 5908
rect 5859 5868 6000 5896
rect 5859 5865 5871 5868
rect 5813 5859 5871 5865
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5896 7343 5899
rect 7558 5896 7564 5908
rect 7331 5868 7564 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 9306 5896 9312 5908
rect 7708 5868 9312 5896
rect 7708 5856 7714 5868
rect 9306 5856 9312 5868
rect 9364 5896 9370 5908
rect 9401 5899 9459 5905
rect 9401 5896 9413 5899
rect 9364 5868 9413 5896
rect 9364 5856 9370 5868
rect 9401 5865 9413 5868
rect 9447 5865 9459 5899
rect 9401 5859 9459 5865
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 10873 5899 10931 5905
rect 9732 5868 9904 5896
rect 9732 5856 9738 5868
rect 3510 5828 3516 5840
rect 3471 5800 3516 5828
rect 3510 5788 3516 5800
rect 3568 5788 3574 5840
rect 3694 5788 3700 5840
rect 3752 5828 3758 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 3752 5800 4261 5828
rect 3752 5788 3758 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 4249 5791 4307 5797
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 6318 5831 6376 5837
rect 6318 5828 6330 5831
rect 5408 5800 6330 5828
rect 5408 5788 5414 5800
rect 6318 5797 6330 5800
rect 6364 5797 6376 5831
rect 6318 5791 6376 5797
rect 6546 5788 6552 5840
rect 6604 5828 6610 5840
rect 7668 5828 7696 5856
rect 8202 5828 8208 5840
rect 6604 5800 7696 5828
rect 8163 5800 8208 5828
rect 6604 5788 6610 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 9876 5837 9904 5868
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11054 5896 11060 5908
rect 10919 5868 11060 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11422 5856 11428 5908
rect 11480 5896 11486 5908
rect 11517 5899 11575 5905
rect 11517 5896 11529 5899
rect 11480 5868 11529 5896
rect 11480 5856 11486 5868
rect 11517 5865 11529 5868
rect 11563 5896 11575 5899
rect 12342 5896 12348 5908
rect 11563 5868 12348 5896
rect 11563 5865 11575 5868
rect 11517 5859 11575 5865
rect 12342 5856 12348 5868
rect 12400 5896 12406 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12400 5868 12817 5896
rect 12400 5856 12406 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 13538 5896 13544 5908
rect 13499 5868 13544 5896
rect 12805 5859 12863 5865
rect 13538 5856 13544 5868
rect 13596 5896 13602 5908
rect 13998 5896 14004 5908
rect 13596 5868 14004 5896
rect 13596 5856 13602 5868
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14608 5868 14657 5896
rect 14608 5856 14614 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 15838 5856 15844 5908
rect 15896 5856 15902 5908
rect 16390 5856 16396 5908
rect 16448 5896 16454 5908
rect 17129 5899 17187 5905
rect 17129 5896 17141 5899
rect 16448 5868 17141 5896
rect 16448 5856 16454 5868
rect 17129 5865 17141 5868
rect 17175 5865 17187 5899
rect 17586 5896 17592 5908
rect 17547 5868 17592 5896
rect 17129 5859 17187 5865
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 19426 5896 19432 5908
rect 19387 5868 19432 5896
rect 19426 5856 19432 5868
rect 19484 5896 19490 5908
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 19484 5868 19809 5896
rect 19484 5856 19490 5868
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 19797 5859 19855 5865
rect 23109 5899 23167 5905
rect 23109 5865 23121 5899
rect 23155 5896 23167 5899
rect 24118 5896 24124 5908
rect 23155 5868 24124 5896
rect 23155 5865 23167 5868
rect 23109 5859 23167 5865
rect 24118 5856 24124 5868
rect 24176 5896 24182 5908
rect 24176 5868 24440 5896
rect 24176 5856 24182 5868
rect 9861 5831 9919 5837
rect 9861 5797 9873 5831
rect 9907 5828 9919 5831
rect 10226 5828 10232 5840
rect 9907 5800 10232 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 15856 5828 15884 5856
rect 15580 5800 17724 5828
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 3292 5732 3801 5760
rect 3292 5720 3298 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 5994 5760 6000 5772
rect 5907 5732 6000 5760
rect 3789 5723 3847 5729
rect 2372 5664 2912 5692
rect 3804 5692 3832 5723
rect 5994 5720 6000 5732
rect 6052 5760 6058 5772
rect 6914 5760 6920 5772
rect 6052 5732 6920 5760
rect 6052 5720 6058 5732
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 11974 5760 11980 5772
rect 11931 5732 11980 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 13814 5760 13820 5772
rect 13775 5732 13820 5760
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 15286 5720 15292 5772
rect 15344 5760 15350 5772
rect 15580 5769 15608 5800
rect 17696 5772 17724 5800
rect 17862 5788 17868 5840
rect 17920 5828 17926 5840
rect 19153 5831 19211 5837
rect 17920 5800 18644 5828
rect 17920 5788 17926 5800
rect 18616 5772 18644 5800
rect 19153 5797 19165 5831
rect 19199 5828 19211 5831
rect 20346 5828 20352 5840
rect 19199 5800 20352 5828
rect 19199 5797 19211 5800
rect 19153 5791 19211 5797
rect 20346 5788 20352 5800
rect 20404 5788 20410 5840
rect 22370 5788 22376 5840
rect 22428 5828 22434 5840
rect 24412 5837 24440 5868
rect 22510 5831 22568 5837
rect 22510 5828 22522 5831
rect 22428 5800 22522 5828
rect 22428 5788 22434 5800
rect 22510 5797 22522 5800
rect 22556 5797 22568 5831
rect 22510 5791 22568 5797
rect 24397 5831 24455 5837
rect 24397 5797 24409 5831
rect 24443 5797 24455 5831
rect 24946 5828 24952 5840
rect 24907 5800 24952 5828
rect 24397 5791 24455 5797
rect 24946 5788 24952 5800
rect 25004 5788 25010 5840
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 15344 5732 15577 5760
rect 15344 5720 15350 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 15712 5732 15853 5760
rect 15712 5720 15718 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 16390 5760 16396 5772
rect 16351 5732 16396 5760
rect 15841 5723 15899 5729
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3804 5664 4169 5692
rect 2372 5652 2378 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4798 5692 4804 5704
rect 4759 5664 4804 5692
rect 4157 5655 4215 5661
rect 4798 5652 4804 5664
rect 4856 5692 4862 5704
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 4856 5664 5181 5692
rect 4856 5652 4862 5664
rect 5169 5661 5181 5664
rect 5215 5692 5227 5695
rect 5258 5692 5264 5704
rect 5215 5664 5264 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8110 5692 8116 5704
rect 7975 5664 8116 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9548 5664 9781 5692
rect 9548 5652 9554 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 9769 5655 9827 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 14550 5692 14556 5704
rect 14415 5664 14556 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 14550 5652 14556 5664
rect 14608 5692 14614 5704
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 14608 5664 15025 5692
rect 14608 5652 14614 5664
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15856 5692 15884 5723
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 16574 5720 16580 5772
rect 16632 5760 16638 5772
rect 16761 5763 16819 5769
rect 16761 5760 16773 5763
rect 16632 5732 16773 5760
rect 16632 5720 16638 5732
rect 16761 5729 16773 5732
rect 16807 5760 16819 5763
rect 17586 5760 17592 5772
rect 16807 5732 17592 5760
rect 16807 5729 16819 5732
rect 16761 5723 16819 5729
rect 17586 5720 17592 5732
rect 17644 5720 17650 5772
rect 17678 5720 17684 5772
rect 17736 5760 17742 5772
rect 17736 5732 17781 5760
rect 17736 5720 17742 5732
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18141 5763 18199 5769
rect 18141 5760 18153 5763
rect 18012 5732 18153 5760
rect 18012 5720 18018 5732
rect 18141 5729 18153 5732
rect 18187 5729 18199 5763
rect 18598 5760 18604 5772
rect 18559 5732 18604 5760
rect 18141 5723 18199 5729
rect 16666 5692 16672 5704
rect 15856 5664 16672 5692
rect 15013 5655 15071 5661
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 16850 5692 16856 5704
rect 16811 5664 16856 5692
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 18156 5692 18184 5723
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 18966 5760 18972 5772
rect 18927 5732 18972 5760
rect 18966 5720 18972 5732
rect 19024 5720 19030 5772
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20496 5732 20913 5760
rect 20496 5720 20502 5732
rect 20901 5729 20913 5732
rect 20947 5760 20959 5763
rect 21821 5763 21879 5769
rect 21821 5760 21833 5763
rect 20947 5732 21833 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 21821 5729 21833 5732
rect 21867 5729 21879 5763
rect 22186 5760 22192 5772
rect 22147 5732 22192 5760
rect 21821 5723 21879 5729
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 18414 5692 18420 5704
rect 18156 5664 18420 5692
rect 18414 5652 18420 5664
rect 18472 5692 18478 5704
rect 19242 5692 19248 5704
rect 18472 5664 19248 5692
rect 18472 5652 18478 5664
rect 19242 5652 19248 5664
rect 19300 5652 19306 5704
rect 24305 5695 24363 5701
rect 24305 5661 24317 5695
rect 24351 5692 24363 5695
rect 25038 5692 25044 5704
rect 24351 5664 25044 5692
rect 24351 5661 24363 5664
rect 24305 5655 24363 5661
rect 25038 5652 25044 5664
rect 25096 5652 25102 5704
rect 8665 5627 8723 5633
rect 8665 5593 8677 5627
rect 8711 5624 8723 5627
rect 12526 5624 12532 5636
rect 8711 5596 9168 5624
rect 12439 5596 12532 5624
rect 8711 5593 8723 5596
rect 8665 5587 8723 5593
rect 9140 5568 9168 5596
rect 12526 5584 12532 5596
rect 12584 5624 12590 5636
rect 13722 5624 13728 5636
rect 12584 5596 13728 5624
rect 12584 5584 12590 5596
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 21450 5624 21456 5636
rect 21411 5596 21456 5624
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 6914 5556 6920 5568
rect 6875 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 9122 5556 9128 5568
rect 9083 5528 9128 5556
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 15746 5516 15752 5568
rect 15804 5556 15810 5568
rect 16114 5556 16120 5568
rect 15804 5528 16120 5556
rect 15804 5516 15810 5528
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 21085 5559 21143 5565
rect 21085 5525 21097 5559
rect 21131 5556 21143 5559
rect 21634 5556 21640 5568
rect 21131 5528 21640 5556
rect 21131 5525 21143 5528
rect 21085 5519 21143 5525
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 24029 5559 24087 5565
rect 24029 5525 24041 5559
rect 24075 5556 24087 5559
rect 24210 5556 24216 5568
rect 24075 5528 24216 5556
rect 24075 5525 24087 5528
rect 24029 5519 24087 5525
rect 24210 5516 24216 5528
rect 24268 5556 24274 5568
rect 24670 5556 24676 5568
rect 24268 5528 24676 5556
rect 24268 5516 24274 5528
rect 24670 5516 24676 5528
rect 24728 5516 24734 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2038 5352 2044 5364
rect 1999 5324 2044 5352
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 3694 5352 3700 5364
rect 3655 5324 3700 5352
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 5994 5352 6000 5364
rect 5767 5324 6000 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8202 5352 8208 5364
rect 7975 5324 8208 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10226 5352 10232 5364
rect 9815 5324 10232 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 13630 5352 13636 5364
rect 13591 5324 13636 5352
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 13740 5324 16252 5352
rect 7282 5244 7288 5296
rect 7340 5284 7346 5296
rect 7469 5287 7527 5293
rect 7469 5284 7481 5287
rect 7340 5256 7481 5284
rect 7340 5244 7346 5256
rect 7469 5253 7481 5256
rect 7515 5253 7527 5287
rect 11882 5284 11888 5296
rect 11843 5256 11888 5284
rect 7469 5247 7527 5253
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 13740 5284 13768 5324
rect 15654 5284 15660 5296
rect 13004 5256 13768 5284
rect 15615 5256 15660 5284
rect 2958 5216 2964 5228
rect 2919 5188 2964 5216
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4522 5216 4528 5228
rect 4479 5188 4528 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4798 5216 4804 5228
rect 4759 5188 4804 5216
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5408 5188 6009 5216
rect 5408 5176 5414 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 7558 5216 7564 5228
rect 6963 5188 7564 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 9122 5216 9128 5228
rect 9035 5188 9128 5216
rect 9122 5176 9128 5188
rect 9180 5216 9186 5228
rect 10042 5216 10048 5228
rect 9180 5188 10048 5216
rect 9180 5176 9186 5188
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 10778 5216 10784 5228
rect 10735 5188 10784 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12492 5188 12537 5216
rect 12492 5176 12498 5188
rect 13004 5160 13032 5256
rect 15654 5244 15660 5256
rect 15712 5284 15718 5296
rect 16114 5284 16120 5296
rect 15712 5256 16120 5284
rect 15712 5244 15718 5256
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 16224 5284 16252 5324
rect 18966 5312 18972 5364
rect 19024 5352 19030 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 19024 5324 19073 5352
rect 19024 5312 19030 5324
rect 19061 5321 19073 5324
rect 19107 5321 19119 5355
rect 19061 5315 19119 5321
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19392 5324 19441 5352
rect 19392 5312 19398 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 22244 5324 22753 5352
rect 22244 5312 22250 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 22741 5315 22799 5321
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 16224 5256 17785 5284
rect 17773 5253 17785 5256
rect 17819 5284 17831 5287
rect 24946 5284 24952 5296
rect 17819 5256 18368 5284
rect 24907 5256 24952 5284
rect 17819 5253 17831 5256
rect 17773 5247 17831 5253
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 14292 5188 16865 5216
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1486 5148 1492 5160
rect 1443 5120 1492 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1486 5108 1492 5120
rect 1544 5108 1550 5160
rect 12250 5148 12256 5160
rect 12163 5120 12256 5148
rect 12250 5108 12256 5120
rect 12308 5148 12314 5160
rect 12986 5148 12992 5160
rect 12308 5120 12992 5148
rect 12308 5108 12314 5120
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14292 5157 14320 5188
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 13872 5120 14289 5148
rect 13872 5108 13878 5120
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 14369 5151 14427 5157
rect 14369 5117 14381 5151
rect 14415 5117 14427 5151
rect 14550 5148 14556 5160
rect 14511 5120 14556 5148
rect 14369 5111 14427 5117
rect 2685 5083 2743 5089
rect 2685 5049 2697 5083
rect 2731 5049 2743 5083
rect 2685 5043 2743 5049
rect 2777 5083 2835 5089
rect 2777 5049 2789 5083
rect 2823 5080 2835 5083
rect 3694 5080 3700 5092
rect 2823 5052 3700 5080
rect 2823 5049 2835 5052
rect 2777 5043 2835 5049
rect 2498 5012 2504 5024
rect 2459 4984 2504 5012
rect 2498 4972 2504 4984
rect 2556 5012 2562 5024
rect 2700 5012 2728 5043
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 4525 5083 4583 5089
rect 4525 5080 4537 5083
rect 4264 5052 4537 5080
rect 4264 5024 4292 5052
rect 4525 5049 4537 5052
rect 4571 5080 4583 5083
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 4571 5052 6561 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 6549 5049 6561 5052
rect 6595 5080 6607 5083
rect 6914 5080 6920 5092
rect 6595 5052 6920 5080
rect 6595 5049 6607 5052
rect 6549 5043 6607 5049
rect 6914 5040 6920 5052
rect 6972 5080 6978 5092
rect 7009 5083 7067 5089
rect 7009 5080 7021 5083
rect 6972 5052 7021 5080
rect 6972 5040 6978 5052
rect 7009 5049 7021 5052
rect 7055 5049 7067 5083
rect 8478 5080 8484 5092
rect 8439 5052 8484 5080
rect 7009 5043 7067 5049
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 8573 5083 8631 5089
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 9398 5080 9404 5092
rect 8619 5052 9404 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 4246 5012 4252 5024
rect 2556 4984 2728 5012
rect 4207 4984 4252 5012
rect 2556 4972 2562 4984
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 8588 5012 8616 5043
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 9858 5040 9864 5092
rect 9916 5080 9922 5092
rect 10137 5083 10195 5089
rect 10137 5080 10149 5083
rect 9916 5052 10149 5080
rect 9916 5040 9922 5052
rect 10137 5049 10149 5052
rect 10183 5049 10195 5083
rect 14090 5080 14096 5092
rect 14051 5052 14096 5080
rect 10137 5043 10195 5049
rect 14090 5040 14096 5052
rect 14148 5080 14154 5092
rect 14384 5080 14412 5111
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 15856 5157 15884 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18141 5219 18199 5225
rect 18141 5216 18153 5219
rect 18012 5188 18153 5216
rect 18012 5176 18018 5188
rect 18141 5185 18153 5188
rect 18187 5185 18199 5219
rect 18141 5179 18199 5185
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5117 15899 5151
rect 15841 5111 15899 5117
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5117 15991 5151
rect 16114 5148 16120 5160
rect 16075 5120 16120 5148
rect 15933 5111 15991 5117
rect 15289 5083 15347 5089
rect 15289 5080 15301 5083
rect 14148 5052 15301 5080
rect 14148 5040 14154 5052
rect 15289 5049 15301 5052
rect 15335 5080 15347 5083
rect 15948 5080 15976 5111
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 18340 5157 18368 5256
rect 24946 5244 24952 5256
rect 25004 5244 25010 5296
rect 18506 5216 18512 5228
rect 18467 5188 18512 5216
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21450 5216 21456 5228
rect 21223 5188 21456 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 21450 5176 21456 5188
rect 21508 5176 21514 5228
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 25317 5219 25375 5225
rect 25317 5216 25329 5219
rect 24176 5188 25329 5216
rect 24176 5176 24182 5188
rect 25317 5185 25329 5188
rect 25363 5185 25375 5219
rect 25317 5179 25375 5185
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5117 18383 5151
rect 18325 5111 18383 5117
rect 20257 5151 20315 5157
rect 20257 5117 20269 5151
rect 20303 5148 20315 5151
rect 20530 5148 20536 5160
rect 20303 5120 20536 5148
rect 20303 5117 20315 5120
rect 20257 5111 20315 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 20714 5148 20720 5160
rect 20675 5120 20720 5148
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 20346 5080 20352 5092
rect 15335 5052 15976 5080
rect 20307 5052 20352 5080
rect 15335 5049 15347 5052
rect 15289 5043 15347 5049
rect 15856 5024 15884 5052
rect 20346 5040 20352 5052
rect 20404 5040 20410 5092
rect 21498 5083 21556 5089
rect 21498 5049 21510 5083
rect 21544 5080 21556 5083
rect 22370 5080 22376 5092
rect 21544 5052 22376 5080
rect 21544 5049 21556 5052
rect 21498 5043 21556 5049
rect 8343 4984 8616 5012
rect 11333 5015 11391 5021
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 11974 5012 11980 5024
rect 11379 4984 11980 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 11974 4972 11980 4984
rect 12032 4972 12038 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14737 5015 14795 5021
rect 14737 5012 14749 5015
rect 14240 4984 14749 5012
rect 14240 4972 14246 4984
rect 14737 4981 14749 4984
rect 14783 4981 14795 5015
rect 14737 4975 14795 4981
rect 15838 4972 15844 5024
rect 15896 4972 15902 5024
rect 16298 5012 16304 5024
rect 16259 4984 16304 5012
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 17497 5015 17555 5021
rect 17497 4981 17509 5015
rect 17543 5012 17555 5015
rect 17678 5012 17684 5024
rect 17543 4984 17684 5012
rect 17543 4981 17555 4984
rect 17497 4975 17555 4981
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20956 4984 21005 5012
rect 20956 4972 20962 4984
rect 20993 4981 21005 4984
rect 21039 5012 21051 5015
rect 21513 5012 21541 5043
rect 22370 5040 22376 5052
rect 22428 5040 22434 5092
rect 23477 5083 23535 5089
rect 23477 5049 23489 5083
rect 23523 5080 23535 5083
rect 23842 5080 23848 5092
rect 23523 5052 23848 5080
rect 23523 5049 23535 5052
rect 23477 5043 23535 5049
rect 23842 5040 23848 5052
rect 23900 5080 23906 5092
rect 24397 5083 24455 5089
rect 24397 5080 24409 5083
rect 23900 5052 24409 5080
rect 23900 5040 23906 5052
rect 24397 5049 24409 5052
rect 24443 5049 24455 5083
rect 24397 5043 24455 5049
rect 24489 5083 24547 5089
rect 24489 5049 24501 5083
rect 24535 5049 24547 5083
rect 24489 5043 24547 5049
rect 21039 4984 21541 5012
rect 22097 5015 22155 5021
rect 21039 4981 21051 4984
rect 20993 4975 21051 4981
rect 22097 4981 22109 5015
rect 22143 5012 22155 5015
rect 22646 5012 22652 5024
rect 22143 4984 22652 5012
rect 22143 4981 22155 4984
rect 22097 4975 22155 4981
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 24210 5012 24216 5024
rect 24171 4984 24216 5012
rect 24210 4972 24216 4984
rect 24268 5012 24274 5024
rect 24504 5012 24532 5043
rect 24268 4984 24532 5012
rect 24268 4972 24274 4984
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1452 4780 1593 4808
rect 1452 4768 1458 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1581 4771 1639 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 3200 4780 3249 4808
rect 3200 4768 3206 4780
rect 3237 4777 3249 4780
rect 3283 4808 3295 4811
rect 3694 4808 3700 4820
rect 3283 4780 3700 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 3694 4768 3700 4780
rect 3752 4808 3758 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3752 4780 3801 4808
rect 3752 4768 3758 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 4580 4780 5089 4808
rect 4580 4768 4586 4780
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 5077 4771 5135 4777
rect 6227 4811 6285 4817
rect 6227 4777 6239 4811
rect 6273 4808 6285 4811
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 6273 4780 8401 4808
rect 6273 4777 6285 4780
rect 6227 4771 6285 4777
rect 8389 4777 8401 4780
rect 8435 4808 8447 4811
rect 8478 4808 8484 4820
rect 8435 4780 8484 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9916 4780 9965 4808
rect 9916 4768 9922 4780
rect 9953 4777 9965 4780
rect 9999 4777 10011 4811
rect 9953 4771 10011 4777
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 10192 4780 10425 4808
rect 10192 4768 10198 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 10413 4771 10471 4777
rect 1762 4700 1768 4752
rect 1820 4740 1826 4752
rect 2222 4740 2228 4752
rect 1820 4712 2228 4740
rect 1820 4700 1826 4712
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 2682 4740 2688 4752
rect 2363 4712 2688 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 2682 4700 2688 4712
rect 2740 4700 2746 4752
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 2958 4740 2964 4752
rect 2915 4712 2964 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 4154 4700 4160 4752
rect 4212 4740 4218 4752
rect 4249 4743 4307 4749
rect 4249 4740 4261 4743
rect 4212 4712 4261 4740
rect 4212 4700 4218 4712
rect 4249 4709 4261 4712
rect 4295 4709 4307 4743
rect 4798 4740 4804 4752
rect 4759 4712 4804 4740
rect 4249 4703 4307 4709
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 7009 4743 7067 4749
rect 7009 4709 7021 4743
rect 7055 4740 7067 4743
rect 7190 4740 7196 4752
rect 7055 4712 7196 4740
rect 7055 4709 7067 4712
rect 7009 4703 7067 4709
rect 7190 4700 7196 4712
rect 7248 4700 7254 4752
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 10428 4740 10456 4771
rect 12526 4768 12532 4820
rect 12584 4808 12590 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 12584 4780 13277 4808
rect 12584 4768 12590 4780
rect 13265 4777 13277 4780
rect 13311 4808 13323 4811
rect 15381 4811 15439 4817
rect 15381 4808 15393 4811
rect 13311 4780 15393 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 15381 4777 15393 4780
rect 15427 4777 15439 4811
rect 15381 4771 15439 4777
rect 16666 4768 16672 4820
rect 16724 4808 16730 4820
rect 17037 4811 17095 4817
rect 17037 4808 17049 4811
rect 16724 4780 17049 4808
rect 16724 4768 16730 4780
rect 17037 4777 17049 4780
rect 17083 4777 17095 4811
rect 17037 4771 17095 4777
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 17497 4811 17555 4817
rect 17497 4808 17509 4811
rect 17276 4780 17509 4808
rect 17276 4768 17282 4780
rect 17497 4777 17509 4780
rect 17543 4808 17555 4811
rect 18874 4808 18880 4820
rect 17543 4780 18880 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 20257 4811 20315 4817
rect 20257 4808 20269 4811
rect 19484 4780 20269 4808
rect 19484 4768 19490 4780
rect 20257 4777 20269 4780
rect 20303 4777 20315 4811
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20257 4771 20315 4777
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 23477 4811 23535 4817
rect 23477 4808 23489 4811
rect 23256 4780 23489 4808
rect 23256 4768 23262 4780
rect 23477 4777 23489 4780
rect 23523 4777 23535 4811
rect 23477 4771 23535 4777
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 24305 4811 24363 4817
rect 24305 4808 24317 4811
rect 24268 4780 24317 4808
rect 24268 4768 24274 4780
rect 24305 4777 24317 4780
rect 24351 4777 24363 4811
rect 25038 4808 25044 4820
rect 24999 4780 25044 4808
rect 24305 4771 24363 4777
rect 25038 4768 25044 4780
rect 25096 4768 25102 4820
rect 10689 4743 10747 4749
rect 10689 4740 10701 4743
rect 7340 4712 7385 4740
rect 10428 4712 10701 4740
rect 7340 4700 7346 4712
rect 10689 4709 10701 4712
rect 10735 4709 10747 4743
rect 10689 4703 10747 4709
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 15105 4743 15163 4749
rect 10836 4712 10881 4740
rect 10836 4700 10842 4712
rect 15105 4709 15117 4743
rect 15151 4740 15163 4743
rect 15286 4740 15292 4752
rect 15151 4712 15292 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 15286 4700 15292 4712
rect 15344 4700 15350 4752
rect 17954 4700 17960 4752
rect 18012 4740 18018 4752
rect 19014 4743 19072 4749
rect 19014 4740 19026 4743
rect 18012 4712 19026 4740
rect 18012 4700 18018 4712
rect 19014 4709 19026 4712
rect 19060 4709 19072 4743
rect 19014 4703 19072 4709
rect 20346 4700 20352 4752
rect 20404 4740 20410 4752
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 20404 4712 21097 4740
rect 20404 4700 20410 4712
rect 21085 4709 21097 4712
rect 21131 4740 21143 4743
rect 21358 4740 21364 4752
rect 21131 4712 21364 4740
rect 21131 4709 21143 4712
rect 21085 4703 21143 4709
rect 21358 4700 21364 4712
rect 21416 4700 21422 4752
rect 22646 4740 22652 4752
rect 22607 4712 22652 4740
rect 22646 4700 22652 4712
rect 22704 4700 22710 4752
rect 6086 4632 6092 4684
rect 6144 4681 6150 4684
rect 6144 4675 6182 4681
rect 6170 4641 6182 4675
rect 12802 4672 12808 4684
rect 12763 4644 12808 4672
rect 6144 4635 6182 4641
rect 6144 4632 6150 4635
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 14056 4644 14105 4672
rect 14056 4632 14062 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4672 15623 4675
rect 15746 4672 15752 4684
rect 15611 4644 15752 4672
rect 15611 4641 15623 4644
rect 15565 4635 15623 4641
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 15930 4672 15936 4684
rect 15891 4644 15936 4672
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16301 4675 16359 4681
rect 16301 4641 16313 4675
rect 16347 4672 16359 4675
rect 16390 4672 16396 4684
rect 16347 4644 16396 4672
rect 16347 4641 16359 4644
rect 16301 4635 16359 4641
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 16574 4672 16580 4684
rect 16535 4644 16580 4672
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 17586 4672 17592 4684
rect 17547 4644 17592 4672
rect 17586 4632 17592 4644
rect 17644 4632 17650 4684
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 18104 4644 18153 4672
rect 18104 4632 18110 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 24118 4672 24124 4684
rect 24079 4644 24124 4672
rect 18141 4635 18199 4641
rect 24118 4632 24124 4644
rect 24176 4632 24182 4684
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4430 4604 4436 4616
rect 4203 4576 4436 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 6972 4576 7481 4604
rect 6972 4564 6978 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4604 11391 4607
rect 11606 4604 11612 4616
rect 11379 4576 11612 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 13872 4576 14657 4604
rect 13872 4564 13878 4576
rect 14645 4573 14657 4576
rect 14691 4573 14703 4607
rect 18690 4604 18696 4616
rect 18651 4576 18696 4604
rect 14645 4567 14703 4573
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 20990 4604 20996 4616
rect 20951 4576 20996 4604
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 21082 4564 21088 4616
rect 21140 4604 21146 4616
rect 21269 4607 21327 4613
rect 21269 4604 21281 4607
rect 21140 4576 21281 4604
rect 21140 4564 21146 4576
rect 21269 4573 21281 4576
rect 21315 4573 21327 4607
rect 22278 4604 22284 4616
rect 22239 4576 22284 4604
rect 21269 4567 21327 4573
rect 22278 4564 22284 4576
rect 22336 4564 22342 4616
rect 22557 4607 22615 4613
rect 22557 4573 22569 4607
rect 22603 4604 22615 4607
rect 23198 4604 23204 4616
rect 22603 4576 23204 4604
rect 22603 4573 22615 4576
rect 22557 4567 22615 4573
rect 23198 4564 23204 4576
rect 23256 4564 23262 4616
rect 4246 4496 4252 4548
rect 4304 4536 4310 4548
rect 5074 4536 5080 4548
rect 4304 4508 5080 4536
rect 4304 4496 4310 4508
rect 5074 4496 5080 4508
rect 5132 4496 5138 4548
rect 8754 4496 8760 4548
rect 8812 4536 8818 4548
rect 9401 4539 9459 4545
rect 9401 4536 9413 4539
rect 8812 4508 9413 4536
rect 8812 4496 8818 4508
rect 9401 4505 9413 4508
rect 9447 4536 9459 4539
rect 9490 4536 9496 4548
rect 9447 4508 9496 4536
rect 9447 4505 9459 4508
rect 9401 4499 9459 4505
rect 9490 4496 9496 4508
rect 9548 4496 9554 4548
rect 14274 4536 14280 4548
rect 14235 4508 14280 4536
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 19613 4539 19671 4545
rect 19613 4505 19625 4539
rect 19659 4536 19671 4539
rect 19981 4539 20039 4545
rect 19981 4536 19993 4539
rect 19659 4508 19993 4536
rect 19659 4505 19671 4508
rect 19613 4499 19671 4505
rect 19981 4505 19993 4508
rect 20027 4536 20039 4539
rect 20530 4536 20536 4548
rect 20027 4508 20536 4536
rect 20027 4505 20039 4508
rect 19981 4499 20039 4505
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 21008 4536 21036 4564
rect 21913 4539 21971 4545
rect 21913 4536 21925 4539
rect 21008 4508 21925 4536
rect 21913 4505 21925 4508
rect 21959 4505 21971 4539
rect 21913 4499 21971 4505
rect 22370 4496 22376 4548
rect 22428 4536 22434 4548
rect 23109 4539 23167 4545
rect 23109 4536 23121 4539
rect 22428 4508 23121 4536
rect 22428 4496 22434 4508
rect 23109 4505 23121 4508
rect 23155 4505 23167 4539
rect 23109 4499 23167 4505
rect 9122 4468 9128 4480
rect 9083 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 11977 4471 12035 4477
rect 11977 4468 11989 4471
rect 11756 4440 11989 4468
rect 11756 4428 11762 4440
rect 11977 4437 11989 4440
rect 12023 4437 12035 4471
rect 12618 4468 12624 4480
rect 12579 4440 12624 4468
rect 11977 4431 12035 4437
rect 12618 4428 12624 4440
rect 12676 4428 12682 4480
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 13722 4468 13728 4480
rect 13679 4440 13728 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 13998 4468 14004 4480
rect 13959 4440 14004 4468
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 17770 4468 17776 4480
rect 17731 4440 17776 4468
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 18506 4468 18512 4480
rect 18467 4440 18512 4468
rect 18506 4428 18512 4440
rect 18564 4428 18570 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 4154 4264 4160 4276
rect 4115 4236 4160 4264
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 4430 4264 4436 4276
rect 4391 4236 4436 4264
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 6086 4224 6092 4276
rect 6144 4264 6150 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 6144 4236 6193 4264
rect 6144 4224 6150 4236
rect 6181 4233 6193 4236
rect 6227 4233 6239 4267
rect 6181 4227 6239 4233
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 12860 4236 13461 4264
rect 12860 4224 12866 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 13449 4227 13507 4233
rect 13909 4267 13967 4273
rect 13909 4233 13921 4267
rect 13955 4264 13967 4267
rect 13998 4264 14004 4276
rect 13955 4236 14004 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 17865 4267 17923 4273
rect 17865 4233 17877 4267
rect 17911 4264 17923 4267
rect 17954 4264 17960 4276
rect 17911 4236 17960 4264
rect 17911 4233 17923 4236
rect 17865 4227 17923 4233
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 21358 4264 21364 4276
rect 21319 4236 21364 4264
rect 21358 4224 21364 4236
rect 21416 4224 21422 4276
rect 22646 4224 22652 4276
rect 22704 4264 22710 4276
rect 23017 4267 23075 4273
rect 23017 4264 23029 4267
rect 22704 4236 23029 4264
rect 22704 4224 22710 4236
rect 23017 4233 23029 4236
rect 23063 4264 23075 4267
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 23063 4236 23397 4264
rect 23063 4233 23075 4236
rect 23017 4227 23075 4233
rect 23385 4233 23397 4236
rect 23431 4233 23443 4267
rect 23385 4227 23443 4233
rect 4338 4156 4344 4208
rect 4396 4156 4402 4208
rect 16853 4199 16911 4205
rect 16853 4196 16865 4199
rect 15948 4168 16865 4196
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3053 4131 3111 4137
rect 2832 4100 2877 4128
rect 2832 4088 2838 4100
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3418 4128 3424 4140
rect 3099 4100 3424 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 4356 4128 4384 4156
rect 15948 4140 15976 4168
rect 16853 4165 16865 4168
rect 16899 4196 16911 4199
rect 17402 4196 17408 4208
rect 16899 4168 17408 4196
rect 16899 4165 16911 4168
rect 16853 4159 16911 4165
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 6546 4128 6552 4140
rect 3743 4100 4384 4128
rect 6507 4100 6552 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 7558 4128 7564 4140
rect 7519 4100 7564 4128
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7834 4128 7840 4140
rect 7795 4100 7840 4128
rect 7834 4088 7840 4100
rect 7892 4128 7898 4140
rect 9122 4128 9128 4140
rect 7892 4100 9128 4128
rect 7892 4088 7898 4100
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9490 4088 9496 4140
rect 9548 4128 9554 4140
rect 9766 4128 9772 4140
rect 9548 4100 9772 4128
rect 9548 4088 9554 4100
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4128 14335 4131
rect 15930 4128 15936 4140
rect 14323 4100 15936 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 1394 4060 1400 4072
rect 1355 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4020 1458 4072
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 2406 4060 2412 4072
rect 1903 4032 2412 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 5123 4032 5825 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5813 4029 5825 4032
rect 5859 4060 5871 4063
rect 6178 4060 6184 4072
rect 5859 4032 6184 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10594 4060 10600 4072
rect 10183 4032 10600 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 11885 4063 11943 4069
rect 11885 4029 11897 4063
rect 11931 4060 11943 4063
rect 12066 4060 12072 4072
rect 11931 4032 12072 4060
rect 11931 4029 11943 4032
rect 11885 4023 11943 4029
rect 12066 4020 12072 4032
rect 12124 4060 12130 4072
rect 12802 4060 12808 4072
rect 12124 4032 12808 4060
rect 12124 4020 12130 4032
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4060 14703 4063
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 14691 4032 15025 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 15013 4029 15025 4032
rect 15059 4060 15071 4063
rect 15102 4060 15108 4072
rect 15059 4032 15108 4060
rect 15059 4029 15071 4032
rect 15013 4023 15071 4029
rect 15102 4020 15108 4032
rect 15160 4060 15166 4072
rect 15381 4063 15439 4069
rect 15381 4060 15393 4063
rect 15160 4032 15393 4060
rect 15160 4020 15166 4032
rect 15381 4029 15393 4032
rect 15427 4060 15439 4063
rect 15746 4060 15752 4072
rect 15427 4032 15752 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 15856 4069 15884 4100
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16390 4128 16396 4140
rect 16132 4100 16396 4128
rect 16132 4069 16160 4100
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 18138 4128 18144 4140
rect 17543 4100 18144 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 18138 4088 18144 4100
rect 18196 4128 18202 4140
rect 18196 4100 18920 4128
rect 18196 4088 18202 4100
rect 18892 4072 18920 4100
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 20441 4131 20499 4137
rect 19024 4100 19380 4128
rect 19024 4088 19030 4100
rect 15841 4063 15899 4069
rect 15841 4029 15853 4063
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 16485 4063 16543 4069
rect 16485 4029 16497 4063
rect 16531 4060 16543 4063
rect 16666 4060 16672 4072
rect 16531 4032 16672 4060
rect 16531 4029 16543 4032
rect 16485 4023 16543 4029
rect 16666 4020 16672 4032
rect 16724 4060 16730 4072
rect 17218 4060 17224 4072
rect 16724 4032 17224 4060
rect 16724 4020 16730 4032
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18472 4032 18521 4060
rect 18472 4020 18478 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18874 4060 18880 4072
rect 18835 4032 18880 4060
rect 18509 4023 18567 4029
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 19352 4069 19380 4100
rect 20441 4097 20453 4131
rect 20487 4128 20499 4131
rect 20622 4128 20628 4140
rect 20487 4100 20628 4128
rect 20487 4097 20499 4100
rect 20441 4091 20499 4097
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 21082 4128 21088 4140
rect 21043 4100 21088 4128
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22370 4128 22376 4140
rect 22152 4100 22197 4128
rect 22331 4100 22376 4128
rect 22152 4088 22158 4100
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 19337 4063 19395 4069
rect 19337 4029 19349 4063
rect 19383 4029 19395 4063
rect 23400 4060 23428 4227
rect 24118 4224 24124 4276
rect 24176 4264 24182 4276
rect 24673 4267 24731 4273
rect 24673 4264 24685 4267
rect 24176 4236 24685 4264
rect 24176 4224 24182 4236
rect 24673 4233 24685 4236
rect 24719 4233 24731 4267
rect 24673 4227 24731 4233
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 25556 4100 25789 4128
rect 25556 4088 25562 4100
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 25777 4091 25835 4097
rect 23753 4063 23811 4069
rect 23753 4060 23765 4063
rect 23400 4032 23765 4060
rect 19337 4023 19395 4029
rect 23753 4029 23765 4032
rect 23799 4029 23811 4063
rect 23753 4023 23811 4029
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 25516 4060 25544 4088
rect 25271 4032 25544 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 3200 3964 3245 3992
rect 3200 3952 3206 3964
rect 5994 3952 6000 4004
rect 6052 3992 6058 4004
rect 7285 3995 7343 4001
rect 7285 3992 7297 3995
rect 6052 3964 7297 3992
rect 6052 3952 6058 3964
rect 7285 3961 7297 3964
rect 7331 3961 7343 3995
rect 7285 3955 7343 3961
rect 7653 3995 7711 4001
rect 7653 3961 7665 3995
rect 7699 3961 7711 3995
rect 7653 3955 7711 3961
rect 5442 3924 5448 3936
rect 5403 3896 5448 3924
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 7300 3924 7328 3955
rect 7668 3924 7696 3955
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 8481 3995 8539 4001
rect 8481 3992 8493 3995
rect 7800 3964 8493 3992
rect 7800 3952 7806 3964
rect 8481 3961 8493 3964
rect 8527 3961 8539 3995
rect 8481 3955 8539 3961
rect 8941 3995 8999 4001
rect 8941 3961 8953 3995
rect 8987 3992 8999 3995
rect 9214 3992 9220 4004
rect 8987 3964 9220 3992
rect 8987 3961 8999 3964
rect 8941 3955 8999 3961
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 10505 3995 10563 4001
rect 10505 3992 10517 3995
rect 9640 3964 10517 3992
rect 9640 3952 9646 3964
rect 10505 3961 10517 3964
rect 10551 3992 10563 3995
rect 10959 3995 11017 4001
rect 10959 3992 10971 3995
rect 10551 3964 10971 3992
rect 10551 3961 10563 3964
rect 10505 3955 10563 3961
rect 10959 3961 10971 3964
rect 11005 3992 11017 3995
rect 12253 3995 12311 4001
rect 12253 3992 12265 3995
rect 11005 3964 12265 3992
rect 11005 3961 11017 3964
rect 10959 3955 11017 3961
rect 12253 3961 12265 3964
rect 12299 3992 12311 3995
rect 12891 3995 12949 4001
rect 12891 3992 12903 3995
rect 12299 3964 12903 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12891 3961 12903 3964
rect 12937 3992 12949 3995
rect 17862 3992 17868 4004
rect 12937 3964 17868 3992
rect 12937 3961 12949 3964
rect 12891 3955 12949 3961
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 18690 3952 18696 4004
rect 18748 3992 18754 4004
rect 19518 3992 19524 4004
rect 18748 3964 19524 3992
rect 18748 3952 18754 3964
rect 19518 3952 19524 3964
rect 19576 3952 19582 4004
rect 20530 3952 20536 4004
rect 20588 3992 20594 4004
rect 22189 3995 22247 4001
rect 20588 3964 20633 3992
rect 20588 3952 20594 3964
rect 22189 3961 22201 3995
rect 22235 3961 22247 3995
rect 23661 3995 23719 4001
rect 23661 3992 23673 3995
rect 22189 3955 22247 3961
rect 22848 3964 23673 3992
rect 11514 3924 11520 3936
rect 7300 3896 7696 3924
rect 11475 3896 11520 3924
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 15194 3924 15200 3936
rect 15155 3896 15200 3924
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 19889 3927 19947 3933
rect 19889 3893 19901 3927
rect 19935 3924 19947 3927
rect 19978 3924 19984 3936
rect 19935 3896 19984 3924
rect 19935 3893 19947 3896
rect 19889 3887 19947 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20162 3924 20168 3936
rect 20123 3896 20168 3924
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 21913 3927 21971 3933
rect 21913 3893 21925 3927
rect 21959 3924 21971 3927
rect 22204 3924 22232 3955
rect 22848 3924 22876 3964
rect 23661 3961 23673 3964
rect 23707 3961 23719 3995
rect 23661 3955 23719 3961
rect 25406 3924 25412 3936
rect 21959 3896 22876 3924
rect 25367 3896 25412 3924
rect 21959 3893 21971 3896
rect 21913 3887 21971 3893
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 2222 3720 2228 3732
rect 2183 3692 2228 3720
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2682 3720 2688 3732
rect 2643 3692 2688 3720
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 3108 3692 3157 3720
rect 3108 3680 3114 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3145 3683 3203 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 6086 3720 6092 3732
rect 5316 3692 6092 3720
rect 5316 3680 5322 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9815 3723 9873 3729
rect 9815 3720 9827 3723
rect 9732 3692 9827 3720
rect 9732 3680 9738 3692
rect 9815 3689 9827 3692
rect 9861 3689 9873 3723
rect 9815 3683 9873 3689
rect 10321 3723 10379 3729
rect 10321 3689 10333 3723
rect 10367 3720 10379 3723
rect 10686 3720 10692 3732
rect 10367 3692 10692 3720
rect 10367 3689 10379 3692
rect 10321 3683 10379 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 12066 3720 12072 3732
rect 12027 3692 12072 3720
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 15102 3720 15108 3732
rect 15063 3692 15108 3720
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 15378 3720 15384 3732
rect 15339 3692 15384 3720
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 16632 3692 17141 3720
rect 16632 3680 16638 3692
rect 17129 3689 17141 3692
rect 17175 3720 17187 3723
rect 17497 3723 17555 3729
rect 17497 3720 17509 3723
rect 17175 3692 17509 3720
rect 17175 3689 17187 3692
rect 17129 3683 17187 3689
rect 17497 3689 17509 3692
rect 17543 3720 17555 3723
rect 17543 3692 18920 3720
rect 17543 3689 17555 3692
rect 17497 3683 17555 3689
rect 5442 3652 5448 3664
rect 4264 3624 5448 3652
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 2130 3584 2136 3596
rect 1443 3556 2136 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 2130 3544 2136 3556
rect 2188 3544 2194 3596
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3142 3584 3148 3596
rect 3007 3556 3148 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3142 3544 3148 3556
rect 3200 3584 3206 3596
rect 3970 3584 3976 3596
rect 3200 3556 3976 3584
rect 3200 3544 3206 3556
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4264 3593 4292 3624
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 5994 3652 6000 3664
rect 5955 3624 6000 3652
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 6549 3655 6607 3661
rect 6549 3621 6561 3655
rect 6595 3652 6607 3655
rect 6914 3652 6920 3664
rect 6595 3624 6920 3652
rect 6595 3621 6607 3624
rect 6549 3615 6607 3621
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7739 3655 7797 3661
rect 7739 3621 7751 3655
rect 7785 3652 7797 3655
rect 8110 3652 8116 3664
rect 7785 3624 8116 3652
rect 7785 3621 7797 3624
rect 7739 3615 7797 3621
rect 8110 3612 8116 3624
rect 8168 3652 8174 3664
rect 8662 3652 8668 3664
rect 8168 3624 8668 3652
rect 8168 3612 8174 3624
rect 8662 3612 8668 3624
rect 8720 3652 8726 3664
rect 9582 3652 9588 3664
rect 8720 3624 9588 3652
rect 8720 3612 8726 3624
rect 9582 3612 9588 3624
rect 9640 3612 9646 3664
rect 11146 3652 11152 3664
rect 11107 3624 11152 3652
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 11698 3652 11704 3664
rect 11659 3624 11704 3652
rect 11698 3612 11704 3624
rect 11756 3612 11762 3664
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 12713 3655 12771 3661
rect 12713 3652 12725 3655
rect 12676 3624 12725 3652
rect 12676 3612 12682 3624
rect 12713 3621 12725 3624
rect 12759 3621 12771 3655
rect 12713 3615 12771 3621
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14737 3655 14795 3661
rect 14737 3652 14749 3655
rect 14056 3624 14749 3652
rect 14056 3612 14062 3624
rect 14737 3621 14749 3624
rect 14783 3652 14795 3655
rect 16390 3652 16396 3664
rect 14783 3624 16396 3652
rect 14783 3621 14795 3624
rect 14737 3615 14795 3621
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 18414 3652 18420 3664
rect 18340 3624 18420 3652
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4614 3584 4620 3596
rect 4571 3556 4620 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4982 3584 4988 3596
rect 4943 3556 4988 3584
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7374 3584 7380 3596
rect 6880 3556 7380 3584
rect 6880 3544 6886 3556
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9712 3587 9770 3593
rect 9712 3584 9724 3587
rect 8996 3556 9724 3584
rect 8996 3544 9002 3556
rect 9712 3553 9724 3556
rect 9758 3584 9770 3587
rect 10042 3584 10048 3596
rect 9758 3556 10048 3584
rect 9758 3553 9770 3556
rect 9712 3547 9770 3553
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 14093 3587 14151 3593
rect 14093 3553 14105 3587
rect 14139 3584 14151 3587
rect 14366 3584 14372 3596
rect 14139 3556 14372 3584
rect 14139 3553 14151 3556
rect 14093 3547 14151 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15160 3556 15301 3584
rect 15160 3544 15166 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15930 3584 15936 3596
rect 15891 3556 15936 3584
rect 15289 3547 15347 3553
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16206 3584 16212 3596
rect 16167 3556 16212 3584
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16666 3584 16672 3596
rect 16627 3556 16672 3584
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 17678 3584 17684 3596
rect 17639 3556 17684 3584
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 18340 3593 18368 3624
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 18325 3587 18383 3593
rect 18325 3553 18337 3587
rect 18371 3553 18383 3587
rect 18506 3584 18512 3596
rect 18419 3556 18512 3584
rect 18325 3547 18383 3553
rect 18506 3544 18512 3556
rect 18564 3544 18570 3596
rect 18892 3593 18920 3692
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19576 3692 19809 3720
rect 19576 3680 19582 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 19797 3683 19855 3689
rect 20441 3723 20499 3729
rect 20441 3689 20453 3723
rect 20487 3720 20499 3723
rect 20530 3720 20536 3732
rect 20487 3692 20536 3720
rect 20487 3689 20499 3692
rect 20441 3683 20499 3689
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 23477 3723 23535 3729
rect 23477 3720 23489 3723
rect 22152 3692 22197 3720
rect 22572 3692 23489 3720
rect 22152 3680 22158 3692
rect 21082 3652 21088 3664
rect 21043 3624 21088 3652
rect 21082 3612 21088 3624
rect 21140 3612 21146 3664
rect 21910 3612 21916 3664
rect 21968 3652 21974 3664
rect 22572 3661 22600 3692
rect 23477 3689 23489 3692
rect 23523 3689 23535 3723
rect 23477 3683 23535 3689
rect 22557 3655 22615 3661
rect 22557 3652 22569 3655
rect 21968 3624 22569 3652
rect 21968 3612 21974 3624
rect 22557 3621 22569 3624
rect 22603 3621 22615 3655
rect 22557 3615 22615 3621
rect 22649 3655 22707 3661
rect 22649 3621 22661 3655
rect 22695 3652 22707 3655
rect 22738 3652 22744 3664
rect 22695 3624 22744 3652
rect 22695 3621 22707 3624
rect 22649 3615 22707 3621
rect 22738 3612 22744 3624
rect 22796 3612 22802 3664
rect 24026 3652 24032 3664
rect 23987 3624 24032 3652
rect 24026 3612 24032 3624
rect 24084 3612 24090 3664
rect 18877 3587 18935 3593
rect 18877 3553 18889 3587
rect 18923 3584 18935 3587
rect 19242 3584 19248 3596
rect 18923 3556 19248 3584
rect 18923 3553 18935 3556
rect 18877 3547 18935 3553
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 24670 3584 24676 3596
rect 24631 3556 24676 3584
rect 24670 3544 24676 3556
rect 24728 3544 24734 3596
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 6362 3516 6368 3528
rect 5951 3488 6368 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 8352 3488 9229 3516
rect 8352 3476 8358 3488
rect 9217 3485 9229 3488
rect 9263 3485 9275 3519
rect 11054 3516 11060 3528
rect 11015 3488 11060 3516
rect 9217 3479 9275 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 12618 3516 12624 3528
rect 12579 3488 12624 3516
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 13078 3516 13084 3528
rect 13039 3488 13084 3516
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 16684 3516 16712 3544
rect 13679 3488 16712 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18524 3516 18552 3544
rect 19150 3516 19156 3528
rect 17920 3488 18552 3516
rect 19111 3488 19156 3516
rect 17920 3476 17926 3488
rect 19150 3476 19156 3488
rect 19208 3476 19214 3528
rect 20070 3476 20076 3528
rect 20128 3516 20134 3528
rect 20990 3516 20996 3528
rect 20128 3488 20996 3516
rect 20128 3476 20134 3488
rect 20990 3476 20996 3488
rect 21048 3476 21054 3528
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3485 21327 3519
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 21269 3479 21327 3485
rect 4338 3448 4344 3460
rect 4299 3420 4344 3448
rect 4338 3408 4344 3420
rect 4396 3408 4402 3460
rect 14274 3448 14280 3460
rect 14235 3420 14280 3448
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 18414 3408 18420 3460
rect 18472 3448 18478 3460
rect 19429 3451 19487 3457
rect 19429 3448 19441 3451
rect 18472 3420 19441 3448
rect 18472 3408 18478 3420
rect 19429 3417 19441 3420
rect 19475 3448 19487 3451
rect 19518 3448 19524 3460
rect 19475 3420 19524 3448
rect 19475 3417 19487 3420
rect 19429 3411 19487 3417
rect 19518 3408 19524 3420
rect 19576 3448 19582 3460
rect 20162 3448 20168 3460
rect 19576 3420 20168 3448
rect 19576 3408 19582 3420
rect 20162 3408 20168 3420
rect 20220 3408 20226 3460
rect 20714 3408 20720 3460
rect 20772 3448 20778 3460
rect 21284 3448 21312 3479
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 21450 3448 21456 3460
rect 20772 3420 21456 3448
rect 20772 3408 20778 3420
rect 21450 3408 21456 3420
rect 21508 3408 21514 3460
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 7098 3380 7104 3392
rect 7059 3352 7104 3380
rect 7098 3340 7104 3352
rect 7156 3380 7162 3392
rect 7282 3380 7288 3392
rect 7156 3352 7288 3380
rect 7156 3340 7162 3352
rect 7282 3340 7288 3352
rect 7340 3380 7346 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 7340 3352 8309 3380
rect 7340 3340 7346 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8846 3380 8852 3392
rect 8807 3352 8852 3380
rect 8297 3343 8355 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 10560 3352 10701 3380
rect 10560 3340 10566 3352
rect 10689 3349 10701 3352
rect 10735 3380 10747 3383
rect 10778 3380 10784 3392
rect 10735 3352 10784 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 10778 3340 10784 3352
rect 10836 3380 10842 3392
rect 11514 3380 11520 3392
rect 10836 3352 11520 3380
rect 10836 3340 10842 3352
rect 11514 3340 11520 3352
rect 11572 3380 11578 3392
rect 12437 3383 12495 3389
rect 12437 3380 12449 3383
rect 11572 3352 12449 3380
rect 11572 3340 11578 3352
rect 12437 3349 12449 3352
rect 12483 3380 12495 3383
rect 12710 3380 12716 3392
rect 12483 3352 12716 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 14001 3383 14059 3389
rect 14001 3380 14013 3383
rect 13780 3352 14013 3380
rect 13780 3340 13786 3352
rect 14001 3349 14013 3352
rect 14047 3380 14059 3383
rect 14826 3380 14832 3392
rect 14047 3352 14832 3380
rect 14047 3349 14059 3352
rect 14001 3343 14059 3349
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1578 3176 1584 3188
rect 1539 3148 1584 3176
rect 1578 3136 1584 3148
rect 1636 3136 1642 3188
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 2317 3179 2375 3185
rect 2317 3176 2329 3179
rect 2188 3148 2329 3176
rect 2188 3136 2194 3148
rect 2317 3145 2329 3148
rect 2363 3145 2375 3179
rect 3142 3176 3148 3188
rect 3103 3148 3148 3176
rect 2317 3139 2375 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 4614 3176 4620 3188
rect 4575 3148 4620 3176
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6512 3148 6561 3176
rect 6512 3136 6518 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8168 3148 8217 3176
rect 8168 3136 8174 3148
rect 8205 3145 8217 3148
rect 8251 3176 8263 3179
rect 8665 3179 8723 3185
rect 8665 3176 8677 3179
rect 8251 3148 8677 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 8665 3145 8677 3148
rect 8711 3145 8723 3179
rect 8665 3139 8723 3145
rect 2777 3111 2835 3117
rect 2777 3077 2789 3111
rect 2823 3108 2835 3111
rect 3510 3108 3516 3120
rect 2823 3080 3516 3108
rect 2823 3077 2835 3080
rect 2777 3071 2835 3077
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 5077 3111 5135 3117
rect 5077 3077 5089 3111
rect 5123 3108 5135 3111
rect 5442 3108 5448 3120
rect 5123 3080 5448 3108
rect 5123 3077 5135 3080
rect 5077 3071 5135 3077
rect 5442 3068 5448 3080
rect 5500 3108 5506 3120
rect 6270 3108 6276 3120
rect 5500 3080 6276 3108
rect 5500 3068 5506 3080
rect 6270 3068 6276 3080
rect 6328 3068 6334 3120
rect 7834 3108 7840 3120
rect 7795 3080 7840 3108
rect 7834 3068 7840 3080
rect 7892 3068 7898 3120
rect 4338 3040 4344 3052
rect 4251 3012 4344 3040
rect 4338 3000 4344 3012
rect 4396 3040 4402 3052
rect 5166 3040 5172 3052
rect 4396 3012 5172 3040
rect 4396 3000 4402 3012
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 5994 3040 6000 3052
rect 5951 3012 6000 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 5994 3000 6000 3012
rect 6052 3040 6058 3052
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 6052 3012 6193 3040
rect 6052 3000 6058 3012
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 6546 3000 6552 3052
rect 6604 3040 6610 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 6604 3012 7297 3040
rect 6604 3000 6610 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 2682 2972 2688 2984
rect 2639 2944 2688 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 4062 2972 4068 2984
rect 3559 2944 4068 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 5350 2972 5356 2984
rect 5311 2944 5356 2972
rect 5350 2932 5356 2944
rect 5408 2972 5414 2984
rect 7009 2975 7067 2981
rect 7009 2972 7021 2975
rect 5408 2944 7021 2972
rect 5408 2932 5414 2944
rect 7009 2941 7021 2944
rect 7055 2972 7067 2975
rect 7098 2972 7104 2984
rect 7055 2944 7104 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7116 2904 7144 2932
rect 7377 2907 7435 2913
rect 7377 2904 7389 2907
rect 7116 2876 7389 2904
rect 7377 2873 7389 2876
rect 7423 2873 7435 2907
rect 8680 2904 8708 3139
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 9582 3176 9588 3188
rect 9272 3148 9588 3176
rect 9272 3136 9278 3148
rect 9582 3136 9588 3148
rect 9640 3176 9646 3188
rect 9769 3179 9827 3185
rect 9769 3176 9781 3179
rect 9640 3148 9781 3176
rect 9640 3136 9646 3148
rect 9769 3145 9781 3148
rect 9815 3145 9827 3179
rect 10042 3176 10048 3188
rect 10003 3148 10048 3176
rect 9769 3139 9827 3145
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10502 3176 10508 3188
rect 10463 3148 10508 3176
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12526 3176 12532 3188
rect 12299 3148 12532 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3176 13510 3188
rect 13504 3148 14136 3176
rect 13504 3136 13510 3148
rect 13078 3108 13084 3120
rect 13039 3080 13084 3108
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 13814 3108 13820 3120
rect 13775 3080 13820 3108
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 14108 3117 14136 3148
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15381 3179 15439 3185
rect 15381 3176 15393 3179
rect 15344 3148 15393 3176
rect 15344 3136 15350 3148
rect 15381 3145 15393 3148
rect 15427 3176 15439 3179
rect 16206 3176 16212 3188
rect 15427 3148 16212 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 17678 3176 17684 3188
rect 17639 3148 17684 3176
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 18046 3136 18052 3188
rect 18104 3176 18110 3188
rect 19797 3179 19855 3185
rect 19797 3176 19809 3179
rect 18104 3148 19809 3176
rect 18104 3136 18110 3148
rect 19797 3145 19809 3148
rect 19843 3176 19855 3179
rect 19978 3176 19984 3188
rect 19843 3148 19984 3176
rect 19843 3145 19855 3148
rect 19797 3139 19855 3145
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 21082 3136 21088 3188
rect 21140 3176 21146 3188
rect 21542 3176 21548 3188
rect 21140 3148 21548 3176
rect 21140 3136 21146 3148
rect 21542 3136 21548 3148
rect 21600 3176 21606 3188
rect 21637 3179 21695 3185
rect 21637 3176 21649 3179
rect 21600 3148 21649 3176
rect 21600 3136 21606 3148
rect 21637 3145 21649 3148
rect 21683 3145 21695 3179
rect 24670 3176 24676 3188
rect 24631 3148 24676 3176
rect 21637 3139 21695 3145
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 25406 3176 25412 3188
rect 25367 3148 25412 3176
rect 25406 3136 25412 3148
rect 25464 3136 25470 3188
rect 14093 3111 14151 3117
rect 14093 3077 14105 3111
rect 14139 3077 14151 3111
rect 14093 3071 14151 3077
rect 23477 3111 23535 3117
rect 23477 3077 23489 3111
rect 23523 3108 23535 3111
rect 23842 3108 23848 3120
rect 23523 3080 23848 3108
rect 23523 3077 23535 3080
rect 23477 3071 23535 3077
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 8846 3040 8852 3052
rect 8807 3012 8852 3040
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 10686 3040 10692 3052
rect 10647 3012 10692 3040
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11698 3040 11704 3052
rect 11379 3012 11704 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11698 3000 11704 3012
rect 11756 3040 11762 3052
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 11756 3012 12541 3040
rect 11756 3000 11762 3012
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 13832 2972 13860 3068
rect 14734 3040 14740 3052
rect 14695 3012 14740 3040
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17000 3012 17417 3040
rect 17000 3000 17006 3012
rect 17405 3009 17417 3012
rect 17451 3040 17463 3043
rect 17451 3012 18920 3040
rect 17451 3009 17463 3012
rect 17405 3003 17463 3009
rect 18892 2984 18920 3012
rect 19150 3000 19156 3052
rect 19208 3040 19214 3052
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 19208 3012 20453 3040
rect 19208 3000 19214 3012
rect 20441 3009 20453 3012
rect 20487 3040 20499 3043
rect 22097 3043 22155 3049
rect 22097 3040 22109 3043
rect 20487 3012 22109 3040
rect 20487 3009 20499 3012
rect 20441 3003 20499 3009
rect 22097 3009 22109 3012
rect 22143 3009 22155 3043
rect 22922 3040 22928 3052
rect 22097 3003 22155 3009
rect 22480 3012 22928 3040
rect 22480 2984 22508 3012
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 23014 3000 23020 3052
rect 23072 3040 23078 3052
rect 24029 3043 24087 3049
rect 24029 3040 24041 3043
rect 23072 3012 24041 3040
rect 23072 3000 23078 3012
rect 24029 3009 24041 3012
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13832 2944 14013 2972
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 14090 2932 14096 2984
rect 14148 2972 14154 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14148 2944 14289 2972
rect 14148 2932 14154 2944
rect 14277 2941 14289 2944
rect 14323 2972 14335 2975
rect 14550 2972 14556 2984
rect 14323 2944 14556 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 15746 2972 15752 2984
rect 15707 2944 15752 2972
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15988 2944 16037 2972
rect 15988 2932 15994 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16025 2935 16083 2941
rect 16206 2932 16212 2984
rect 16264 2972 16270 2984
rect 16393 2975 16451 2981
rect 16393 2972 16405 2975
rect 16264 2944 16405 2972
rect 16264 2932 16270 2944
rect 16393 2941 16405 2944
rect 16439 2941 16451 2975
rect 16393 2935 16451 2941
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 16632 2944 16773 2972
rect 16632 2932 16638 2944
rect 16761 2941 16773 2944
rect 16807 2941 16819 2975
rect 18046 2972 18052 2984
rect 17959 2944 18052 2972
rect 16761 2935 16819 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18472 2944 18521 2972
rect 18472 2932 18478 2944
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 18874 2972 18880 2984
rect 18835 2944 18880 2972
rect 18509 2935 18567 2941
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 19242 2972 19248 2984
rect 19203 2944 19248 2972
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 22462 2972 22468 2984
rect 22375 2944 22468 2972
rect 22462 2932 22468 2944
rect 22520 2932 22526 2984
rect 22830 2932 22836 2984
rect 22888 2972 22894 2984
rect 25225 2975 25283 2981
rect 22888 2944 23336 2972
rect 22888 2932 22894 2944
rect 9170 2907 9228 2913
rect 9170 2904 9182 2907
rect 8680 2876 9182 2904
rect 7377 2867 7435 2873
rect 9170 2873 9182 2876
rect 9216 2873 9228 2907
rect 9170 2867 9228 2873
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 12621 2907 12679 2913
rect 10836 2876 10881 2904
rect 10836 2864 10842 2876
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 12802 2904 12808 2916
rect 12667 2876 12808 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 15764 2904 15792 2932
rect 18064 2904 18092 2932
rect 15764 2876 18092 2904
rect 20762 2907 20820 2913
rect 20762 2873 20774 2907
rect 20808 2904 20820 2907
rect 20898 2904 20904 2916
rect 20808 2876 20904 2904
rect 20808 2873 20820 2876
rect 20762 2867 20820 2873
rect 11698 2836 11704 2848
rect 11659 2808 11704 2836
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 16758 2836 16764 2848
rect 16719 2808 16764 2836
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 19242 2836 19248 2848
rect 19203 2808 19248 2836
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 19426 2796 19432 2848
rect 19484 2836 19490 2848
rect 20257 2839 20315 2845
rect 20257 2836 20269 2839
rect 19484 2808 20269 2836
rect 19484 2796 19490 2808
rect 20257 2805 20269 2808
rect 20303 2836 20315 2839
rect 20777 2836 20805 2867
rect 20898 2864 20904 2876
rect 20956 2864 20962 2916
rect 22738 2904 22744 2916
rect 22480 2876 22744 2904
rect 20303 2808 20805 2836
rect 21361 2839 21419 2845
rect 20303 2805 20315 2808
rect 20257 2799 20315 2805
rect 21361 2805 21373 2839
rect 21407 2836 21419 2839
rect 22480 2836 22508 2876
rect 22738 2864 22744 2876
rect 22796 2904 22802 2916
rect 23308 2904 23336 2944
rect 25225 2941 25237 2975
rect 25271 2972 25283 2975
rect 25682 2972 25688 2984
rect 25271 2944 25688 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 25682 2932 25688 2944
rect 25740 2972 25746 2984
rect 25777 2975 25835 2981
rect 25777 2972 25789 2975
rect 25740 2944 25789 2972
rect 25740 2932 25746 2944
rect 25777 2941 25789 2944
rect 25823 2941 25835 2975
rect 25777 2935 25835 2941
rect 23750 2904 23756 2916
rect 22796 2876 23152 2904
rect 23308 2876 23756 2904
rect 22796 2864 22802 2876
rect 22646 2836 22652 2848
rect 21407 2808 22508 2836
rect 22607 2808 22652 2836
rect 21407 2805 21419 2808
rect 21361 2799 21419 2805
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 23124 2845 23152 2876
rect 23750 2864 23756 2876
rect 23808 2864 23814 2916
rect 23842 2864 23848 2916
rect 23900 2904 23906 2916
rect 23900 2876 23945 2904
rect 23900 2864 23906 2876
rect 23109 2839 23167 2845
rect 23109 2805 23121 2839
rect 23155 2836 23167 2839
rect 23382 2836 23388 2848
rect 23155 2808 23388 2836
rect 23155 2805 23167 2808
rect 23109 2799 23167 2805
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2498 2632 2504 2644
rect 2459 2604 2504 2632
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 5166 2632 5172 2644
rect 5127 2604 5172 2632
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 6362 2632 6368 2644
rect 5920 2604 6368 2632
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 4706 2564 4712 2576
rect 2087 2536 4712 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 2056 2496 2084 2527
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 1443 2468 2084 2496
rect 4249 2499 4307 2505
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4798 2496 4804 2508
rect 4295 2468 4804 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5920 2505 5948 2604
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 6733 2635 6791 2641
rect 6733 2601 6745 2635
rect 6779 2632 6791 2635
rect 6822 2632 6828 2644
rect 6779 2604 6828 2632
rect 6779 2601 6791 2604
rect 6733 2595 6791 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7239 2635 7297 2641
rect 7239 2601 7251 2635
rect 7285 2632 7297 2635
rect 8754 2632 8760 2644
rect 7285 2604 8760 2632
rect 7285 2601 7297 2604
rect 7239 2595 7297 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 9456 2604 9505 2632
rect 9456 2592 9462 2604
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 9493 2595 9551 2601
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 10686 2632 10692 2644
rect 10459 2604 10692 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 8202 2564 8208 2576
rect 8163 2536 8208 2564
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 8352 2536 8397 2564
rect 8352 2524 8358 2536
rect 5905 2499 5963 2505
rect 5905 2465 5917 2499
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 7136 2499 7194 2505
rect 7136 2496 7148 2499
rect 7055 2468 7148 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 7136 2465 7148 2468
rect 7182 2465 7194 2499
rect 7136 2459 7194 2465
rect 8849 2499 8907 2505
rect 8849 2465 8861 2499
rect 8895 2496 8907 2499
rect 9490 2496 9496 2508
rect 8895 2468 9496 2496
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10428 2496 10456 2595
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11698 2632 11704 2644
rect 11164 2604 11704 2632
rect 11164 2576 11192 2604
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 13630 2632 13636 2644
rect 12483 2604 13636 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14090 2632 14096 2644
rect 14051 2604 14096 2632
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15746 2632 15752 2644
rect 15335 2604 15752 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 16577 2635 16635 2641
rect 16577 2601 16589 2635
rect 16623 2632 16635 2635
rect 16666 2632 16672 2644
rect 16623 2604 16672 2632
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 17862 2632 17868 2644
rect 17819 2604 17868 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 19426 2632 19432 2644
rect 18800 2604 19432 2632
rect 10781 2567 10839 2573
rect 10781 2533 10793 2567
rect 10827 2564 10839 2567
rect 11057 2567 11115 2573
rect 11057 2564 11069 2567
rect 10827 2536 11069 2564
rect 10827 2533 10839 2536
rect 10781 2527 10839 2533
rect 11057 2533 11069 2536
rect 11103 2564 11115 2567
rect 11146 2564 11152 2576
rect 11103 2536 11152 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11606 2564 11612 2576
rect 11567 2536 11612 2564
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 11716 2564 11744 2592
rect 18800 2576 18828 2604
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19613 2635 19671 2641
rect 19613 2632 19625 2635
rect 19576 2604 19625 2632
rect 19576 2592 19582 2604
rect 19613 2601 19625 2604
rect 19659 2601 19671 2635
rect 20990 2632 20996 2644
rect 20951 2604 20996 2632
rect 19613 2595 19671 2601
rect 20990 2592 20996 2604
rect 21048 2592 21054 2644
rect 22462 2592 22468 2644
rect 22520 2632 22526 2644
rect 22557 2635 22615 2641
rect 22557 2632 22569 2635
rect 22520 2604 22569 2632
rect 22520 2592 22526 2604
rect 22557 2601 22569 2604
rect 22603 2601 22615 2635
rect 23750 2632 23756 2644
rect 23711 2604 23756 2632
rect 22557 2595 22615 2601
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 25406 2632 25412 2644
rect 25367 2604 25412 2632
rect 25406 2592 25412 2604
rect 25464 2592 25470 2644
rect 12621 2567 12679 2573
rect 12621 2564 12633 2567
rect 11716 2536 12633 2564
rect 12621 2533 12633 2536
rect 12667 2533 12679 2567
rect 12621 2527 12679 2533
rect 17954 2524 17960 2576
rect 18012 2564 18018 2576
rect 18782 2573 18788 2576
rect 18141 2567 18199 2573
rect 18141 2564 18153 2567
rect 18012 2536 18153 2564
rect 18012 2524 18018 2536
rect 18141 2533 18153 2536
rect 18187 2564 18199 2567
rect 18779 2564 18788 2573
rect 18187 2536 18788 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 18779 2527 18788 2536
rect 18782 2524 18788 2527
rect 18840 2524 18846 2576
rect 21361 2567 21419 2573
rect 21361 2564 21373 2567
rect 20548 2536 21373 2564
rect 12710 2496 12716 2508
rect 9907 2468 10456 2496
rect 12671 2468 12716 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 14274 2496 14280 2508
rect 14235 2468 14280 2496
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 15562 2496 15568 2508
rect 15523 2468 15568 2496
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 20548 2505 20576 2536
rect 21361 2533 21373 2536
rect 21407 2533 21419 2567
rect 22186 2564 22192 2576
rect 22147 2536 22192 2564
rect 21361 2527 21419 2533
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 23658 2564 23664 2576
rect 22848 2536 23664 2564
rect 22848 2505 22876 2536
rect 23658 2524 23664 2536
rect 23716 2524 23722 2576
rect 23842 2524 23848 2576
rect 23900 2564 23906 2576
rect 24029 2567 24087 2573
rect 24029 2564 24041 2567
rect 23900 2536 24041 2564
rect 23900 2524 23906 2536
rect 24029 2533 24041 2536
rect 24075 2533 24087 2567
rect 24029 2527 24087 2533
rect 17313 2499 17371 2505
rect 17313 2465 17325 2499
rect 17359 2496 17371 2499
rect 19337 2499 19395 2505
rect 19337 2496 19349 2499
rect 17359 2468 19349 2496
rect 17359 2465 17371 2468
rect 17313 2459 17371 2465
rect 19337 2465 19349 2468
rect 19383 2496 19395 2499
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19383 2468 19993 2496
rect 19383 2465 19395 2468
rect 19337 2459 19395 2465
rect 19981 2465 19993 2468
rect 20027 2496 20039 2499
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20027 2468 20545 2496
rect 20027 2465 20039 2468
rect 19981 2459 20039 2465
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 24121 2499 24179 2505
rect 24121 2496 24133 2499
rect 23532 2468 24133 2496
rect 23532 2456 23538 2468
rect 24121 2465 24133 2468
rect 24167 2496 24179 2499
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24167 2468 25053 2496
rect 24167 2465 24179 2468
rect 24121 2459 24179 2465
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 25660 2499 25718 2505
rect 25660 2465 25672 2499
rect 25706 2496 25718 2499
rect 26142 2496 26148 2508
rect 25706 2468 26148 2496
rect 25706 2465 25718 2468
rect 25660 2459 25718 2465
rect 26142 2456 26148 2468
rect 26200 2456 26206 2508
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 6043 2400 7941 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 7929 2397 7941 2400
rect 7975 2428 7987 2431
rect 8294 2428 8300 2440
rect 7975 2400 8300 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9214 2428 9220 2440
rect 9175 2400 9220 2428
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 10962 2428 10968 2440
rect 10875 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2428 11026 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11020 2400 11897 2428
rect 11020 2388 11026 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 15286 2388 15292 2440
rect 15344 2428 15350 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15344 2400 16129 2428
rect 15344 2388 15350 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 17402 2428 17408 2440
rect 17363 2400 17408 2428
rect 16117 2391 16175 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2428 18475 2431
rect 19242 2428 19248 2440
rect 18463 2400 19248 2428
rect 18463 2397 18475 2400
rect 18417 2391 18475 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 21266 2428 21272 2440
rect 21227 2400 21272 2428
rect 21266 2388 21272 2400
rect 21324 2388 21330 2440
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 21545 2431 21603 2437
rect 21545 2428 21557 2431
rect 21508 2400 21557 2428
rect 21508 2388 21514 2400
rect 21545 2397 21557 2400
rect 21591 2397 21603 2431
rect 21545 2391 21603 2397
rect 3602 2320 3608 2372
rect 3660 2360 3666 2372
rect 7009 2363 7067 2369
rect 7009 2360 7021 2363
rect 3660 2332 7021 2360
rect 3660 2320 3666 2332
rect 7009 2329 7021 2332
rect 7055 2360 7067 2363
rect 7561 2363 7619 2369
rect 7561 2360 7573 2363
rect 7055 2332 7573 2360
rect 7055 2329 7067 2332
rect 7009 2323 7067 2329
rect 7561 2329 7573 2332
rect 7607 2329 7619 2363
rect 7561 2323 7619 2329
rect 24854 2320 24860 2372
rect 24912 2360 24918 2372
rect 25731 2363 25789 2369
rect 25731 2360 25743 2363
rect 24912 2332 25743 2360
rect 24912 2320 24918 2332
rect 25731 2329 25743 2332
rect 25777 2329 25789 2363
rect 25731 2323 25789 2329
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 4430 2292 4436 2304
rect 4391 2264 4436 2292
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 10045 2295 10103 2301
rect 10045 2261 10057 2295
rect 10091 2292 10103 2295
rect 10226 2292 10232 2304
rect 10091 2264 10232 2292
rect 10091 2261 10103 2264
rect 10045 2255 10103 2261
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 14458 2292 14464 2304
rect 14419 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 23014 2292 23020 2304
rect 22975 2264 23020 2292
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 26142 2292 26148 2304
rect 26103 2264 26148 2292
rect 26142 2252 26148 2264
rect 26200 2252 26206 2304
rect 26418 2292 26424 2304
rect 26379 2264 26424 2292
rect 26418 2252 26424 2264
rect 26476 2252 26482 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 2314 1232 2320 1284
rect 2372 1272 2378 1284
rect 3602 1272 3608 1284
rect 2372 1244 3608 1272
rect 2372 1232 2378 1244
rect 3602 1232 3608 1244
rect 3660 1232 3666 1284
rect 7190 552 7196 604
rect 7248 592 7254 604
rect 7926 592 7932 604
rect 7248 564 7932 592
rect 7248 552 7254 564
rect 7926 552 7932 564
rect 7984 552 7990 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 24768 23808 24820 23860
rect 13544 23715 13596 23724
rect 13544 23681 13553 23715
rect 13553 23681 13587 23715
rect 13587 23681 13596 23715
rect 13544 23672 13596 23681
rect 1400 23647 1452 23656
rect 1400 23613 1444 23647
rect 1444 23613 1452 23647
rect 1400 23604 1452 23613
rect 24768 23604 24820 23656
rect 1768 23468 1820 23520
rect 13360 23468 13412 23520
rect 23480 23468 23532 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 24676 22720 24728 22772
rect 24676 22559 24728 22568
rect 24676 22525 24694 22559
rect 24694 22525 24728 22559
rect 24676 22516 24728 22525
rect 23664 22380 23716 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 13452 21403 13504 21412
rect 13452 21369 13461 21403
rect 13461 21369 13495 21403
rect 13495 21369 13504 21403
rect 13452 21360 13504 21369
rect 13544 21292 13596 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1860 20952 1912 21004
rect 2688 20952 2740 21004
rect 2780 20952 2832 21004
rect 24676 20995 24728 21004
rect 24676 20961 24694 20995
rect 24694 20961 24728 20995
rect 24676 20952 24728 20961
rect 2136 20816 2188 20868
rect 3424 20748 3476 20800
rect 23480 20748 23532 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2780 20544 2832 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 2044 20476 2096 20528
rect 1584 20340 1636 20392
rect 1584 20204 1636 20256
rect 1860 20247 1912 20256
rect 1860 20213 1869 20247
rect 1869 20213 1903 20247
rect 1903 20213 1912 20247
rect 1860 20204 1912 20213
rect 3148 20272 3200 20324
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1400 19907 1452 19916
rect 1400 19873 1444 19907
rect 1444 19873 1452 19907
rect 1400 19864 1452 19873
rect 4344 19864 4396 19916
rect 2504 19796 2556 19848
rect 2320 19660 2372 19712
rect 4988 19660 5040 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1400 19456 1452 19508
rect 1400 19295 1452 19304
rect 1400 19261 1444 19295
rect 1444 19261 1452 19295
rect 1400 19252 1452 19261
rect 2964 19295 3016 19304
rect 2964 19261 2973 19295
rect 2973 19261 3007 19295
rect 3007 19261 3016 19295
rect 2964 19252 3016 19261
rect 3608 19252 3660 19304
rect 5080 19252 5132 19304
rect 2136 19184 2188 19236
rect 2412 19116 2464 19168
rect 3148 19116 3200 19168
rect 4344 19159 4396 19168
rect 4344 19125 4353 19159
rect 4353 19125 4387 19159
rect 4387 19125 4396 19159
rect 4344 19116 4396 19125
rect 4528 19116 4580 19168
rect 5080 19116 5132 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1952 18776 2004 18828
rect 2688 18776 2740 18828
rect 3332 18776 3384 18828
rect 5172 18819 5224 18828
rect 5172 18785 5190 18819
rect 5190 18785 5224 18819
rect 5172 18776 5224 18785
rect 5448 18708 5500 18760
rect 3884 18640 3936 18692
rect 1676 18572 1728 18624
rect 2136 18572 2188 18624
rect 4160 18572 4212 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2596 18368 2648 18420
rect 3332 18411 3384 18420
rect 3332 18377 3341 18411
rect 3341 18377 3375 18411
rect 3375 18377 3384 18411
rect 3332 18368 3384 18377
rect 1308 18300 1360 18352
rect 1216 18164 1268 18216
rect 2596 18164 2648 18216
rect 8116 18300 8168 18352
rect 5172 18275 5224 18284
rect 5172 18241 5181 18275
rect 5181 18241 5215 18275
rect 5215 18241 5224 18275
rect 5172 18232 5224 18241
rect 8576 18232 8628 18284
rect 6000 18096 6052 18148
rect 1584 18028 1636 18080
rect 2596 18028 2648 18080
rect 3516 18028 3568 18080
rect 3792 18028 3844 18080
rect 4436 18028 4488 18080
rect 7472 18139 7524 18148
rect 7472 18105 7481 18139
rect 7481 18105 7515 18139
rect 7515 18105 7524 18139
rect 7472 18096 7524 18105
rect 6184 18028 6236 18080
rect 6920 18028 6972 18080
rect 7656 18028 7708 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 1400 17620 1452 17672
rect 4804 17688 4856 17740
rect 6276 17688 6328 17740
rect 8944 17688 8996 17740
rect 9956 17688 10008 17740
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 2228 17620 2280 17629
rect 6460 17620 6512 17672
rect 10968 17620 11020 17672
rect 2688 17484 2740 17536
rect 3700 17484 3752 17536
rect 4712 17484 4764 17536
rect 6092 17484 6144 17536
rect 8300 17484 8352 17536
rect 9864 17484 9916 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 6276 17280 6328 17332
rect 1400 17144 1452 17196
rect 6920 17212 6972 17264
rect 3240 17119 3292 17128
rect 3240 17085 3284 17119
rect 3284 17085 3292 17119
rect 3240 17076 3292 17085
rect 2964 17008 3016 17060
rect 7380 17008 7432 17060
rect 10048 17076 10100 17128
rect 11152 17076 11204 17128
rect 13084 17119 13136 17128
rect 13084 17085 13102 17119
rect 13102 17085 13136 17119
rect 13084 17076 13136 17085
rect 14740 17076 14792 17128
rect 9036 17051 9088 17060
rect 9036 17017 9045 17051
rect 9045 17017 9079 17051
rect 9079 17017 9088 17051
rect 9036 17008 9088 17017
rect 10876 17008 10928 17060
rect 1860 16940 1912 16992
rect 3976 16940 4028 16992
rect 4804 16940 4856 16992
rect 4896 16940 4948 16992
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 7472 16940 7524 16992
rect 8392 16940 8444 16992
rect 8944 16940 8996 16992
rect 9956 16940 10008 16992
rect 11244 16940 11296 16992
rect 12808 16940 12860 16992
rect 16304 16940 16356 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1952 16736 2004 16788
rect 2044 16736 2096 16788
rect 4712 16779 4764 16788
rect 4712 16745 4721 16779
rect 4721 16745 4755 16779
rect 4755 16745 4764 16779
rect 4712 16736 4764 16745
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 13268 16779 13320 16788
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 15936 16736 15988 16788
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 2688 16668 2740 16720
rect 8208 16668 8260 16720
rect 2044 16532 2096 16584
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 4344 16600 4396 16652
rect 4620 16532 4672 16584
rect 5264 16600 5316 16652
rect 6828 16600 6880 16652
rect 8484 16643 8536 16652
rect 8484 16609 8528 16643
rect 8528 16609 8536 16643
rect 8484 16600 8536 16609
rect 9588 16600 9640 16652
rect 10140 16600 10192 16652
rect 11888 16600 11940 16652
rect 12348 16600 12400 16652
rect 16120 16668 16172 16720
rect 5540 16532 5592 16584
rect 12256 16532 12308 16584
rect 13636 16600 13688 16652
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 16948 16600 17000 16652
rect 6736 16439 6788 16448
rect 6736 16405 6745 16439
rect 6745 16405 6779 16439
rect 6779 16405 6788 16439
rect 6736 16396 6788 16405
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 14372 16396 14424 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2688 16192 2740 16244
rect 4712 16124 4764 16176
rect 2872 16099 2924 16108
rect 2872 16065 2881 16099
rect 2881 16065 2915 16099
rect 2915 16065 2924 16099
rect 2872 16056 2924 16065
rect 5080 16099 5132 16108
rect 5080 16065 5089 16099
rect 5089 16065 5123 16099
rect 5123 16065 5132 16099
rect 5080 16056 5132 16065
rect 4620 15988 4672 16040
rect 2688 15963 2740 15972
rect 2688 15929 2697 15963
rect 2697 15929 2731 15963
rect 2731 15929 2740 15963
rect 2688 15920 2740 15929
rect 1400 15852 1452 15904
rect 8484 16192 8536 16244
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 24768 16192 24820 16244
rect 9588 16056 9640 16108
rect 6276 15920 6328 15972
rect 5632 15852 5684 15904
rect 5724 15852 5776 15904
rect 6552 15852 6604 15904
rect 6828 15852 6880 15904
rect 7288 15852 7340 15904
rect 8116 16031 8168 16040
rect 8116 15997 8160 16031
rect 8160 15997 8168 16031
rect 8116 15988 8168 15997
rect 9128 16031 9180 16040
rect 9128 15997 9137 16031
rect 9137 15997 9171 16031
rect 9171 15997 9180 16031
rect 9128 15988 9180 15997
rect 12440 16056 12492 16108
rect 14648 16099 14700 16108
rect 11336 15988 11388 16040
rect 11520 15988 11572 16040
rect 12164 15988 12216 16040
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 14280 16031 14332 16040
rect 11428 15963 11480 15972
rect 11428 15929 11437 15963
rect 11437 15929 11471 15963
rect 11471 15929 11480 15963
rect 11428 15920 11480 15929
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 14372 15988 14424 16040
rect 13820 15920 13872 15972
rect 16856 15963 16908 15972
rect 16856 15929 16865 15963
rect 16865 15929 16899 15963
rect 16899 15929 16908 15963
rect 16856 15920 16908 15929
rect 7932 15852 7984 15904
rect 8116 15852 8168 15904
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 11888 15852 11940 15904
rect 12624 15852 12676 15904
rect 14280 15852 14332 15904
rect 14464 15852 14516 15904
rect 15292 15852 15344 15904
rect 15752 15852 15804 15904
rect 16948 15852 17000 15904
rect 18512 15852 18564 15904
rect 24768 15988 24820 16040
rect 18788 15852 18840 15904
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 23480 15852 23532 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1216 15648 1268 15700
rect 1492 15648 1544 15700
rect 2044 15648 2096 15700
rect 2688 15648 2740 15700
rect 2964 15648 3016 15700
rect 2320 15623 2372 15632
rect 2320 15589 2329 15623
rect 2329 15589 2363 15623
rect 2363 15589 2372 15623
rect 2320 15580 2372 15589
rect 2872 15623 2924 15632
rect 2872 15589 2881 15623
rect 2881 15589 2915 15623
rect 2915 15589 2924 15623
rect 5172 15648 5224 15700
rect 5632 15648 5684 15700
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 11796 15691 11848 15700
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 2872 15580 2924 15589
rect 6092 15623 6144 15632
rect 6092 15589 6101 15623
rect 6101 15589 6135 15623
rect 6135 15589 6144 15623
rect 6092 15580 6144 15589
rect 6276 15580 6328 15632
rect 10232 15580 10284 15632
rect 13820 15623 13872 15632
rect 13820 15589 13829 15623
rect 13829 15589 13863 15623
rect 13863 15589 13872 15623
rect 13820 15580 13872 15589
rect 15844 15580 15896 15632
rect 17776 15623 17828 15632
rect 17776 15589 17785 15623
rect 17785 15589 17819 15623
rect 17819 15589 17828 15623
rect 17776 15580 17828 15589
rect 17868 15623 17920 15632
rect 17868 15589 17877 15623
rect 17877 15589 17911 15623
rect 17911 15589 17920 15623
rect 17868 15580 17920 15589
rect 7840 15512 7892 15564
rect 11888 15555 11940 15564
rect 2412 15444 2464 15496
rect 4068 15376 4120 15428
rect 4252 15444 4304 15496
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 6920 15444 6972 15496
rect 8024 15376 8076 15428
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12256 15512 12308 15521
rect 12440 15512 12492 15564
rect 9680 15444 9732 15496
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 16212 15487 16264 15496
rect 16212 15453 16221 15487
rect 16221 15453 16255 15487
rect 16255 15453 16264 15487
rect 16212 15444 16264 15453
rect 16488 15444 16540 15496
rect 16856 15487 16908 15496
rect 16856 15453 16865 15487
rect 16865 15453 16899 15487
rect 16899 15453 16908 15487
rect 16856 15444 16908 15453
rect 20076 15444 20128 15496
rect 21732 15444 21784 15496
rect 10140 15376 10192 15428
rect 11060 15376 11112 15428
rect 11336 15308 11388 15360
rect 13636 15376 13688 15428
rect 13912 15376 13964 15428
rect 12716 15308 12768 15360
rect 14556 15308 14608 15360
rect 15844 15308 15896 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2780 15104 2832 15156
rect 6092 15104 6144 15156
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 12256 15147 12308 15156
rect 12256 15113 12265 15147
rect 12265 15113 12299 15147
rect 12299 15113 12308 15147
rect 12256 15104 12308 15113
rect 13636 15147 13688 15156
rect 13636 15113 13645 15147
rect 13645 15113 13679 15147
rect 13679 15113 13688 15147
rect 13636 15104 13688 15113
rect 15292 15104 15344 15156
rect 17776 15104 17828 15156
rect 2320 15079 2372 15088
rect 2320 15045 2329 15079
rect 2329 15045 2363 15079
rect 2363 15045 2372 15079
rect 2320 15036 2372 15045
rect 2964 15036 3016 15088
rect 2872 14968 2924 15020
rect 3240 14832 3292 14884
rect 4436 14968 4488 15020
rect 6920 15011 6972 15020
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 7196 15011 7248 15020
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 9588 14968 9640 15020
rect 11244 14968 11296 15020
rect 2412 14764 2464 14816
rect 5080 14832 5132 14884
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 3884 14764 3936 14816
rect 6092 14807 6144 14816
rect 6092 14773 6101 14807
rect 6101 14773 6135 14807
rect 6135 14773 6144 14807
rect 6092 14764 6144 14773
rect 6276 14764 6328 14816
rect 7840 14764 7892 14816
rect 9496 14832 9548 14884
rect 11060 14832 11112 14884
rect 12716 14968 12768 15020
rect 14556 14968 14608 15020
rect 17868 14968 17920 15020
rect 12256 14832 12308 14884
rect 12716 14875 12768 14884
rect 12716 14841 12725 14875
rect 12725 14841 12759 14875
rect 12759 14841 12768 14875
rect 12716 14832 12768 14841
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 14372 14832 14424 14884
rect 14832 14875 14884 14884
rect 14832 14841 14841 14875
rect 14841 14841 14875 14875
rect 14875 14841 14884 14875
rect 14832 14832 14884 14841
rect 15384 14764 15436 14816
rect 15844 14875 15896 14884
rect 15844 14841 15853 14875
rect 15853 14841 15887 14875
rect 15887 14841 15896 14875
rect 15844 14832 15896 14841
rect 20168 15036 20220 15088
rect 20720 14900 20772 14952
rect 23940 14900 23992 14952
rect 18328 14764 18380 14816
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 18972 14764 19024 14816
rect 20260 14764 20312 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 21456 14764 21508 14816
rect 22284 14807 22336 14816
rect 22284 14773 22293 14807
rect 22293 14773 22327 14807
rect 22327 14773 22336 14807
rect 22284 14764 22336 14773
rect 24124 14764 24176 14816
rect 24952 14764 25004 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2228 14560 2280 14612
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 3240 14603 3292 14612
rect 3240 14569 3249 14603
rect 3249 14569 3283 14603
rect 3283 14569 3292 14603
rect 3240 14560 3292 14569
rect 4068 14560 4120 14612
rect 6092 14560 6144 14612
rect 8024 14560 8076 14612
rect 4252 14535 4304 14544
rect 1860 14424 1912 14476
rect 4252 14501 4261 14535
rect 4261 14501 4295 14535
rect 4295 14501 4304 14535
rect 4252 14492 4304 14501
rect 4804 14535 4856 14544
rect 4804 14501 4813 14535
rect 4813 14501 4847 14535
rect 4847 14501 4856 14535
rect 4804 14492 4856 14501
rect 6276 14492 6328 14544
rect 8668 14492 8720 14544
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 8484 14424 8536 14476
rect 9588 14560 9640 14612
rect 12256 14560 12308 14612
rect 14372 14603 14424 14612
rect 14372 14569 14381 14603
rect 14381 14569 14415 14603
rect 14415 14569 14424 14603
rect 14372 14560 14424 14569
rect 15292 14560 15344 14612
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 10232 14492 10284 14544
rect 13544 14535 13596 14544
rect 13544 14501 13547 14535
rect 13547 14501 13581 14535
rect 13581 14501 13596 14535
rect 13544 14492 13596 14501
rect 16488 14535 16540 14544
rect 16488 14501 16497 14535
rect 16497 14501 16531 14535
rect 16531 14501 16540 14535
rect 16488 14492 16540 14501
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 10876 14424 10928 14476
rect 11428 14467 11480 14476
rect 11428 14433 11437 14467
rect 11437 14433 11471 14467
rect 11471 14433 11480 14467
rect 11428 14424 11480 14433
rect 13268 14424 13320 14476
rect 15476 14424 15528 14476
rect 17408 14424 17460 14476
rect 18144 14424 18196 14476
rect 19524 14467 19576 14476
rect 19524 14433 19568 14467
rect 19568 14433 19576 14467
rect 19524 14424 19576 14433
rect 20904 14467 20956 14476
rect 20904 14433 20948 14467
rect 20948 14433 20956 14467
rect 20904 14424 20956 14433
rect 22008 14467 22060 14476
rect 22008 14433 22026 14467
rect 22026 14433 22060 14467
rect 22008 14424 22060 14433
rect 23940 14467 23992 14476
rect 23940 14433 23984 14467
rect 23984 14433 23992 14467
rect 23940 14424 23992 14433
rect 24860 14424 24912 14476
rect 2320 14356 2372 14408
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 6644 14356 6696 14408
rect 9312 14356 9364 14408
rect 16856 14356 16908 14408
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17040 14356 17092 14365
rect 22192 14356 22244 14408
rect 10140 14288 10192 14340
rect 5080 14220 5132 14272
rect 10692 14220 10744 14272
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 12992 14263 13044 14272
rect 12992 14229 13001 14263
rect 13001 14229 13035 14263
rect 13035 14229 13044 14263
rect 12992 14220 13044 14229
rect 20720 14220 20772 14272
rect 21548 14220 21600 14272
rect 22008 14220 22060 14272
rect 23204 14220 23256 14272
rect 25320 14220 25372 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 3240 14016 3292 14068
rect 4252 14016 4304 14068
rect 7012 14016 7064 14068
rect 8300 14016 8352 14068
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 11244 14016 11296 14068
rect 11428 14016 11480 14068
rect 12716 14016 12768 14068
rect 15476 14016 15528 14068
rect 16488 14016 16540 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 19616 14016 19668 14068
rect 20904 14016 20956 14068
rect 21364 14016 21416 14068
rect 21916 14016 21968 14068
rect 24860 14016 24912 14068
rect 1860 13948 1912 14000
rect 10600 13991 10652 14000
rect 10600 13957 10609 13991
rect 10609 13957 10643 13991
rect 10643 13957 10652 13991
rect 10600 13948 10652 13957
rect 10876 13991 10928 14000
rect 10876 13957 10885 13991
rect 10885 13957 10919 13991
rect 10919 13957 10928 13991
rect 10876 13948 10928 13957
rect 13268 13948 13320 14000
rect 16580 13948 16632 14000
rect 18144 13948 18196 14000
rect 19524 13948 19576 14000
rect 24216 13948 24268 14000
rect 2228 13880 2280 13932
rect 4068 13880 4120 13932
rect 2964 13812 3016 13864
rect 1400 13744 1452 13796
rect 1860 13744 1912 13796
rect 2320 13744 2372 13796
rect 5080 13880 5132 13932
rect 5448 13880 5500 13932
rect 7196 13880 7248 13932
rect 9772 13880 9824 13932
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 12992 13880 13044 13932
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 23756 13880 23808 13932
rect 6828 13855 6880 13864
rect 6828 13821 6833 13855
rect 6833 13821 6867 13855
rect 6867 13821 6880 13855
rect 6828 13812 6880 13821
rect 8576 13855 8628 13864
rect 8576 13821 8620 13855
rect 8620 13821 8628 13855
rect 8576 13812 8628 13821
rect 2044 13676 2096 13728
rect 4068 13676 4120 13728
rect 5540 13744 5592 13796
rect 6276 13787 6328 13796
rect 6276 13753 6285 13787
rect 6285 13753 6319 13787
rect 6319 13753 6328 13787
rect 6276 13744 6328 13753
rect 10232 13744 10284 13796
rect 11428 13719 11480 13728
rect 11428 13685 11437 13719
rect 11437 13685 11471 13719
rect 11471 13685 11480 13719
rect 13544 13744 13596 13796
rect 15384 13812 15436 13864
rect 15936 13812 15988 13864
rect 16396 13812 16448 13864
rect 17224 13812 17276 13864
rect 18696 13812 18748 13864
rect 19984 13744 20036 13796
rect 21180 13812 21232 13864
rect 23112 13812 23164 13864
rect 23940 13855 23992 13864
rect 23940 13821 23949 13855
rect 23949 13821 23983 13855
rect 23983 13821 23992 13855
rect 23940 13812 23992 13821
rect 11428 13676 11480 13685
rect 15384 13676 15436 13728
rect 20904 13676 20956 13728
rect 22560 13676 22612 13728
rect 25596 13719 25648 13728
rect 25596 13685 25605 13719
rect 25605 13685 25639 13719
rect 25639 13685 25648 13719
rect 25596 13676 25648 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2780 13472 2832 13524
rect 4160 13472 4212 13524
rect 5264 13472 5316 13524
rect 5540 13472 5592 13524
rect 6644 13515 6696 13524
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 9588 13472 9640 13524
rect 16856 13472 16908 13524
rect 17316 13515 17368 13524
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 18696 13472 18748 13524
rect 18880 13472 18932 13524
rect 2044 13404 2096 13456
rect 5448 13404 5500 13456
rect 6276 13404 6328 13456
rect 3884 13336 3936 13388
rect 4712 13336 4764 13388
rect 8300 13404 8352 13456
rect 9680 13404 9732 13456
rect 10048 13404 10100 13456
rect 10232 13447 10284 13456
rect 10232 13413 10241 13447
rect 10241 13413 10275 13447
rect 10275 13413 10284 13447
rect 10232 13404 10284 13413
rect 10692 13404 10744 13456
rect 10876 13404 10928 13456
rect 13820 13447 13872 13456
rect 13820 13413 13829 13447
rect 13829 13413 13863 13447
rect 13863 13413 13872 13447
rect 13820 13404 13872 13413
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 12532 13379 12584 13388
rect 12532 13345 12541 13379
rect 12541 13345 12575 13379
rect 12575 13345 12584 13379
rect 12532 13336 12584 13345
rect 2688 13268 2740 13320
rect 5540 13268 5592 13320
rect 11060 13268 11112 13320
rect 13268 13268 13320 13320
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 13912 13268 13964 13320
rect 4620 13200 4672 13252
rect 15476 13404 15528 13456
rect 16764 13404 16816 13456
rect 17684 13447 17736 13456
rect 17684 13413 17693 13447
rect 17693 13413 17727 13447
rect 17727 13413 17736 13447
rect 17684 13404 17736 13413
rect 19156 13379 19208 13388
rect 19156 13345 19174 13379
rect 19174 13345 19208 13379
rect 19156 13336 19208 13345
rect 20996 13379 21048 13388
rect 20996 13345 21014 13379
rect 21014 13345 21048 13379
rect 20996 13336 21048 13345
rect 23388 13336 23440 13388
rect 23572 13379 23624 13388
rect 23572 13345 23616 13379
rect 23616 13345 23624 13379
rect 23572 13336 23624 13345
rect 24032 13336 24084 13388
rect 25136 13336 25188 13388
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 17316 13268 17368 13320
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 23480 13200 23532 13252
rect 1860 13132 1912 13184
rect 2228 13132 2280 13184
rect 4988 13132 5040 13184
rect 5448 13132 5500 13184
rect 6828 13132 6880 13184
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 9772 13132 9824 13184
rect 11060 13132 11112 13184
rect 15384 13132 15436 13184
rect 21088 13132 21140 13184
rect 22836 13132 22888 13184
rect 24216 13132 24268 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2780 12928 2832 12980
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 2688 12724 2740 12776
rect 4712 12928 4764 12980
rect 6276 12928 6328 12980
rect 8300 12928 8352 12980
rect 10140 12928 10192 12980
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 13544 12928 13596 12980
rect 13820 12928 13872 12980
rect 16028 12928 16080 12980
rect 16764 12971 16816 12980
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 17500 12928 17552 12980
rect 17684 12928 17736 12980
rect 4068 12903 4120 12912
rect 4068 12869 4077 12903
rect 4077 12869 4111 12903
rect 4111 12869 4120 12903
rect 4068 12860 4120 12869
rect 10876 12903 10928 12912
rect 10876 12869 10885 12903
rect 10885 12869 10919 12903
rect 10919 12869 10928 12903
rect 10876 12860 10928 12869
rect 18052 12860 18104 12912
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 5264 12792 5316 12844
rect 7104 12792 7156 12844
rect 7748 12792 7800 12844
rect 8024 12792 8076 12844
rect 12348 12792 12400 12844
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 16028 12792 16080 12844
rect 16304 12835 16356 12844
rect 16304 12801 16313 12835
rect 16313 12801 16347 12835
rect 16347 12801 16356 12835
rect 16304 12792 16356 12801
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 7656 12724 7708 12776
rect 8760 12767 8812 12776
rect 8760 12733 8804 12767
rect 8804 12733 8812 12767
rect 8760 12724 8812 12733
rect 11152 12724 11204 12776
rect 12440 12724 12492 12776
rect 5724 12699 5776 12708
rect 2044 12588 2096 12640
rect 4804 12588 4856 12640
rect 5724 12665 5733 12699
rect 5733 12665 5767 12699
rect 5767 12665 5776 12699
rect 5724 12656 5776 12665
rect 7104 12588 7156 12640
rect 8576 12631 8628 12640
rect 8576 12597 8585 12631
rect 8585 12597 8619 12631
rect 8619 12597 8628 12631
rect 8576 12588 8628 12597
rect 10692 12656 10744 12708
rect 11060 12588 11112 12640
rect 12348 12656 12400 12708
rect 13636 12656 13688 12708
rect 17592 12724 17644 12776
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 14280 12699 14332 12708
rect 14280 12665 14289 12699
rect 14289 12665 14323 12699
rect 14323 12665 14332 12699
rect 14280 12656 14332 12665
rect 14372 12699 14424 12708
rect 14372 12665 14381 12699
rect 14381 12665 14415 12699
rect 14415 12665 14424 12699
rect 14372 12656 14424 12665
rect 12532 12588 12584 12640
rect 12716 12588 12768 12640
rect 15292 12588 15344 12640
rect 18052 12588 18104 12640
rect 18696 12724 18748 12776
rect 20628 12928 20680 12980
rect 20996 12928 21048 12980
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 23572 12928 23624 12980
rect 24216 12928 24268 12980
rect 25136 12971 25188 12980
rect 20812 12767 20864 12776
rect 20812 12733 20856 12767
rect 20856 12733 20864 12767
rect 20812 12724 20864 12733
rect 22652 12767 22704 12776
rect 22652 12733 22670 12767
rect 22670 12733 22704 12767
rect 25136 12937 25145 12971
rect 25145 12937 25179 12971
rect 25179 12937 25188 12971
rect 25136 12928 25188 12937
rect 22652 12724 22704 12733
rect 25044 12656 25096 12708
rect 18420 12588 18472 12640
rect 18696 12588 18748 12640
rect 19156 12631 19208 12640
rect 19156 12597 19165 12631
rect 19165 12597 19199 12631
rect 19199 12597 19208 12631
rect 19156 12588 19208 12597
rect 19340 12588 19392 12640
rect 20996 12588 21048 12640
rect 23388 12588 23440 12640
rect 25136 12588 25188 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2780 12384 2832 12436
rect 3516 12427 3568 12436
rect 3516 12393 3525 12427
rect 3525 12393 3559 12427
rect 3559 12393 3568 12427
rect 3516 12384 3568 12393
rect 4988 12384 5040 12436
rect 5356 12384 5408 12436
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 7840 12384 7892 12436
rect 9496 12427 9548 12436
rect 9496 12393 9505 12427
rect 9505 12393 9539 12427
rect 9539 12393 9548 12427
rect 9496 12384 9548 12393
rect 9772 12384 9824 12436
rect 9864 12384 9916 12436
rect 1584 12316 1636 12368
rect 2320 12316 2372 12368
rect 4160 12316 4212 12368
rect 6092 12291 6144 12300
rect 2964 12180 3016 12232
rect 3976 12180 4028 12232
rect 4252 12180 4304 12232
rect 5448 12180 5500 12232
rect 5724 12180 5776 12232
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 7656 12316 7708 12368
rect 6092 12248 6144 12257
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 6000 12180 6052 12232
rect 7656 12180 7708 12232
rect 11060 12384 11112 12436
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 14280 12384 14332 12436
rect 18144 12384 18196 12436
rect 22284 12384 22336 12436
rect 22468 12384 22520 12436
rect 8484 12248 8536 12300
rect 9128 12248 9180 12300
rect 10784 12316 10836 12368
rect 12532 12316 12584 12368
rect 14372 12316 14424 12368
rect 16212 12359 16264 12368
rect 16212 12325 16221 12359
rect 16221 12325 16255 12359
rect 16255 12325 16264 12359
rect 16212 12316 16264 12325
rect 17776 12359 17828 12368
rect 17776 12325 17785 12359
rect 17785 12325 17819 12359
rect 17819 12325 17828 12359
rect 17776 12316 17828 12325
rect 18420 12316 18472 12368
rect 11428 12248 11480 12300
rect 12164 12248 12216 12300
rect 14280 12248 14332 12300
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 20812 12248 20864 12300
rect 22284 12291 22336 12300
rect 22284 12257 22302 12291
rect 22302 12257 22336 12291
rect 22284 12248 22336 12257
rect 24124 12248 24176 12300
rect 24768 12291 24820 12300
rect 24768 12257 24786 12291
rect 24786 12257 24820 12291
rect 24768 12248 24820 12257
rect 7932 12180 7984 12232
rect 9312 12180 9364 12232
rect 1400 12112 1452 12164
rect 8668 12112 8720 12164
rect 10140 12180 10192 12232
rect 10600 12112 10652 12164
rect 1860 12044 1912 12096
rect 2136 12044 2188 12096
rect 10692 12044 10744 12096
rect 16304 12180 16356 12232
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 16764 12180 16816 12189
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 14832 12112 14884 12164
rect 22100 12112 22152 12164
rect 16028 12044 16080 12096
rect 18144 12044 18196 12096
rect 19432 12087 19484 12096
rect 19432 12053 19441 12087
rect 19441 12053 19475 12087
rect 19475 12053 19484 12087
rect 19432 12044 19484 12053
rect 20720 12044 20772 12096
rect 22928 12044 22980 12096
rect 24952 12044 25004 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 2320 11840 2372 11892
rect 2780 11840 2832 11892
rect 6092 11840 6144 11892
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 6920 11840 6972 11892
rect 7380 11840 7432 11892
rect 10600 11883 10652 11892
rect 10600 11849 10609 11883
rect 10609 11849 10643 11883
rect 10643 11849 10652 11883
rect 10600 11840 10652 11849
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 17684 11840 17736 11892
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 24768 11840 24820 11892
rect 1308 11704 1360 11756
rect 1584 11704 1636 11756
rect 1676 11704 1728 11756
rect 3516 11772 3568 11824
rect 3700 11772 3752 11824
rect 6000 11772 6052 11824
rect 6736 11772 6788 11824
rect 8484 11772 8536 11824
rect 10324 11815 10376 11824
rect 10324 11781 10333 11815
rect 10333 11781 10367 11815
rect 10367 11781 10376 11815
rect 10324 11772 10376 11781
rect 12348 11772 12400 11824
rect 2412 11704 2464 11756
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 7288 11704 7340 11756
rect 9496 11704 9548 11756
rect 12624 11704 12676 11756
rect 14648 11704 14700 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 18144 11704 18196 11713
rect 18236 11704 18288 11756
rect 7840 11636 7892 11688
rect 14280 11679 14332 11688
rect 2228 11568 2280 11620
rect 2964 11568 3016 11620
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 5816 11568 5868 11620
rect 3608 11500 3660 11509
rect 4160 11500 4212 11552
rect 6368 11500 6420 11552
rect 6552 11568 6604 11620
rect 6920 11568 6972 11620
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 9588 11568 9640 11620
rect 9036 11500 9088 11552
rect 9496 11500 9548 11552
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 14832 11636 14884 11688
rect 16764 11679 16816 11688
rect 16764 11645 16773 11679
rect 16773 11645 16807 11679
rect 16807 11645 16816 11679
rect 16764 11636 16816 11645
rect 21272 11679 21324 11688
rect 21272 11645 21281 11679
rect 21281 11645 21315 11679
rect 21315 11645 21324 11679
rect 21272 11636 21324 11645
rect 23480 11636 23532 11688
rect 23940 11704 23992 11756
rect 15384 11568 15436 11620
rect 15844 11568 15896 11620
rect 17132 11568 17184 11620
rect 19432 11568 19484 11620
rect 20352 11611 20404 11620
rect 20352 11577 20361 11611
rect 20361 11577 20395 11611
rect 20395 11577 20404 11611
rect 20352 11568 20404 11577
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 13268 11500 13320 11552
rect 16212 11500 16264 11552
rect 16396 11500 16448 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 20812 11500 20864 11552
rect 21640 11543 21692 11552
rect 21640 11509 21649 11543
rect 21649 11509 21683 11543
rect 21683 11509 21692 11543
rect 21640 11500 21692 11509
rect 23664 11500 23716 11552
rect 24124 11679 24176 11688
rect 24124 11645 24133 11679
rect 24133 11645 24167 11679
rect 24167 11645 24176 11679
rect 24124 11636 24176 11645
rect 24308 11636 24360 11688
rect 24124 11500 24176 11552
rect 24400 11500 24452 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1952 11296 2004 11348
rect 2228 11339 2280 11348
rect 2228 11305 2237 11339
rect 2237 11305 2271 11339
rect 2271 11305 2280 11339
rect 2228 11296 2280 11305
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 5816 11296 5868 11348
rect 7288 11296 7340 11348
rect 9496 11339 9548 11348
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 15016 11339 15068 11348
rect 15016 11305 15025 11339
rect 15025 11305 15059 11339
rect 15059 11305 15068 11339
rect 15016 11296 15068 11305
rect 16304 11339 16356 11348
rect 16304 11305 16313 11339
rect 16313 11305 16347 11339
rect 16347 11305 16356 11339
rect 16304 11296 16356 11305
rect 18420 11339 18472 11348
rect 2504 11271 2556 11280
rect 2504 11237 2513 11271
rect 2513 11237 2547 11271
rect 2547 11237 2556 11271
rect 2504 11228 2556 11237
rect 3148 11228 3200 11280
rect 3608 11228 3660 11280
rect 4160 11228 4212 11280
rect 4804 11271 4856 11280
rect 4804 11237 4813 11271
rect 4813 11237 4847 11271
rect 4847 11237 4856 11271
rect 4804 11228 4856 11237
rect 5356 11271 5408 11280
rect 5356 11237 5365 11271
rect 5365 11237 5399 11271
rect 5399 11237 5408 11271
rect 5356 11228 5408 11237
rect 6552 11271 6604 11280
rect 6552 11237 6555 11271
rect 6555 11237 6589 11271
rect 6589 11237 6604 11271
rect 6552 11228 6604 11237
rect 8116 11228 8168 11280
rect 8392 11228 8444 11280
rect 12256 11228 12308 11280
rect 12624 11228 12676 11280
rect 13268 11228 13320 11280
rect 14372 11271 14424 11280
rect 14372 11237 14381 11271
rect 14381 11237 14415 11271
rect 14415 11237 14424 11271
rect 14372 11228 14424 11237
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 17408 11228 17460 11280
rect 18420 11305 18429 11339
rect 18429 11305 18463 11339
rect 18463 11305 18472 11339
rect 18420 11296 18472 11305
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 19248 11228 19300 11280
rect 20352 11228 20404 11280
rect 21640 11228 21692 11280
rect 1676 11160 1728 11212
rect 6920 11160 6972 11212
rect 9404 11160 9456 11212
rect 11796 11160 11848 11212
rect 4160 11092 4212 11144
rect 4896 11092 4948 11144
rect 2964 11024 3016 11076
rect 8208 11092 8260 11144
rect 9772 11092 9824 11144
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 4252 10956 4304 11008
rect 7288 11024 7340 11076
rect 8484 11024 8536 11076
rect 16580 11092 16632 11144
rect 18236 11092 18288 11144
rect 22100 11092 22152 11144
rect 6920 10956 6972 11008
rect 11060 10956 11112 11008
rect 13820 10956 13872 11008
rect 24216 11160 24268 11212
rect 24676 11160 24728 11212
rect 23940 11092 23992 11144
rect 24400 11092 24452 11144
rect 21824 10956 21876 11008
rect 23020 10956 23072 11008
rect 24860 11024 24912 11076
rect 24768 10999 24820 11008
rect 24768 10965 24777 10999
rect 24777 10965 24811 10999
rect 24811 10965 24820 10999
rect 24768 10956 24820 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 3148 10752 3200 10804
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 9496 10752 9548 10804
rect 10692 10752 10744 10804
rect 11796 10752 11848 10804
rect 13268 10795 13320 10804
rect 13268 10761 13277 10795
rect 13277 10761 13311 10795
rect 13311 10761 13320 10795
rect 13268 10752 13320 10761
rect 15476 10752 15528 10804
rect 15844 10752 15896 10804
rect 17132 10795 17184 10804
rect 2504 10684 2556 10736
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 2044 10480 2096 10489
rect 2504 10480 2556 10532
rect 5172 10684 5224 10736
rect 7748 10684 7800 10736
rect 9772 10684 9824 10736
rect 5356 10616 5408 10668
rect 6000 10616 6052 10668
rect 6184 10616 6236 10668
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 7104 10548 7156 10557
rect 8208 10616 8260 10668
rect 9680 10616 9732 10668
rect 10140 10616 10192 10668
rect 13820 10616 13872 10668
rect 15384 10616 15436 10668
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 20996 10795 21048 10804
rect 20996 10761 21005 10795
rect 21005 10761 21039 10795
rect 21039 10761 21048 10795
rect 20996 10752 21048 10761
rect 21272 10684 21324 10736
rect 7840 10548 7892 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 7656 10480 7708 10532
rect 3608 10412 3660 10464
rect 3792 10412 3844 10464
rect 5172 10412 5224 10464
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 6552 10412 6604 10464
rect 6920 10455 6972 10464
rect 6920 10421 6929 10455
rect 6929 10421 6963 10455
rect 6963 10421 6972 10455
rect 6920 10412 6972 10421
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 7840 10412 7892 10421
rect 8300 10412 8352 10464
rect 13912 10523 13964 10532
rect 13912 10489 13921 10523
rect 13921 10489 13955 10523
rect 13955 10489 13964 10523
rect 13912 10480 13964 10489
rect 15108 10480 15160 10532
rect 17408 10523 17460 10532
rect 17408 10489 17417 10523
rect 17417 10489 17451 10523
rect 17451 10489 17460 10523
rect 17408 10480 17460 10489
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 12256 10412 12308 10464
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 16948 10412 17000 10464
rect 21640 10752 21692 10804
rect 22100 10752 22152 10804
rect 23020 10795 23072 10804
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 21824 10616 21876 10668
rect 24676 10616 24728 10668
rect 25136 10616 25188 10668
rect 18328 10591 18380 10600
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 18236 10480 18288 10532
rect 23848 10548 23900 10600
rect 24860 10548 24912 10600
rect 18512 10455 18564 10464
rect 18512 10421 18521 10455
rect 18521 10421 18555 10455
rect 18555 10421 18564 10455
rect 18512 10412 18564 10421
rect 19524 10412 19576 10464
rect 20352 10412 20404 10464
rect 21272 10412 21324 10464
rect 25044 10480 25096 10532
rect 23112 10412 23164 10464
rect 23480 10412 23532 10464
rect 25412 10455 25464 10464
rect 25412 10421 25421 10455
rect 25421 10421 25455 10455
rect 25455 10421 25464 10455
rect 25412 10412 25464 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2780 10208 2832 10260
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 4068 10208 4120 10260
rect 5448 10208 5500 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8392 10208 8444 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 10140 10208 10192 10260
rect 11520 10251 11572 10260
rect 11520 10217 11529 10251
rect 11529 10217 11563 10251
rect 11563 10217 11572 10251
rect 13360 10251 13412 10260
rect 11520 10208 11572 10217
rect 2504 10140 2556 10192
rect 3976 10140 4028 10192
rect 6000 10140 6052 10192
rect 6184 10183 6236 10192
rect 6184 10149 6187 10183
rect 6187 10149 6221 10183
rect 6221 10149 6236 10183
rect 6184 10140 6236 10149
rect 5356 10072 5408 10124
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 10416 10140 10468 10192
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13820 10208 13872 10260
rect 15384 10251 15436 10260
rect 15384 10217 15393 10251
rect 15393 10217 15427 10251
rect 15427 10217 15436 10251
rect 15384 10208 15436 10217
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 18604 10208 18656 10260
rect 21272 10208 21324 10260
rect 21640 10208 21692 10260
rect 22560 10208 22612 10260
rect 23388 10208 23440 10260
rect 23756 10208 23808 10260
rect 8208 10072 8260 10124
rect 12072 10072 12124 10124
rect 19892 10140 19944 10192
rect 20168 10140 20220 10192
rect 20536 10140 20588 10192
rect 21916 10183 21968 10192
rect 21916 10149 21925 10183
rect 21925 10149 21959 10183
rect 21959 10149 21968 10183
rect 21916 10140 21968 10149
rect 23480 10183 23532 10192
rect 23480 10149 23489 10183
rect 23489 10149 23523 10183
rect 23523 10149 23532 10183
rect 23480 10140 23532 10149
rect 24952 10183 25004 10192
rect 24952 10149 24961 10183
rect 24961 10149 24995 10183
rect 24995 10149 25004 10183
rect 24952 10140 25004 10149
rect 25044 10183 25096 10192
rect 25044 10149 25053 10183
rect 25053 10149 25087 10183
rect 25087 10149 25096 10183
rect 25044 10140 25096 10149
rect 13176 10072 13228 10124
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 14096 10072 14148 10124
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 15568 10072 15620 10124
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 19984 10115 20036 10124
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 4252 10004 4304 10056
rect 6184 10004 6236 10056
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 10876 10004 10928 10056
rect 13452 10004 13504 10056
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 20168 10004 20220 10056
rect 20536 10004 20588 10056
rect 21364 10004 21416 10056
rect 21824 10047 21876 10056
rect 21824 10013 21833 10047
rect 21833 10013 21867 10047
rect 21867 10013 21876 10047
rect 21824 10004 21876 10013
rect 23388 10047 23440 10056
rect 23388 10013 23397 10047
rect 23397 10013 23431 10047
rect 23431 10013 23440 10047
rect 23388 10004 23440 10013
rect 10324 9979 10376 9988
rect 10324 9945 10333 9979
rect 10333 9945 10367 9979
rect 10367 9945 10376 9979
rect 10324 9936 10376 9945
rect 10692 9936 10744 9988
rect 11336 9936 11388 9988
rect 12992 9979 13044 9988
rect 12992 9945 13001 9979
rect 13001 9945 13035 9979
rect 13035 9945 13044 9979
rect 12992 9936 13044 9945
rect 18236 9936 18288 9988
rect 18972 9936 19024 9988
rect 23296 9936 23348 9988
rect 25136 10004 25188 10056
rect 3608 9868 3660 9920
rect 4160 9868 4212 9920
rect 12164 9911 12216 9920
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 12164 9868 12216 9877
rect 13820 9868 13872 9920
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 16396 9868 16448 9877
rect 17224 9868 17276 9920
rect 17684 9868 17736 9920
rect 18328 9868 18380 9920
rect 20444 9911 20496 9920
rect 20444 9877 20453 9911
rect 20453 9877 20487 9911
rect 20487 9877 20496 9911
rect 20444 9868 20496 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 7288 9664 7340 9716
rect 7748 9664 7800 9716
rect 8116 9664 8168 9716
rect 14096 9664 14148 9716
rect 15292 9707 15344 9716
rect 15292 9673 15301 9707
rect 15301 9673 15335 9707
rect 15335 9673 15344 9707
rect 15292 9664 15344 9673
rect 18328 9664 18380 9716
rect 18696 9664 18748 9716
rect 21824 9664 21876 9716
rect 3976 9596 4028 9648
rect 3516 9528 3568 9580
rect 4712 9596 4764 9648
rect 6828 9596 6880 9648
rect 7104 9596 7156 9648
rect 5448 9528 5500 9580
rect 6000 9528 6052 9580
rect 7012 9528 7064 9580
rect 2504 9435 2556 9444
rect 2504 9401 2507 9435
rect 2507 9401 2541 9435
rect 2541 9401 2556 9435
rect 2504 9392 2556 9401
rect 7288 9460 7340 9512
rect 9220 9639 9272 9648
rect 9220 9605 9229 9639
rect 9229 9605 9263 9639
rect 9263 9605 9272 9639
rect 9220 9596 9272 9605
rect 10324 9639 10376 9648
rect 10324 9605 10333 9639
rect 10333 9605 10367 9639
rect 10367 9605 10376 9639
rect 10324 9596 10376 9605
rect 10876 9596 10928 9648
rect 11796 9639 11848 9648
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 12992 9596 13044 9648
rect 16396 9596 16448 9648
rect 10416 9460 10468 9512
rect 11060 9460 11112 9512
rect 13360 9528 13412 9580
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 14832 9528 14884 9580
rect 16856 9528 16908 9580
rect 19248 9596 19300 9648
rect 19340 9596 19392 9648
rect 19524 9639 19576 9648
rect 19524 9605 19533 9639
rect 19533 9605 19567 9639
rect 19567 9605 19576 9639
rect 19524 9596 19576 9605
rect 20168 9596 20220 9648
rect 21916 9596 21968 9648
rect 18420 9528 18472 9580
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 20812 9528 20864 9580
rect 23296 9664 23348 9716
rect 23204 9596 23256 9648
rect 23480 9664 23532 9716
rect 24124 9664 24176 9716
rect 25044 9664 25096 9716
rect 14464 9503 14516 9512
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 8300 9392 8352 9444
rect 5816 9324 5868 9376
rect 6000 9324 6052 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 9588 9392 9640 9444
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 10876 9392 10928 9444
rect 12164 9392 12216 9444
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 15292 9460 15344 9512
rect 15844 9503 15896 9512
rect 14372 9392 14424 9444
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 17132 9460 17184 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18604 9503 18656 9512
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 18144 9392 18196 9444
rect 19248 9460 19300 9512
rect 19432 9460 19484 9512
rect 20444 9503 20496 9512
rect 20444 9469 20453 9503
rect 20453 9469 20487 9503
rect 20487 9469 20496 9503
rect 20444 9460 20496 9469
rect 20812 9435 20864 9444
rect 20812 9401 20815 9435
rect 20815 9401 20849 9435
rect 20849 9401 20864 9435
rect 20812 9392 20864 9401
rect 23204 9460 23256 9512
rect 24308 9596 24360 9648
rect 23756 9571 23808 9580
rect 23756 9537 23765 9571
rect 23765 9537 23799 9571
rect 23799 9537 23808 9571
rect 23756 9528 23808 9537
rect 24124 9528 24176 9580
rect 25136 9528 25188 9580
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 23848 9435 23900 9444
rect 23848 9401 23857 9435
rect 23857 9401 23891 9435
rect 23891 9401 23900 9435
rect 23848 9392 23900 9401
rect 24032 9392 24084 9444
rect 12072 9367 12124 9376
rect 9496 9324 9548 9333
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15200 9324 15252 9376
rect 15936 9324 15988 9376
rect 23296 9324 23348 9376
rect 23756 9324 23808 9376
rect 24860 9324 24912 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1952 9120 2004 9172
rect 4252 9163 4304 9172
rect 4252 9129 4261 9163
rect 4261 9129 4295 9163
rect 4295 9129 4304 9163
rect 4252 9120 4304 9129
rect 5816 9163 5868 9172
rect 5816 9129 5825 9163
rect 5825 9129 5859 9163
rect 5859 9129 5868 9163
rect 5816 9120 5868 9129
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 6920 9120 6972 9172
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 9772 9120 9824 9172
rect 12532 9120 12584 9172
rect 13728 9120 13780 9172
rect 14188 9120 14240 9172
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 19340 9120 19392 9172
rect 20168 9163 20220 9172
rect 20168 9129 20177 9163
rect 20177 9129 20211 9163
rect 20211 9129 20220 9163
rect 20168 9120 20220 9129
rect 21364 9163 21416 9172
rect 21364 9129 21373 9163
rect 21373 9129 21407 9163
rect 21407 9129 21416 9163
rect 21364 9120 21416 9129
rect 23204 9120 23256 9172
rect 1676 8984 1728 9036
rect 2136 9052 2188 9104
rect 4988 9052 5040 9104
rect 5172 9052 5224 9104
rect 6000 9052 6052 9104
rect 6828 9095 6880 9104
rect 6828 9061 6837 9095
rect 6837 9061 6871 9095
rect 6871 9061 6880 9095
rect 6828 9052 6880 9061
rect 2044 9027 2096 9036
rect 2044 8993 2053 9027
rect 2053 8993 2087 9027
rect 2087 8993 2096 9027
rect 2044 8984 2096 8993
rect 6184 8984 6236 9036
rect 9312 9052 9364 9104
rect 9680 9052 9732 9104
rect 12256 9052 12308 9104
rect 12716 9052 12768 9104
rect 13176 9095 13228 9104
rect 13176 9061 13185 9095
rect 13185 9061 13219 9095
rect 13219 9061 13228 9095
rect 13176 9052 13228 9061
rect 14464 9052 14516 9104
rect 15660 9052 15712 9104
rect 11980 9027 12032 9036
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 14280 8984 14332 9036
rect 16304 9052 16356 9104
rect 21732 9052 21784 9104
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 16396 9027 16448 9036
rect 16396 8993 16405 9027
rect 16405 8993 16439 9027
rect 16439 8993 16448 9027
rect 16396 8984 16448 8993
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 18788 9027 18840 9036
rect 18788 8993 18797 9027
rect 18797 8993 18831 9027
rect 18831 8993 18840 9027
rect 18788 8984 18840 8993
rect 18972 9027 19024 9036
rect 18972 8993 18981 9027
rect 18981 8993 19015 9027
rect 19015 8993 19024 9027
rect 18972 8984 19024 8993
rect 19340 9027 19392 9036
rect 19340 8993 19349 9027
rect 19349 8993 19383 9027
rect 19383 8993 19392 9027
rect 19340 8984 19392 8993
rect 23848 9120 23900 9172
rect 23940 9120 23992 9172
rect 24124 9095 24176 9104
rect 24124 9061 24133 9095
rect 24133 9061 24167 9095
rect 24167 9061 24176 9095
rect 24124 9052 24176 9061
rect 24952 9120 25004 9172
rect 1400 8916 1452 8968
rect 2136 8916 2188 8968
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 8208 8916 8260 8968
rect 9496 8916 9548 8968
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 10692 8916 10744 8968
rect 11152 8916 11204 8968
rect 13912 8916 13964 8968
rect 14372 8916 14424 8968
rect 15568 8916 15620 8968
rect 21916 8916 21968 8968
rect 24216 8916 24268 8968
rect 15200 8848 15252 8900
rect 572 8780 624 8832
rect 7012 8780 7064 8832
rect 9680 8780 9732 8832
rect 10692 8780 10744 8832
rect 12900 8823 12952 8832
rect 12900 8789 12909 8823
rect 12909 8789 12943 8823
rect 12943 8789 12952 8823
rect 12900 8780 12952 8789
rect 15384 8780 15436 8832
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 17868 8780 17920 8832
rect 21640 8780 21692 8832
rect 24032 8780 24084 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2780 8576 2832 8628
rect 4896 8576 4948 8628
rect 6276 8576 6328 8628
rect 7012 8619 7064 8628
rect 5724 8508 5776 8560
rect 6368 8508 6420 8560
rect 4344 8440 4396 8492
rect 5448 8440 5500 8492
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 9312 8619 9364 8628
rect 9312 8585 9321 8619
rect 9321 8585 9355 8619
rect 9355 8585 9364 8619
rect 9312 8576 9364 8585
rect 10600 8576 10652 8628
rect 10876 8576 10928 8628
rect 14280 8576 14332 8628
rect 19340 8576 19392 8628
rect 23572 8576 23624 8628
rect 25136 8576 25188 8628
rect 13820 8508 13872 8560
rect 14464 8508 14516 8560
rect 17132 8508 17184 8560
rect 18788 8508 18840 8560
rect 23940 8508 23992 8560
rect 9772 8483 9824 8492
rect 7932 8372 7984 8424
rect 6276 8347 6328 8356
rect 6276 8313 6285 8347
rect 6285 8313 6319 8347
rect 6319 8313 6328 8347
rect 6276 8304 6328 8313
rect 9404 8372 9456 8424
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 12256 8440 12308 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14004 8440 14056 8492
rect 11060 8372 11112 8424
rect 14372 8415 14424 8424
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 4988 8236 5040 8288
rect 9772 8304 9824 8356
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 14832 8372 14884 8424
rect 16856 8440 16908 8492
rect 24216 8440 24268 8492
rect 15936 8415 15988 8424
rect 15936 8381 15945 8415
rect 15945 8381 15979 8415
rect 15979 8381 15988 8415
rect 15936 8372 15988 8381
rect 16396 8415 16448 8424
rect 16396 8381 16405 8415
rect 16405 8381 16439 8415
rect 16439 8381 16448 8415
rect 16396 8372 16448 8381
rect 16580 8415 16632 8424
rect 16580 8381 16589 8415
rect 16589 8381 16623 8415
rect 16623 8381 16632 8415
rect 16580 8372 16632 8381
rect 18236 8415 18288 8424
rect 15292 8304 15344 8356
rect 12164 8236 12216 8288
rect 18236 8381 18245 8415
rect 18245 8381 18279 8415
rect 18279 8381 18288 8415
rect 18236 8372 18288 8381
rect 18788 8415 18840 8424
rect 18788 8381 18797 8415
rect 18797 8381 18831 8415
rect 18831 8381 18840 8415
rect 18788 8372 18840 8381
rect 18972 8415 19024 8424
rect 18972 8381 18981 8415
rect 18981 8381 19015 8415
rect 19015 8381 19024 8415
rect 18972 8372 19024 8381
rect 19524 8415 19576 8424
rect 19524 8381 19533 8415
rect 19533 8381 19567 8415
rect 19567 8381 19576 8415
rect 19524 8372 19576 8381
rect 19984 8372 20036 8424
rect 16488 8236 16540 8288
rect 17868 8304 17920 8356
rect 20260 8347 20312 8356
rect 20260 8313 20269 8347
rect 20269 8313 20303 8347
rect 20303 8313 20312 8347
rect 23940 8372 23992 8424
rect 20260 8304 20312 8313
rect 21732 8304 21784 8356
rect 23572 8304 23624 8356
rect 18052 8236 18104 8288
rect 20812 8236 20864 8288
rect 24032 8279 24084 8288
rect 24032 8245 24041 8279
rect 24041 8245 24075 8279
rect 24075 8245 24084 8279
rect 24032 8236 24084 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 8032 1452 8084
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 4160 8075 4212 8084
rect 4160 8041 4169 8075
rect 4169 8041 4203 8075
rect 4203 8041 4212 8075
rect 4160 8032 4212 8041
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 7288 8075 7340 8084
rect 7288 8041 7297 8075
rect 7297 8041 7331 8075
rect 7331 8041 7340 8075
rect 7288 8032 7340 8041
rect 9496 8075 9548 8084
rect 9496 8041 9505 8075
rect 9505 8041 9539 8075
rect 9539 8041 9548 8075
rect 9496 8032 9548 8041
rect 9680 8032 9732 8084
rect 11980 8075 12032 8084
rect 11980 8041 11989 8075
rect 11989 8041 12023 8075
rect 12023 8041 12032 8075
rect 11980 8032 12032 8041
rect 12348 8032 12400 8084
rect 12532 8032 12584 8084
rect 13636 8032 13688 8084
rect 14096 8032 14148 8084
rect 16396 8075 16448 8084
rect 16396 8041 16405 8075
rect 16405 8041 16439 8075
rect 16439 8041 16448 8075
rect 16396 8032 16448 8041
rect 17132 8032 17184 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 21916 8075 21968 8084
rect 21916 8041 21925 8075
rect 21925 8041 21959 8075
rect 21959 8041 21968 8075
rect 21916 8032 21968 8041
rect 2320 7964 2372 8016
rect 2504 7964 2556 8016
rect 6828 7964 6880 8016
rect 7104 7964 7156 8016
rect 2228 7939 2280 7948
rect 2228 7905 2237 7939
rect 2237 7905 2271 7939
rect 2271 7905 2280 7939
rect 2228 7896 2280 7905
rect 4160 7939 4212 7948
rect 4160 7905 4169 7939
rect 4169 7905 4203 7939
rect 4203 7905 4212 7939
rect 4160 7896 4212 7905
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 6000 7896 6052 7948
rect 6184 7939 6236 7948
rect 6184 7905 6193 7939
rect 6193 7905 6227 7939
rect 6227 7905 6236 7939
rect 6184 7896 6236 7905
rect 10232 7964 10284 8016
rect 12716 7964 12768 8016
rect 12900 7964 12952 8016
rect 13176 7964 13228 8016
rect 14372 7964 14424 8016
rect 8852 7896 8904 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 14464 7896 14516 7948
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 16580 7964 16632 8016
rect 20996 7964 21048 8016
rect 22560 7964 22612 8016
rect 24032 8007 24084 8016
rect 24032 7973 24041 8007
rect 24041 7973 24075 8007
rect 24075 7973 24084 8007
rect 24032 7964 24084 7973
rect 15936 7896 15988 7948
rect 16764 7896 16816 7948
rect 16948 7896 17000 7948
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 18604 7896 18656 7948
rect 19524 7939 19576 7948
rect 2044 7828 2096 7837
rect 8116 7828 8168 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 12348 7828 12400 7880
rect 12992 7828 13044 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 18144 7828 18196 7880
rect 19524 7905 19533 7939
rect 19533 7905 19567 7939
rect 19567 7905 19576 7939
rect 19524 7896 19576 7905
rect 22100 7896 22152 7948
rect 21088 7828 21140 7880
rect 23940 7896 23992 7948
rect 23296 7828 23348 7880
rect 2412 7760 2464 7812
rect 6828 7803 6880 7812
rect 6828 7769 6837 7803
rect 6837 7769 6871 7803
rect 6871 7769 6880 7803
rect 6828 7760 6880 7769
rect 12164 7760 12216 7812
rect 15660 7760 15712 7812
rect 16856 7760 16908 7812
rect 22008 7760 22060 7812
rect 23204 7760 23256 7812
rect 24032 7760 24084 7812
rect 3056 7692 3108 7744
rect 4804 7692 4856 7744
rect 5540 7692 5592 7744
rect 7932 7692 7984 7744
rect 9772 7692 9824 7744
rect 10416 7692 10468 7744
rect 10692 7692 10744 7744
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 15844 7692 15896 7744
rect 17868 7692 17920 7744
rect 20168 7735 20220 7744
rect 20168 7701 20177 7735
rect 20177 7701 20211 7735
rect 20211 7701 20220 7735
rect 20168 7692 20220 7701
rect 23756 7692 23808 7744
rect 24124 7692 24176 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2320 7488 2372 7540
rect 4988 7488 5040 7540
rect 6000 7488 6052 7540
rect 6736 7488 6788 7540
rect 8116 7488 8168 7540
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8300 7488 8352 7497
rect 9404 7488 9456 7540
rect 10232 7488 10284 7540
rect 11428 7531 11480 7540
rect 11428 7497 11437 7531
rect 11437 7497 11471 7531
rect 11471 7497 11480 7531
rect 11428 7488 11480 7497
rect 12256 7488 12308 7540
rect 12440 7488 12492 7540
rect 2688 7420 2740 7472
rect 4160 7420 4212 7472
rect 10876 7463 10928 7472
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 4068 7352 4120 7404
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 10876 7429 10885 7463
rect 10885 7429 10919 7463
rect 10919 7429 10928 7463
rect 10876 7420 10928 7429
rect 12808 7488 12860 7540
rect 13268 7488 13320 7540
rect 13636 7488 13688 7540
rect 15936 7488 15988 7540
rect 18052 7488 18104 7540
rect 19524 7488 19576 7540
rect 23940 7488 23992 7540
rect 14096 7463 14148 7472
rect 14096 7429 14105 7463
rect 14105 7429 14139 7463
rect 14139 7429 14148 7463
rect 14096 7420 14148 7429
rect 7748 7352 7800 7404
rect 10140 7352 10192 7404
rect 14832 7420 14884 7472
rect 20996 7420 21048 7472
rect 22008 7420 22060 7472
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 15292 7352 15344 7404
rect 17868 7352 17920 7404
rect 22100 7352 22152 7404
rect 23480 7352 23532 7404
rect 23756 7395 23808 7404
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 23756 7352 23808 7361
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 7104 7284 7156 7336
rect 8300 7284 8352 7336
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 12532 7284 12584 7336
rect 14004 7327 14056 7336
rect 2964 7259 3016 7268
rect 2964 7225 2973 7259
rect 2973 7225 3007 7259
rect 3007 7225 3016 7259
rect 2964 7216 3016 7225
rect 3056 7259 3108 7268
rect 3056 7225 3065 7259
rect 3065 7225 3099 7259
rect 3099 7225 3108 7259
rect 3056 7216 3108 7225
rect 4988 7216 5040 7268
rect 5356 7216 5408 7268
rect 10416 7259 10468 7268
rect 10416 7225 10425 7259
rect 10425 7225 10459 7259
rect 10459 7225 10468 7259
rect 10416 7216 10468 7225
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 16580 7327 16632 7336
rect 16580 7293 16589 7327
rect 16589 7293 16623 7327
rect 16623 7293 16632 7327
rect 16580 7284 16632 7293
rect 19156 7327 19208 7336
rect 19156 7293 19165 7327
rect 19165 7293 19199 7327
rect 19199 7293 19208 7327
rect 19156 7284 19208 7293
rect 19432 7284 19484 7336
rect 20168 7327 20220 7336
rect 20168 7293 20177 7327
rect 20177 7293 20211 7327
rect 20211 7293 20220 7327
rect 20168 7284 20220 7293
rect 25228 7327 25280 7336
rect 25228 7293 25237 7327
rect 25237 7293 25271 7327
rect 25271 7293 25280 7327
rect 25228 7284 25280 7293
rect 17132 7259 17184 7268
rect 2044 7148 2096 7200
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 17132 7225 17141 7259
rect 17141 7225 17175 7259
rect 17175 7225 17184 7259
rect 17132 7216 17184 7225
rect 20812 7216 20864 7268
rect 20904 7216 20956 7268
rect 21548 7216 21600 7268
rect 22008 7259 22060 7268
rect 22008 7225 22017 7259
rect 22017 7225 22051 7259
rect 22051 7225 22060 7259
rect 22008 7216 22060 7225
rect 22100 7259 22152 7268
rect 22100 7225 22109 7259
rect 22109 7225 22143 7259
rect 22143 7225 22152 7259
rect 23480 7259 23532 7268
rect 22100 7216 22152 7225
rect 23480 7225 23489 7259
rect 23489 7225 23523 7259
rect 23523 7225 23532 7259
rect 23480 7216 23532 7225
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 5540 7148 5592 7200
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 12256 7191 12308 7200
rect 12256 7157 12265 7191
rect 12265 7157 12299 7191
rect 12299 7157 12308 7191
rect 12256 7148 12308 7157
rect 12440 7148 12492 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14464 7148 14516 7200
rect 15200 7148 15252 7200
rect 16764 7148 16816 7200
rect 18144 7148 18196 7200
rect 18604 7148 18656 7200
rect 20260 7148 20312 7200
rect 20996 7148 21048 7200
rect 22560 7148 22612 7200
rect 25412 7191 25464 7200
rect 25412 7157 25421 7191
rect 25421 7157 25455 7191
rect 25455 7157 25464 7191
rect 25412 7148 25464 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2228 6944 2280 6996
rect 2320 6919 2372 6928
rect 2320 6885 2329 6919
rect 2329 6885 2363 6919
rect 2363 6885 2372 6919
rect 2320 6876 2372 6885
rect 4160 6876 4212 6928
rect 4896 6944 4948 6996
rect 6184 6944 6236 6996
rect 6828 6944 6880 6996
rect 7104 6944 7156 6996
rect 9772 6987 9824 6996
rect 9772 6953 9781 6987
rect 9781 6953 9815 6987
rect 9815 6953 9824 6987
rect 9772 6944 9824 6953
rect 13176 6987 13228 6996
rect 13176 6953 13185 6987
rect 13185 6953 13219 6987
rect 13219 6953 13228 6987
rect 13176 6944 13228 6953
rect 14004 6987 14056 6996
rect 14004 6953 14013 6987
rect 14013 6953 14047 6987
rect 14047 6953 14056 6987
rect 14004 6944 14056 6953
rect 16948 6987 17000 6996
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 1860 6740 1912 6792
rect 2964 6740 3016 6792
rect 3516 6672 3568 6724
rect 4344 6740 4396 6792
rect 5356 6740 5408 6792
rect 7380 6808 7432 6860
rect 9588 6808 9640 6860
rect 10048 6808 10100 6860
rect 12164 6851 12216 6860
rect 7288 6740 7340 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 9312 6740 9364 6792
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 14188 6851 14240 6860
rect 12440 6808 12492 6817
rect 14188 6817 14197 6851
rect 14197 6817 14231 6851
rect 14231 6817 14240 6851
rect 14188 6808 14240 6817
rect 15292 6876 15344 6928
rect 16948 6953 16957 6987
rect 16957 6953 16991 6987
rect 16991 6953 17000 6987
rect 16948 6944 17000 6953
rect 18328 6944 18380 6996
rect 15844 6851 15896 6860
rect 12348 6740 12400 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 5264 6672 5316 6724
rect 12256 6715 12308 6724
rect 12256 6681 12265 6715
rect 12265 6681 12299 6715
rect 12299 6681 12308 6715
rect 12256 6672 12308 6681
rect 12532 6672 12584 6724
rect 15844 6817 15853 6851
rect 15853 6817 15887 6851
rect 15887 6817 15896 6851
rect 15844 6808 15896 6817
rect 15660 6740 15712 6792
rect 16396 6808 16448 6860
rect 16672 6808 16724 6860
rect 18236 6808 18288 6860
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 17592 6740 17644 6792
rect 18972 6808 19024 6860
rect 21088 6944 21140 6996
rect 21640 6987 21692 6996
rect 21640 6953 21649 6987
rect 21649 6953 21683 6987
rect 21683 6953 21692 6987
rect 21640 6944 21692 6953
rect 22008 6987 22060 6996
rect 22008 6953 22017 6987
rect 22017 6953 22051 6987
rect 22051 6953 22060 6987
rect 22008 6944 22060 6953
rect 23296 6987 23348 6996
rect 23296 6953 23305 6987
rect 23305 6953 23339 6987
rect 23339 6953 23348 6987
rect 23296 6944 23348 6953
rect 23756 6987 23808 6996
rect 23756 6953 23765 6987
rect 23765 6953 23799 6987
rect 23799 6953 23808 6987
rect 23756 6944 23808 6953
rect 19340 6808 19392 6860
rect 20904 6808 20956 6860
rect 22468 6919 22520 6928
rect 22468 6885 22471 6919
rect 22471 6885 22505 6919
rect 22505 6885 22520 6919
rect 22468 6876 22520 6885
rect 24216 6876 24268 6928
rect 21732 6808 21784 6860
rect 18880 6740 18932 6792
rect 24124 6740 24176 6792
rect 25044 6740 25096 6792
rect 19248 6715 19300 6724
rect 19248 6681 19257 6715
rect 19257 6681 19291 6715
rect 19291 6681 19300 6715
rect 19248 6672 19300 6681
rect 1492 6604 1544 6656
rect 1952 6604 2004 6656
rect 4712 6604 4764 6656
rect 6644 6604 6696 6656
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 12440 6604 12492 6656
rect 17408 6604 17460 6656
rect 18236 6604 18288 6656
rect 19432 6604 19484 6656
rect 21180 6647 21232 6656
rect 21180 6613 21189 6647
rect 21189 6613 21223 6647
rect 21223 6613 21232 6647
rect 21180 6604 21232 6613
rect 24216 6604 24268 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 6920 6400 6972 6452
rect 7380 6400 7432 6452
rect 10048 6443 10100 6452
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 5356 6332 5408 6384
rect 8668 6332 8720 6384
rect 10876 6375 10928 6384
rect 10876 6341 10885 6375
rect 10885 6341 10919 6375
rect 10919 6341 10928 6375
rect 10876 6332 10928 6341
rect 12164 6400 12216 6452
rect 13912 6443 13964 6452
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 7840 6264 7892 6316
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 3700 6196 3752 6248
rect 4712 6196 4764 6248
rect 2044 6128 2096 6180
rect 5264 6171 5316 6180
rect 5264 6137 5273 6171
rect 5273 6137 5307 6171
rect 5307 6137 5316 6171
rect 5264 6128 5316 6137
rect 2320 6060 2372 6112
rect 4160 6060 4212 6112
rect 5448 6128 5500 6180
rect 7104 6196 7156 6248
rect 8760 6239 8812 6248
rect 8760 6205 8769 6239
rect 8769 6205 8803 6239
rect 8803 6205 8812 6239
rect 8760 6196 8812 6205
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 6920 6103 6972 6112
rect 6920 6069 6929 6103
rect 6929 6069 6963 6103
rect 6963 6069 6972 6103
rect 6920 6060 6972 6069
rect 7288 6060 7340 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 11704 6128 11756 6180
rect 11980 6128 12032 6180
rect 12348 6196 12400 6248
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 13820 6196 13872 6248
rect 13912 6196 13964 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 16212 6332 16264 6384
rect 17592 6400 17644 6452
rect 20904 6400 20956 6452
rect 21732 6443 21784 6452
rect 21732 6409 21741 6443
rect 21741 6409 21775 6443
rect 21775 6409 21784 6443
rect 21732 6400 21784 6409
rect 23388 6400 23440 6452
rect 24124 6400 24176 6452
rect 25320 6443 25372 6452
rect 25320 6409 25329 6443
rect 25329 6409 25363 6443
rect 25363 6409 25372 6443
rect 25320 6400 25372 6409
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 15752 6196 15804 6248
rect 15292 6128 15344 6180
rect 17500 6196 17552 6248
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 17408 6128 17460 6180
rect 18604 6196 18656 6248
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 19064 6196 19116 6248
rect 20352 6239 20404 6248
rect 20352 6205 20361 6239
rect 20361 6205 20395 6239
rect 20395 6205 20404 6239
rect 20352 6196 20404 6205
rect 21272 6196 21324 6248
rect 25044 6171 25096 6180
rect 8668 6060 8720 6069
rect 9864 6060 9916 6112
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 15752 6060 15804 6112
rect 16764 6060 16816 6112
rect 17684 6060 17736 6112
rect 19248 6103 19300 6112
rect 19248 6069 19257 6103
rect 19257 6069 19291 6103
rect 19291 6069 19300 6103
rect 19248 6060 19300 6069
rect 20260 6103 20312 6112
rect 20260 6069 20269 6103
rect 20269 6069 20303 6103
rect 20303 6069 20312 6103
rect 20260 6060 20312 6069
rect 20904 6060 20956 6112
rect 22376 6060 22428 6112
rect 24032 6060 24084 6112
rect 25044 6137 25053 6171
rect 25053 6137 25087 6171
rect 25087 6137 25096 6171
rect 25044 6128 25096 6137
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 2044 5788 2096 5840
rect 1584 5720 1636 5772
rect 1768 5720 1820 5772
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2320 5652 2372 5704
rect 4160 5856 4212 5908
rect 6000 5856 6052 5908
rect 7564 5856 7616 5908
rect 7656 5856 7708 5908
rect 9312 5856 9364 5908
rect 9680 5856 9732 5908
rect 3516 5831 3568 5840
rect 3516 5797 3525 5831
rect 3525 5797 3559 5831
rect 3559 5797 3568 5831
rect 3516 5788 3568 5797
rect 3700 5788 3752 5840
rect 5356 5788 5408 5840
rect 6552 5788 6604 5840
rect 8208 5831 8260 5840
rect 8208 5797 8217 5831
rect 8217 5797 8251 5831
rect 8251 5797 8260 5831
rect 8208 5788 8260 5797
rect 11060 5856 11112 5908
rect 11428 5856 11480 5908
rect 12348 5856 12400 5908
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 14004 5856 14056 5908
rect 14556 5856 14608 5908
rect 15844 5856 15896 5908
rect 16396 5856 16448 5908
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 24124 5856 24176 5908
rect 10232 5788 10284 5840
rect 3240 5720 3292 5772
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 6920 5720 6972 5772
rect 11980 5720 12032 5772
rect 13820 5763 13872 5772
rect 13820 5729 13829 5763
rect 13829 5729 13863 5763
rect 13863 5729 13872 5763
rect 13820 5720 13872 5729
rect 15292 5720 15344 5772
rect 17868 5788 17920 5840
rect 20352 5831 20404 5840
rect 20352 5797 20361 5831
rect 20361 5797 20395 5831
rect 20395 5797 20404 5831
rect 20352 5788 20404 5797
rect 22376 5788 22428 5840
rect 24952 5831 25004 5840
rect 24952 5797 24961 5831
rect 24961 5797 24995 5831
rect 24995 5797 25004 5831
rect 24952 5788 25004 5797
rect 15660 5720 15712 5772
rect 16396 5763 16448 5772
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 5264 5652 5316 5704
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 9496 5652 9548 5704
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 14556 5652 14608 5704
rect 16396 5729 16405 5763
rect 16405 5729 16439 5763
rect 16439 5729 16448 5763
rect 16396 5720 16448 5729
rect 16580 5720 16632 5772
rect 17592 5720 17644 5772
rect 17684 5763 17736 5772
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 17960 5720 18012 5772
rect 18604 5763 18656 5772
rect 16672 5652 16724 5704
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 18604 5729 18613 5763
rect 18613 5729 18647 5763
rect 18647 5729 18656 5763
rect 18604 5720 18656 5729
rect 18972 5763 19024 5772
rect 18972 5729 18981 5763
rect 18981 5729 19015 5763
rect 19015 5729 19024 5763
rect 18972 5720 19024 5729
rect 20444 5720 20496 5772
rect 22192 5763 22244 5772
rect 22192 5729 22201 5763
rect 22201 5729 22235 5763
rect 22235 5729 22244 5763
rect 22192 5720 22244 5729
rect 18420 5652 18472 5704
rect 19248 5652 19300 5704
rect 25044 5652 25096 5704
rect 12532 5627 12584 5636
rect 12532 5593 12541 5627
rect 12541 5593 12575 5627
rect 12575 5593 12584 5627
rect 12532 5584 12584 5593
rect 13728 5584 13780 5636
rect 21456 5627 21508 5636
rect 21456 5593 21465 5627
rect 21465 5593 21499 5627
rect 21499 5593 21508 5627
rect 21456 5584 21508 5593
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 9128 5559 9180 5568
rect 9128 5525 9137 5559
rect 9137 5525 9171 5559
rect 9171 5525 9180 5559
rect 9128 5516 9180 5525
rect 15752 5516 15804 5568
rect 16120 5516 16172 5568
rect 21640 5516 21692 5568
rect 24216 5516 24268 5568
rect 24676 5516 24728 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2044 5355 2096 5364
rect 2044 5321 2053 5355
rect 2053 5321 2087 5355
rect 2087 5321 2096 5355
rect 2044 5312 2096 5321
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 6000 5312 6052 5364
rect 8208 5312 8260 5364
rect 10232 5312 10284 5364
rect 13636 5355 13688 5364
rect 13636 5321 13645 5355
rect 13645 5321 13679 5355
rect 13679 5321 13688 5355
rect 13636 5312 13688 5321
rect 7288 5244 7340 5296
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 11888 5244 11940 5253
rect 15660 5287 15712 5296
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 4528 5176 4580 5228
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 5356 5176 5408 5228
rect 7564 5176 7616 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 10048 5219 10100 5228
rect 9128 5176 9180 5185
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 10784 5176 10836 5228
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 15660 5253 15669 5287
rect 15669 5253 15703 5287
rect 15703 5253 15712 5287
rect 15660 5244 15712 5253
rect 16120 5244 16172 5296
rect 18972 5312 19024 5364
rect 19340 5312 19392 5364
rect 22192 5312 22244 5364
rect 24952 5287 25004 5296
rect 1492 5108 1544 5160
rect 12256 5151 12308 5160
rect 12256 5117 12265 5151
rect 12265 5117 12299 5151
rect 12299 5117 12308 5151
rect 12992 5151 13044 5160
rect 12256 5108 12308 5117
rect 12992 5117 13001 5151
rect 13001 5117 13035 5151
rect 13035 5117 13044 5151
rect 12992 5108 13044 5117
rect 13820 5108 13872 5160
rect 14556 5151 14608 5160
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 3700 5040 3752 5092
rect 6920 5040 6972 5092
rect 8484 5083 8536 5092
rect 8484 5049 8493 5083
rect 8493 5049 8527 5083
rect 8527 5049 8536 5083
rect 8484 5040 8536 5049
rect 4252 5015 4304 5024
rect 2504 4972 2556 4981
rect 4252 4981 4261 5015
rect 4261 4981 4295 5015
rect 4295 4981 4304 5015
rect 4252 4972 4304 4981
rect 9404 5040 9456 5092
rect 9864 5040 9916 5092
rect 14096 5083 14148 5092
rect 14096 5049 14105 5083
rect 14105 5049 14139 5083
rect 14139 5049 14148 5083
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 17960 5176 18012 5228
rect 16120 5151 16172 5160
rect 14096 5040 14148 5049
rect 16120 5117 16129 5151
rect 16129 5117 16163 5151
rect 16163 5117 16172 5151
rect 16120 5108 16172 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 24952 5253 24961 5287
rect 24961 5253 24995 5287
rect 24995 5253 25004 5287
rect 24952 5244 25004 5253
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 21456 5176 21508 5228
rect 24124 5176 24176 5228
rect 20536 5108 20588 5160
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 20352 5083 20404 5092
rect 20352 5049 20361 5083
rect 20361 5049 20395 5083
rect 20395 5049 20404 5083
rect 20352 5040 20404 5049
rect 22376 5083 22428 5092
rect 11980 4972 12032 5024
rect 14188 4972 14240 5024
rect 15844 4972 15896 5024
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 17684 4972 17736 5024
rect 20904 4972 20956 5024
rect 22376 5049 22385 5083
rect 22385 5049 22419 5083
rect 22419 5049 22428 5083
rect 22376 5040 22428 5049
rect 23848 5040 23900 5092
rect 22652 4972 22704 5024
rect 24216 5015 24268 5024
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 24216 4972 24268 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1400 4768 1452 4820
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 3148 4768 3200 4820
rect 3700 4768 3752 4820
rect 4528 4768 4580 4820
rect 8484 4768 8536 4820
rect 9864 4768 9916 4820
rect 10140 4768 10192 4820
rect 1768 4700 1820 4752
rect 2228 4743 2280 4752
rect 2228 4709 2237 4743
rect 2237 4709 2271 4743
rect 2271 4709 2280 4743
rect 2228 4700 2280 4709
rect 2688 4700 2740 4752
rect 2964 4700 3016 4752
rect 4160 4700 4212 4752
rect 4804 4743 4856 4752
rect 4804 4709 4813 4743
rect 4813 4709 4847 4743
rect 4847 4709 4856 4743
rect 4804 4700 4856 4709
rect 7196 4743 7248 4752
rect 7196 4709 7205 4743
rect 7205 4709 7239 4743
rect 7239 4709 7248 4743
rect 7196 4700 7248 4709
rect 7288 4743 7340 4752
rect 7288 4709 7297 4743
rect 7297 4709 7331 4743
rect 7331 4709 7340 4743
rect 12532 4768 12584 4820
rect 16672 4768 16724 4820
rect 17224 4768 17276 4820
rect 18880 4768 18932 4820
rect 19432 4768 19484 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 23204 4768 23256 4820
rect 24216 4768 24268 4820
rect 25044 4811 25096 4820
rect 25044 4777 25053 4811
rect 25053 4777 25087 4811
rect 25087 4777 25096 4811
rect 25044 4768 25096 4777
rect 7288 4700 7340 4709
rect 10784 4743 10836 4752
rect 10784 4709 10793 4743
rect 10793 4709 10827 4743
rect 10827 4709 10836 4743
rect 10784 4700 10836 4709
rect 15292 4700 15344 4752
rect 17960 4700 18012 4752
rect 20352 4700 20404 4752
rect 21364 4700 21416 4752
rect 22652 4743 22704 4752
rect 22652 4709 22661 4743
rect 22661 4709 22695 4743
rect 22695 4709 22704 4743
rect 22652 4700 22704 4709
rect 6092 4675 6144 4684
rect 6092 4641 6136 4675
rect 6136 4641 6144 4675
rect 12808 4675 12860 4684
rect 6092 4632 6144 4641
rect 12808 4641 12817 4675
rect 12817 4641 12851 4675
rect 12851 4641 12860 4675
rect 12808 4632 12860 4641
rect 14004 4632 14056 4684
rect 15752 4632 15804 4684
rect 15936 4675 15988 4684
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 16396 4632 16448 4684
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 17592 4675 17644 4684
rect 17592 4641 17601 4675
rect 17601 4641 17635 4675
rect 17635 4641 17644 4675
rect 17592 4632 17644 4641
rect 18052 4632 18104 4684
rect 24124 4675 24176 4684
rect 24124 4641 24133 4675
rect 24133 4641 24167 4675
rect 24167 4641 24176 4675
rect 24124 4632 24176 4641
rect 4436 4564 4488 4616
rect 6920 4564 6972 4616
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 13820 4564 13872 4616
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 21088 4564 21140 4616
rect 22284 4607 22336 4616
rect 22284 4573 22293 4607
rect 22293 4573 22327 4607
rect 22327 4573 22336 4607
rect 22284 4564 22336 4573
rect 23204 4564 23256 4616
rect 4252 4496 4304 4548
rect 5080 4496 5132 4548
rect 8760 4496 8812 4548
rect 9496 4496 9548 4548
rect 14280 4539 14332 4548
rect 14280 4505 14289 4539
rect 14289 4505 14323 4539
rect 14323 4505 14332 4539
rect 14280 4496 14332 4505
rect 20536 4496 20588 4548
rect 22376 4496 22428 4548
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 11704 4428 11756 4480
rect 12624 4471 12676 4480
rect 12624 4437 12633 4471
rect 12633 4437 12667 4471
rect 12667 4437 12676 4471
rect 12624 4428 12676 4437
rect 13728 4428 13780 4480
rect 14004 4471 14056 4480
rect 14004 4437 14013 4471
rect 14013 4437 14047 4471
rect 14047 4437 14056 4471
rect 14004 4428 14056 4437
rect 17776 4471 17828 4480
rect 17776 4437 17785 4471
rect 17785 4437 17819 4471
rect 17819 4437 17828 4471
rect 17776 4428 17828 4437
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 4160 4267 4212 4276
rect 4160 4233 4169 4267
rect 4169 4233 4203 4267
rect 4203 4233 4212 4267
rect 4160 4224 4212 4233
rect 4436 4267 4488 4276
rect 4436 4233 4445 4267
rect 4445 4233 4479 4267
rect 4479 4233 4488 4267
rect 4436 4224 4488 4233
rect 6092 4224 6144 4276
rect 12808 4224 12860 4276
rect 14004 4224 14056 4276
rect 17960 4224 18012 4276
rect 21364 4267 21416 4276
rect 21364 4233 21373 4267
rect 21373 4233 21407 4267
rect 21407 4233 21416 4267
rect 21364 4224 21416 4233
rect 22652 4224 22704 4276
rect 4344 4156 4396 4208
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 3424 4088 3476 4140
rect 17408 4156 17460 4208
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 9128 4131 9180 4140
rect 7840 4088 7892 4097
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 9496 4088 9548 4140
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 2412 4063 2464 4072
rect 2412 4029 2421 4063
rect 2421 4029 2455 4063
rect 2455 4029 2464 4063
rect 2412 4020 2464 4029
rect 6184 4020 6236 4072
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 12072 4020 12124 4072
rect 12808 4020 12860 4072
rect 15108 4020 15160 4072
rect 15752 4020 15804 4072
rect 15936 4088 15988 4140
rect 16396 4088 16448 4140
rect 18144 4088 18196 4140
rect 18972 4088 19024 4140
rect 16672 4020 16724 4072
rect 17224 4020 17276 4072
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 18420 4020 18472 4072
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 18880 4020 18932 4029
rect 20628 4088 20680 4140
rect 21088 4131 21140 4140
rect 21088 4097 21097 4131
rect 21097 4097 21131 4131
rect 21131 4097 21140 4131
rect 21088 4088 21140 4097
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22376 4131 22428 4140
rect 22100 4088 22152 4097
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 24124 4224 24176 4276
rect 25504 4088 25556 4140
rect 3148 3995 3200 4004
rect 3148 3961 3157 3995
rect 3157 3961 3191 3995
rect 3191 3961 3200 3995
rect 3148 3952 3200 3961
rect 6000 3952 6052 4004
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 7748 3952 7800 4004
rect 9220 3995 9272 4004
rect 9220 3961 9229 3995
rect 9229 3961 9263 3995
rect 9263 3961 9272 3995
rect 9220 3952 9272 3961
rect 9588 3952 9640 4004
rect 17868 3952 17920 4004
rect 18696 3952 18748 4004
rect 19524 3995 19576 4004
rect 19524 3961 19533 3995
rect 19533 3961 19567 3995
rect 19567 3961 19576 3995
rect 19524 3952 19576 3961
rect 20536 3995 20588 4004
rect 20536 3961 20545 3995
rect 20545 3961 20579 3995
rect 20579 3961 20588 3995
rect 20536 3952 20588 3961
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 19984 3884 20036 3936
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 2228 3723 2280 3732
rect 2228 3689 2237 3723
rect 2237 3689 2271 3723
rect 2271 3689 2280 3723
rect 2228 3680 2280 3689
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 3056 3680 3108 3732
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 5264 3680 5316 3732
rect 6092 3680 6144 3732
rect 9680 3680 9732 3732
rect 10692 3680 10744 3732
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 15108 3723 15160 3732
rect 15108 3689 15117 3723
rect 15117 3689 15151 3723
rect 15151 3689 15160 3723
rect 15108 3680 15160 3689
rect 15384 3723 15436 3732
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 16580 3680 16632 3732
rect 2136 3544 2188 3596
rect 3148 3544 3200 3596
rect 3976 3544 4028 3596
rect 5448 3612 5500 3664
rect 6000 3655 6052 3664
rect 6000 3621 6009 3655
rect 6009 3621 6043 3655
rect 6043 3621 6052 3655
rect 6000 3612 6052 3621
rect 6920 3612 6972 3664
rect 8116 3612 8168 3664
rect 8668 3612 8720 3664
rect 9588 3612 9640 3664
rect 11152 3655 11204 3664
rect 11152 3621 11161 3655
rect 11161 3621 11195 3655
rect 11195 3621 11204 3655
rect 11152 3612 11204 3621
rect 11704 3655 11756 3664
rect 11704 3621 11713 3655
rect 11713 3621 11747 3655
rect 11747 3621 11756 3655
rect 11704 3612 11756 3621
rect 12624 3612 12676 3664
rect 14004 3612 14056 3664
rect 16396 3612 16448 3664
rect 4620 3544 4672 3596
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 6828 3544 6880 3596
rect 7380 3587 7432 3596
rect 7380 3553 7389 3587
rect 7389 3553 7423 3587
rect 7423 3553 7432 3587
rect 7380 3544 7432 3553
rect 8944 3544 8996 3596
rect 10048 3544 10100 3596
rect 14372 3544 14424 3596
rect 15108 3544 15160 3596
rect 15936 3587 15988 3596
rect 15936 3553 15945 3587
rect 15945 3553 15979 3587
rect 15979 3553 15988 3587
rect 15936 3544 15988 3553
rect 16212 3587 16264 3596
rect 16212 3553 16221 3587
rect 16221 3553 16255 3587
rect 16255 3553 16264 3587
rect 16212 3544 16264 3553
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 17684 3587 17736 3596
rect 17684 3553 17693 3587
rect 17693 3553 17727 3587
rect 17727 3553 17736 3587
rect 17684 3544 17736 3553
rect 18420 3612 18472 3664
rect 18512 3587 18564 3596
rect 18512 3553 18521 3587
rect 18521 3553 18555 3587
rect 18555 3553 18564 3587
rect 18512 3544 18564 3553
rect 19524 3680 19576 3732
rect 20536 3680 20588 3732
rect 22100 3723 22152 3732
rect 22100 3689 22109 3723
rect 22109 3689 22143 3723
rect 22143 3689 22152 3723
rect 22100 3680 22152 3689
rect 21088 3655 21140 3664
rect 21088 3621 21097 3655
rect 21097 3621 21131 3655
rect 21131 3621 21140 3655
rect 21088 3612 21140 3621
rect 21916 3612 21968 3664
rect 22744 3612 22796 3664
rect 24032 3655 24084 3664
rect 24032 3621 24041 3655
rect 24041 3621 24075 3655
rect 24075 3621 24084 3655
rect 24032 3612 24084 3621
rect 19248 3544 19300 3596
rect 24676 3587 24728 3596
rect 24676 3553 24685 3587
rect 24685 3553 24719 3587
rect 24719 3553 24728 3587
rect 24676 3544 24728 3553
rect 6368 3476 6420 3528
rect 8300 3476 8352 3528
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 17868 3476 17920 3528
rect 19156 3519 19208 3528
rect 19156 3485 19165 3519
rect 19165 3485 19199 3519
rect 19199 3485 19208 3519
rect 19156 3476 19208 3485
rect 20076 3476 20128 3528
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 23020 3519 23072 3528
rect 4344 3451 4396 3460
rect 4344 3417 4353 3451
rect 4353 3417 4387 3451
rect 4387 3417 4396 3451
rect 4344 3408 4396 3417
rect 14280 3451 14332 3460
rect 14280 3417 14289 3451
rect 14289 3417 14323 3451
rect 14323 3417 14332 3451
rect 14280 3408 14332 3417
rect 18420 3408 18472 3460
rect 19524 3408 19576 3460
rect 20168 3408 20220 3460
rect 20720 3408 20772 3460
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 21456 3408 21508 3460
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 7288 3340 7340 3392
rect 8852 3383 8904 3392
rect 8852 3349 8861 3383
rect 8861 3349 8895 3383
rect 8895 3349 8904 3383
rect 8852 3340 8904 3349
rect 10508 3340 10560 3392
rect 10784 3340 10836 3392
rect 11520 3340 11572 3392
rect 12716 3340 12768 3392
rect 13728 3340 13780 3392
rect 14832 3340 14884 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1584 3179 1636 3188
rect 1584 3145 1593 3179
rect 1593 3145 1627 3179
rect 1627 3145 1636 3179
rect 1584 3136 1636 3145
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2136 3136 2188 3188
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 6460 3136 6512 3188
rect 8116 3136 8168 3188
rect 3516 3068 3568 3120
rect 5448 3068 5500 3120
rect 6276 3068 6328 3120
rect 7840 3111 7892 3120
rect 7840 3077 7849 3111
rect 7849 3077 7883 3111
rect 7883 3077 7892 3111
rect 7840 3068 7892 3077
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 5172 3000 5224 3052
rect 6000 3000 6052 3052
rect 6552 3000 6604 3052
rect 2044 2932 2096 2984
rect 2688 2932 2740 2984
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 7104 2932 7156 2984
rect 9220 3136 9272 3188
rect 9588 3136 9640 3188
rect 10048 3179 10100 3188
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 10508 3179 10560 3188
rect 10508 3145 10517 3179
rect 10517 3145 10551 3179
rect 10551 3145 10560 3179
rect 10508 3136 10560 3145
rect 12532 3136 12584 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13084 3111 13136 3120
rect 13084 3077 13093 3111
rect 13093 3077 13127 3111
rect 13127 3077 13136 3111
rect 13084 3068 13136 3077
rect 13820 3111 13872 3120
rect 13820 3077 13829 3111
rect 13829 3077 13863 3111
rect 13863 3077 13872 3111
rect 13820 3068 13872 3077
rect 15292 3136 15344 3188
rect 16212 3136 16264 3188
rect 17684 3179 17736 3188
rect 17684 3145 17693 3179
rect 17693 3145 17727 3179
rect 17727 3145 17736 3179
rect 17684 3136 17736 3145
rect 18052 3136 18104 3188
rect 19984 3136 20036 3188
rect 21088 3136 21140 3188
rect 21548 3136 21600 3188
rect 24676 3179 24728 3188
rect 24676 3145 24685 3179
rect 24685 3145 24719 3179
rect 24719 3145 24728 3179
rect 24676 3136 24728 3145
rect 25412 3179 25464 3188
rect 25412 3145 25421 3179
rect 25421 3145 25455 3179
rect 25455 3145 25464 3179
rect 25412 3136 25464 3145
rect 23848 3068 23900 3120
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 11704 3000 11756 3052
rect 14740 3043 14792 3052
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 16948 3000 17000 3052
rect 19156 3000 19208 3052
rect 22928 3000 22980 3052
rect 23020 3000 23072 3052
rect 14096 2932 14148 2984
rect 14556 2932 14608 2984
rect 15752 2975 15804 2984
rect 15752 2941 15761 2975
rect 15761 2941 15795 2975
rect 15795 2941 15804 2975
rect 15752 2932 15804 2941
rect 15936 2932 15988 2984
rect 16212 2932 16264 2984
rect 16580 2932 16632 2984
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 18420 2932 18472 2984
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 19248 2975 19300 2984
rect 19248 2941 19257 2975
rect 19257 2941 19291 2975
rect 19291 2941 19300 2975
rect 19248 2932 19300 2941
rect 22468 2975 22520 2984
rect 22468 2941 22477 2975
rect 22477 2941 22511 2975
rect 22511 2941 22520 2975
rect 22468 2932 22520 2941
rect 22836 2932 22888 2984
rect 10784 2907 10836 2916
rect 10784 2873 10793 2907
rect 10793 2873 10827 2907
rect 10827 2873 10836 2907
rect 10784 2864 10836 2873
rect 12808 2864 12860 2916
rect 11704 2839 11756 2848
rect 11704 2805 11713 2839
rect 11713 2805 11747 2839
rect 11747 2805 11756 2839
rect 11704 2796 11756 2805
rect 16764 2839 16816 2848
rect 16764 2805 16773 2839
rect 16773 2805 16807 2839
rect 16807 2805 16816 2839
rect 16764 2796 16816 2805
rect 19248 2839 19300 2848
rect 19248 2805 19257 2839
rect 19257 2805 19291 2839
rect 19291 2805 19300 2839
rect 19248 2796 19300 2805
rect 19432 2796 19484 2848
rect 20904 2864 20956 2916
rect 22744 2864 22796 2916
rect 25688 2932 25740 2984
rect 23756 2907 23808 2916
rect 22652 2839 22704 2848
rect 22652 2805 22661 2839
rect 22661 2805 22695 2839
rect 22695 2805 22704 2839
rect 22652 2796 22704 2805
rect 23756 2873 23765 2907
rect 23765 2873 23799 2907
rect 23799 2873 23808 2907
rect 23756 2864 23808 2873
rect 23848 2907 23900 2916
rect 23848 2873 23857 2907
rect 23857 2873 23891 2907
rect 23891 2873 23900 2907
rect 23848 2864 23900 2873
rect 23388 2796 23440 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2504 2635 2556 2644
rect 2504 2601 2513 2635
rect 2513 2601 2547 2635
rect 2547 2601 2556 2635
rect 2504 2592 2556 2601
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 6368 2635 6420 2644
rect 4712 2524 4764 2576
rect 4804 2499 4856 2508
rect 4804 2465 4813 2499
rect 4813 2465 4847 2499
rect 4847 2465 4856 2499
rect 4804 2456 4856 2465
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 6828 2592 6880 2644
rect 8760 2592 8812 2644
rect 9404 2592 9456 2644
rect 8208 2567 8260 2576
rect 8208 2533 8217 2567
rect 8217 2533 8251 2567
rect 8251 2533 8260 2567
rect 8208 2524 8260 2533
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 8300 2524 8352 2533
rect 9496 2456 9548 2508
rect 10692 2592 10744 2644
rect 11704 2592 11756 2644
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 15752 2592 15804 2644
rect 16672 2592 16724 2644
rect 17868 2592 17920 2644
rect 11152 2524 11204 2576
rect 11612 2567 11664 2576
rect 11612 2533 11621 2567
rect 11621 2533 11655 2567
rect 11655 2533 11664 2567
rect 11612 2524 11664 2533
rect 19432 2592 19484 2644
rect 19524 2592 19576 2644
rect 20996 2635 21048 2644
rect 20996 2601 21005 2635
rect 21005 2601 21039 2635
rect 21039 2601 21048 2635
rect 20996 2592 21048 2601
rect 22468 2592 22520 2644
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 25412 2635 25464 2644
rect 25412 2601 25421 2635
rect 25421 2601 25455 2635
rect 25455 2601 25464 2635
rect 25412 2592 25464 2601
rect 17960 2524 18012 2576
rect 18788 2567 18840 2576
rect 18788 2533 18791 2567
rect 18791 2533 18825 2567
rect 18825 2533 18840 2567
rect 18788 2524 18840 2533
rect 12716 2499 12768 2508
rect 12716 2465 12725 2499
rect 12725 2465 12759 2499
rect 12759 2465 12768 2499
rect 12716 2456 12768 2465
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 22192 2567 22244 2576
rect 22192 2533 22201 2567
rect 22201 2533 22235 2567
rect 22235 2533 22244 2567
rect 22192 2524 22244 2533
rect 23664 2524 23716 2576
rect 23848 2524 23900 2576
rect 23480 2456 23532 2508
rect 26148 2456 26200 2508
rect 8300 2388 8352 2440
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 15292 2388 15344 2440
rect 17408 2431 17460 2440
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 19248 2388 19300 2440
rect 21272 2431 21324 2440
rect 21272 2397 21281 2431
rect 21281 2397 21315 2431
rect 21315 2397 21324 2431
rect 21272 2388 21324 2397
rect 21456 2388 21508 2440
rect 3608 2320 3660 2372
rect 24860 2320 24912 2372
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 4436 2295 4488 2304
rect 4436 2261 4445 2295
rect 4445 2261 4479 2295
rect 4479 2261 4488 2295
rect 4436 2252 4488 2261
rect 10232 2252 10284 2304
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 26148 2295 26200 2304
rect 26148 2261 26157 2295
rect 26157 2261 26191 2295
rect 26191 2261 26200 2295
rect 26148 2252 26200 2261
rect 26424 2295 26476 2304
rect 26424 2261 26433 2295
rect 26433 2261 26467 2295
rect 26467 2261 26476 2295
rect 26424 2252 26476 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 2320 1232 2372 1284
rect 3608 1232 3660 1284
rect 7196 552 7248 604
rect 7932 552 7984 604
<< metal2 >>
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 24766 27432 24822 27441
rect 24766 27367 24822 27376
rect 1398 25392 1454 25401
rect 1398 25327 1454 25336
rect 1412 23662 1440 25327
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1214 23216 1270 23225
rect 1214 23151 1270 23160
rect 386 18320 442 18329
rect 386 18255 442 18264
rect 400 2972 428 18255
rect 1228 18222 1256 23151
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1412 19922 1440 21111
rect 1596 20398 1624 27367
rect 2594 26344 2650 26353
rect 2594 26279 2650 26288
rect 23478 26344 23534 26353
rect 23478 26279 23534 26288
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1412 19514 1440 19858
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1308 18352 1360 18358
rect 1308 18294 1360 18300
rect 1216 18216 1268 18222
rect 1216 18158 1268 18164
rect 1216 15700 1268 15706
rect 1216 15642 1268 15648
rect 1228 12481 1256 15642
rect 1214 12472 1270 12481
rect 1214 12407 1270 12416
rect 1320 11762 1348 18294
rect 1412 18057 1440 19246
rect 1596 18170 1624 20198
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1504 18142 1624 18170
rect 1398 18048 1454 18057
rect 1398 17983 1454 17992
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 17202 1440 17614
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 15910 1440 17138
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 13802 1440 15846
rect 1504 15706 1532 18142
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1400 13796 1452 13802
rect 1400 13738 1452 13744
rect 1490 12472 1546 12481
rect 1490 12407 1546 12416
rect 1400 12164 1452 12170
rect 1400 12106 1452 12112
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 570 9752 626 9761
rect 570 9687 626 9696
rect 584 8838 612 9687
rect 1412 8974 1440 12106
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 572 8832 624 8838
rect 572 8774 624 8780
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1412 4826 1440 8026
rect 1504 6746 1532 12407
rect 1596 12374 1624 18022
rect 1584 12368 1636 12374
rect 1584 12310 1636 12316
rect 1596 11898 1624 12310
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1688 11762 1716 18566
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1596 7970 1624 11698
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1688 10985 1716 11154
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1688 10810 1716 10911
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8090 1716 8978
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1596 7942 1716 7970
rect 1582 7712 1638 7721
rect 1582 7647 1638 7656
rect 1596 7546 1624 7647
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1504 6718 1624 6746
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 5166 1532 6598
rect 1596 5778 1624 6718
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1596 5370 1624 5607
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1412 4078 1440 4762
rect 1582 4584 1638 4593
rect 1582 4519 1638 4528
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1596 3738 1624 4519
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1688 3618 1716 7942
rect 1780 6746 1808 23462
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 1872 20262 1900 20946
rect 2134 20904 2190 20913
rect 2134 20839 2136 20848
rect 2188 20839 2190 20848
rect 2136 20810 2188 20816
rect 2044 20528 2096 20534
rect 2044 20470 2096 20476
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 1872 19417 1900 20198
rect 1858 19408 1914 19417
rect 1858 19343 1914 19352
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 18426 1992 18770
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1950 17776 2006 17785
rect 1950 17711 1952 17720
rect 2004 17711 2006 17720
rect 1952 17682 2004 17688
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1872 14482 1900 16934
rect 1964 16794 1992 17682
rect 2056 16794 2084 20470
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2134 19272 2190 19281
rect 2134 19207 2136 19216
rect 2188 19207 2190 19216
rect 2136 19178 2188 19184
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2148 16674 2176 18566
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 1964 16646 2176 16674
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1872 14006 1900 14418
rect 1860 14000 1912 14006
rect 1860 13942 1912 13948
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 1872 13190 1900 13738
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1860 12776 1912 12782
rect 1964 12753 1992 16646
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2134 16552 2190 16561
rect 2056 15706 2084 16526
rect 2134 16487 2190 16496
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 13462 2084 13670
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 1860 12718 1912 12724
rect 1950 12744 2006 12753
rect 1872 12102 1900 12718
rect 1950 12679 2006 12688
rect 2056 12646 2084 13398
rect 2044 12640 2096 12646
rect 1950 12608 2006 12617
rect 2044 12582 2096 12588
rect 1950 12543 2006 12552
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1964 11354 1992 12543
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2056 10538 2084 12582
rect 2148 12481 2176 16487
rect 2240 14618 2268 17614
rect 2332 16153 2360 19654
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2318 16144 2374 16153
rect 2318 16079 2374 16088
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 2332 15094 2360 15574
rect 2424 15502 2452 19110
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2240 13938 2268 14554
rect 2332 14521 2360 15030
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2318 14512 2374 14521
rect 2318 14447 2374 14456
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2332 13802 2360 14350
rect 2320 13796 2372 13802
rect 2320 13738 2372 13744
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12782 2268 13126
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2134 12472 2190 12481
rect 2134 12407 2190 12416
rect 2320 12368 2372 12374
rect 2226 12336 2282 12345
rect 2320 12310 2372 12316
rect 2226 12271 2282 12280
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1952 10056 2004 10062
rect 1858 10024 1914 10033
rect 1952 9998 2004 10004
rect 1858 9959 1914 9968
rect 1872 6882 1900 9959
rect 1964 9178 1992 9998
rect 2148 9897 2176 12038
rect 2240 11626 2268 12271
rect 2332 11898 2360 12310
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2424 11762 2452 14758
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2240 11354 2268 11562
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2516 11286 2544 19790
rect 2608 18426 2636 26279
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 2962 24304 3018 24313
rect 2962 24239 3018 24248
rect 2686 21992 2742 22001
rect 2686 21927 2742 21936
rect 2700 21010 2728 21927
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2792 20602 2820 20946
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2778 20088 2834 20097
rect 2778 20023 2834 20032
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2594 18320 2650 18329
rect 2594 18255 2650 18264
rect 2608 18222 2636 18255
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2516 10742 2544 11222
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2516 10198 2544 10474
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2134 9888 2190 9897
rect 2134 9823 2190 9832
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2148 9110 2176 9823
rect 2516 9450 2544 10134
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2226 9072 2282 9081
rect 2044 9036 2096 9042
rect 2226 9007 2282 9016
rect 2044 8978 2096 8984
rect 2056 7886 2084 8978
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1872 6854 1992 6882
rect 1860 6792 1912 6798
rect 1780 6740 1860 6746
rect 1780 6734 1912 6740
rect 1780 6718 1900 6734
rect 1872 5914 1900 6718
rect 1964 6662 1992 6854
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 2056 6186 2084 7142
rect 2044 6180 2096 6186
rect 2044 6122 2096 6128
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2056 5846 2084 6122
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1780 4758 1808 5714
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1964 4826 1992 5646
rect 2056 5370 2084 5782
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1768 4752 1820 4758
rect 1768 4694 1820 4700
rect 1964 4146 1992 4762
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1412 3590 1716 3618
rect 2148 3602 2176 8910
rect 2240 8430 2268 9007
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2240 7954 2268 8230
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2240 7002 2268 7890
rect 2332 7546 2360 7958
rect 2424 7818 2452 8366
rect 2516 8022 2544 9386
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2332 7206 2360 7482
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2332 6118 2360 6870
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2332 5710 2360 6054
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 2240 3738 2268 4694
rect 2424 4078 2452 7754
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2136 3596 2188 3602
rect 400 2944 520 2972
rect 492 480 520 2944
rect 1412 480 1440 3590
rect 2136 3538 2188 3544
rect 1582 3496 1638 3505
rect 1582 3431 1638 3440
rect 1596 3194 1624 3431
rect 2042 3224 2098 3233
rect 1584 3188 1636 3194
rect 2148 3194 2176 3538
rect 2042 3159 2044 3168
rect 1584 3130 1636 3136
rect 2096 3159 2098 3168
rect 2136 3188 2188 3194
rect 2044 3130 2096 3136
rect 2136 3130 2188 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2516 2650 2544 4966
rect 2608 4185 2636 18022
rect 2700 17542 2728 18770
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2700 16250 2728 16662
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15706 2728 15914
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2792 15162 2820 20023
rect 2976 19310 3004 24239
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 23492 23769 23520 26279
rect 23846 25392 23902 25401
rect 23846 25327 23902 25336
rect 13542 23760 13598 23769
rect 13542 23695 13544 23704
rect 13596 23695 13598 23704
rect 23478 23760 23534 23769
rect 23478 23695 23534 23704
rect 13544 23666 13596 23672
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 7102 20904 7158 20913
rect 7102 20839 7158 20848
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3148 20324 3200 20330
rect 3148 20266 3200 20272
rect 3160 19394 3188 20266
rect 3068 19366 3188 19394
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2976 16969 3004 17002
rect 2962 16960 3018 16969
rect 2962 16895 3018 16904
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 16114 2912 16526
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2884 15638 2912 16050
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2884 15026 2912 15574
rect 2976 15094 3004 15642
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2976 14618 3004 15030
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2686 14512 2742 14521
rect 3068 14498 3096 19366
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 2686 14447 2742 14456
rect 2884 14470 3096 14498
rect 2700 13818 2728 14447
rect 2700 13790 2820 13818
rect 2792 13530 2820 13790
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2700 12782 2728 13262
rect 2792 12986 2820 13466
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2688 12776 2740 12782
rect 2740 12736 2820 12764
rect 2688 12718 2740 12724
rect 2686 12472 2742 12481
rect 2792 12442 2820 12736
rect 2686 12407 2742 12416
rect 2780 12436 2832 12442
rect 2700 7478 2728 12407
rect 2780 12378 2832 12384
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2792 11257 2820 11834
rect 2778 11248 2834 11257
rect 2778 11183 2834 11192
rect 2792 10266 2820 11183
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2792 8634 2820 10202
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2688 4752 2740 4758
rect 2778 4720 2834 4729
rect 2740 4700 2778 4706
rect 2688 4694 2778 4700
rect 2700 4678 2778 4694
rect 2778 4655 2834 4664
rect 2686 4584 2742 4593
rect 2686 4519 2742 4528
rect 2594 4176 2650 4185
rect 2594 4111 2650 4120
rect 2700 3738 2728 4519
rect 2792 4146 2820 4655
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2700 2990 2728 3674
rect 2884 3176 2912 14470
rect 2962 13968 3018 13977
rect 3160 13954 3188 19110
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3344 18426 3372 18770
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3240 17128 3292 17134
rect 3292 17076 3372 17082
rect 3240 17070 3372 17076
rect 3252 17054 3372 17070
rect 3344 16833 3372 17054
rect 3330 16824 3386 16833
rect 3330 16759 3386 16768
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3252 14618 3280 14826
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3252 14074 3280 14554
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3160 13926 3280 13954
rect 2962 13903 3018 13912
rect 2976 13870 3004 13903
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11626 3004 12174
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2976 11082 3004 11562
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3160 10810 3188 11222
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3160 10266 3188 10746
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7274 3096 7686
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2976 6798 3004 7210
rect 3054 7168 3110 7177
rect 3054 7103 3110 7112
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 5234 3004 6734
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2976 4758 3004 5170
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 3068 3738 3096 7103
rect 3252 5778 3280 13926
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3160 4010 3188 4762
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3160 3194 3188 3538
rect 2792 3148 2912 3176
rect 3148 3188 3200 3194
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 1465 1624 2246
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 2320 1284 2372 1290
rect 2320 1226 2372 1232
rect 2332 480 2360 1226
rect 2792 513 2820 3148
rect 3148 3130 3200 3136
rect 2778 504 2834 513
rect 478 0 534 480
rect 1398 0 1454 480
rect 2318 0 2374 480
rect 3344 480 3372 16759
rect 3436 4146 3464 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 4344 19916 4396 19922
rect 4344 19858 4396 19864
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3528 12850 3556 18022
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3528 12442 3556 12786
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3528 9738 3556 11766
rect 3620 11642 3648 19246
rect 4356 19174 4384 19858
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 3884 18692 3936 18698
rect 3884 18634 3936 18640
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3712 11830 3740 17478
rect 3804 13274 3832 18022
rect 3896 14929 3924 18634
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3882 14920 3938 14929
rect 3882 14855 3938 14864
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 13394 3924 14758
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3882 13288 3938 13297
rect 3804 13246 3882 13274
rect 3882 13223 3938 13232
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3620 11614 3740 11642
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11286 3648 11494
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 9926 3648 10406
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3528 9710 3648 9738
rect 3514 9616 3570 9625
rect 3514 9551 3516 9560
rect 3568 9551 3570 9560
rect 3516 9522 3568 9528
rect 3620 7410 3648 9710
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3528 5846 3556 6666
rect 3712 6338 3740 11614
rect 3804 11354 3832 11698
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3620 6310 3740 6338
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3514 5672 3570 5681
rect 3514 5607 3570 5616
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3436 3738 3464 4082
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3528 3126 3556 5607
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3620 2378 3648 6310
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3712 5846 3740 6190
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3712 5370 3740 5782
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3712 5098 3740 5306
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3712 4826 3740 5034
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3804 2802 3832 10406
rect 3896 3233 3924 13223
rect 3988 12238 4016 16934
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4080 14618 4108 15370
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4172 14414 4200 18566
rect 4356 17105 4384 19110
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4342 17096 4398 17105
rect 4342 17031 4398 17040
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4250 16144 4306 16153
rect 4250 16079 4306 16088
rect 4264 15502 4292 16079
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4252 14544 4304 14550
rect 4250 14512 4252 14521
rect 4304 14512 4306 14521
rect 4250 14447 4306 14456
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4080 13841 4108 13874
rect 4066 13832 4122 13841
rect 4066 13767 4122 13776
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 12918 4108 13670
rect 4172 13530 4200 14350
rect 4264 14074 4292 14447
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4172 11558 4200 12310
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4264 11354 4292 12174
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4160 11280 4212 11286
rect 4158 11248 4160 11257
rect 4212 11248 4214 11257
rect 4158 11183 4214 11192
rect 4160 11144 4212 11150
rect 4080 11092 4160 11098
rect 4080 11086 4212 11092
rect 4080 11070 4200 11086
rect 4080 10266 4108 11070
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3988 9654 4016 10134
rect 4264 10062 4292 10950
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 8809 4108 9318
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4172 8090 4200 9862
rect 4264 9178 4292 9998
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4356 8498 4384 16594
rect 4448 15026 4476 18022
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4434 14920 4490 14929
rect 4434 14855 4490 14864
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7478 4200 7890
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3974 7304 4030 7313
rect 3974 7239 4030 7248
rect 3988 3602 4016 7239
rect 4080 6225 4108 7346
rect 4172 7206 4200 7414
rect 4160 7200 4212 7206
rect 4158 7168 4160 7177
rect 4212 7168 4214 7177
rect 4158 7103 4214 7112
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4172 6118 4200 6870
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4250 6624 4306 6633
rect 4250 6559 4306 6568
rect 4264 6458 4292 6559
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5914 4200 6054
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4066 4992 4122 5001
rect 4066 4927 4122 4936
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3882 3224 3938 3233
rect 3882 3159 3938 3168
rect 4080 2990 4108 4927
rect 4172 4758 4200 5850
rect 4356 5273 4384 6734
rect 4342 5264 4398 5273
rect 4342 5199 4398 5208
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4160 4752 4212 4758
rect 4264 4729 4292 4966
rect 4160 4694 4212 4700
rect 4250 4720 4306 4729
rect 4172 4282 4200 4694
rect 4250 4655 4306 4664
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 3804 2774 3924 2802
rect 3896 2553 3924 2774
rect 3882 2544 3938 2553
rect 3882 2479 3938 2488
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 3620 1290 3648 2314
rect 3608 1284 3660 1290
rect 3608 1226 3660 1232
rect 4264 480 4292 4490
rect 4356 4214 4384 5199
rect 4448 4622 4476 14855
rect 4540 5234 4568 19110
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4724 16794 4752 17478
rect 4816 16998 4844 17682
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 16046 4660 16526
rect 4724 16182 4752 16730
rect 4816 16561 4844 16934
rect 4802 16552 4858 16561
rect 4802 16487 4858 16496
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4802 15872 4858 15881
rect 4802 15807 4858 15816
rect 4816 15722 4844 15807
rect 4724 15694 4844 15722
rect 4724 13546 4752 15694
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4816 14550 4844 15438
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4724 13518 4844 13546
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4632 10033 4660 13194
rect 4724 12986 4752 13330
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4816 12866 4844 13518
rect 4724 12838 4844 12866
rect 4618 10024 4674 10033
rect 4618 9959 4674 9968
rect 4724 9654 4752 12838
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4816 12345 4844 12582
rect 4802 12336 4858 12345
rect 4802 12271 4858 12280
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4816 10810 4844 11222
rect 4908 11150 4936 16934
rect 5000 13190 5028 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 19174 5120 19246
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 5092 17241 5120 19110
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5184 18290 5212 18770
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5078 17232 5134 17241
rect 5078 17167 5134 17176
rect 5092 16232 5120 17167
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5092 16204 5212 16232
rect 5080 16108 5132 16114
rect 5080 16050 5132 16056
rect 5092 14890 5120 16050
rect 5184 15881 5212 16204
rect 5170 15872 5226 15881
rect 5170 15807 5226 15816
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5092 14278 5120 14826
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 13938 5120 14214
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5078 13696 5134 13705
rect 5078 13631 5134 13640
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 5000 10985 5028 12378
rect 4986 10976 5042 10985
rect 4986 10911 5042 10920
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5000 10169 5028 10911
rect 4986 10160 5042 10169
rect 4986 10095 5042 10104
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4908 8634 4936 8910
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5000 8294 5028 9046
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 6458 4752 6598
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4724 6254 4752 6394
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4816 5794 4844 7686
rect 5000 7546 5028 8230
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4894 7440 4950 7449
rect 4894 7375 4896 7384
rect 4948 7375 4950 7384
rect 4896 7346 4948 7352
rect 4908 7002 4936 7346
rect 5000 7274 5028 7482
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4986 6352 5042 6361
rect 4986 6287 5042 6296
rect 4724 5766 4844 5794
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4540 4826 4568 5170
rect 4618 5128 4674 5137
rect 4618 5063 4674 5072
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4448 4282 4476 4558
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4632 3602 4660 5063
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4356 3058 4384 3402
rect 4632 3194 4660 3538
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4724 2582 4752 5766
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 5234 4844 5646
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4816 4758 4844 5170
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 5000 3602 5028 6287
rect 5092 4554 5120 13631
rect 5184 10742 5212 15642
rect 5276 13530 5304 16594
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5276 12850 5304 13466
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5368 12442 5396 16934
rect 5460 14056 5488 18702
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5552 16232 5580 16526
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5552 16204 5764 16232
rect 5736 15910 5764 16204
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5644 15706 5672 15846
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5460 14028 5672 14056
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 13462 5488 13874
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13530 5580 13738
rect 5644 13705 5672 14028
rect 5630 13696 5686 13705
rect 5630 13631 5686 13640
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5460 12322 5488 13126
rect 5552 12442 5580 13262
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12866 6040 18090
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 15638 6132 17478
rect 6092 15632 6144 15638
rect 6092 15574 6144 15580
rect 6104 15162 6132 15574
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6104 14618 6132 14758
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 5644 12838 6040 12866
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5276 12294 5488 12322
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 9110 5212 10406
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5276 6730 5304 12294
rect 5448 12232 5500 12238
rect 5644 12186 5672 12838
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5736 12238 5764 12650
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5448 12174 5500 12180
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5368 10674 5396 11222
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 10130 5396 10474
rect 5460 10266 5488 12174
rect 5552 12158 5672 12186
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5460 9586 5488 10202
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5460 8498 5488 9522
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5552 7750 5580 12158
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11830 6040 12174
rect 6104 11898 6132 12242
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6090 11656 6146 11665
rect 5816 11620 5868 11626
rect 6090 11591 6146 11600
rect 5816 11562 5868 11568
rect 5828 11354 5856 11562
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6012 10198 6040 10610
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9586 6040 10134
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5828 9178 5856 9318
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 6012 9110 6040 9318
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5736 8090 5764 8502
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7546 6040 7890
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 6798 5396 7210
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 5368 6390 5396 6734
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5276 5710 5304 6122
rect 5368 5846 5396 6326
rect 5448 6180 5500 6186
rect 5552 6168 5580 7142
rect 5722 7032 5778 7041
rect 5722 6967 5778 6976
rect 5998 7032 6054 7041
rect 5998 6967 6054 6976
rect 5736 6866 5764 6967
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5736 6225 5764 6258
rect 5500 6140 5580 6168
rect 5722 6216 5778 6225
rect 5722 6151 5778 6160
rect 5448 6122 5500 6128
rect 6012 5914 6040 6967
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5368 5234 5396 5782
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5370 6040 5714
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 6104 4690 6132 11591
rect 6196 10674 6224 18022
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6288 17338 6316 17682
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6288 16096 6316 17274
rect 6288 16068 6408 16096
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6288 15638 6316 15914
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6288 14822 6316 15574
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6288 13802 6316 14486
rect 6380 13977 6408 16068
rect 6366 13968 6422 13977
rect 6366 13903 6422 13912
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6288 13462 6316 13738
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6288 12986 6316 13398
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6274 12744 6330 12753
rect 6274 12679 6330 12688
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10198 6224 10406
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 9178 6224 9998
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 7954 6224 8978
rect 6288 8634 6316 12679
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 10849 6408 11494
rect 6366 10840 6422 10849
rect 6366 10775 6422 10784
rect 6366 10024 6422 10033
rect 6366 9959 6422 9968
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 8566 6408 9959
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6274 8392 6330 8401
rect 6274 8327 6276 8336
rect 6328 8327 6330 8336
rect 6276 8298 6328 8304
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6196 7002 6224 7890
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6104 4282 6132 4626
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5170 3088 5226 3097
rect 5170 3023 5172 3032
rect 5224 3023 5226 3032
rect 5172 2994 5224 3000
rect 5184 2650 5212 2994
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4802 2544 4858 2553
rect 4802 2479 4804 2488
rect 4856 2479 4858 2488
rect 4804 2450 4856 2456
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4448 1601 4476 2246
rect 4434 1592 4490 1601
rect 4434 1527 4490 1536
rect 5276 480 5304 3674
rect 5460 3670 5488 3878
rect 6012 3670 6040 3946
rect 6104 3738 6132 4218
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 2990 5396 3334
rect 5460 3126 5488 3606
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 6012 3058 6040 3606
rect 6196 3369 6224 4014
rect 6368 3528 6420 3534
rect 6472 3516 6500 17614
rect 6932 17270 6960 18022
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 14521 6592 15846
rect 6550 14512 6606 14521
rect 6550 14447 6606 14456
rect 6564 13410 6592 14447
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6656 13530 6684 14350
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6564 13382 6684 13410
rect 6550 12336 6606 12345
rect 6550 12271 6606 12280
rect 6564 11898 6592 12271
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6564 11626 6592 11834
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6564 10470 6592 11222
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6550 10160 6606 10169
rect 6550 10095 6606 10104
rect 6564 6202 6592 10095
rect 6656 6662 6684 13382
rect 6748 12458 6776 16390
rect 6840 15910 6868 16594
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 14906 6868 15846
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6932 15026 6960 15438
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6840 14878 6960 14906
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13190 6868 13806
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6748 12430 6868 12458
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6748 7546 6776 11766
rect 6840 9654 6868 12430
rect 6932 11898 6960 14878
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7024 14074 7052 14826
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7116 13818 7144 20839
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 7470 18184 7526 18193
rect 7470 18119 7472 18128
rect 7524 18119 7526 18128
rect 7472 18090 7524 18096
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 13938 7236 14962
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7116 13790 7236 13818
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12850 7144 13126
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7012 12776 7064 12782
rect 7010 12744 7012 12753
rect 7064 12744 7066 12753
rect 7010 12679 7066 12688
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 11218 6960 11562
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10470 6960 10950
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 7024 9586 7052 12679
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 10606 7144 12582
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7116 9761 7144 10542
rect 7102 9752 7158 9761
rect 7102 9687 7158 9696
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6920 9376 6972 9382
rect 6826 9344 6882 9353
rect 6920 9318 6972 9324
rect 6826 9279 6882 9288
rect 6840 9110 6868 9279
rect 6932 9178 6960 9318
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8634 7052 8774
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7116 8022 7144 9590
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 6840 7818 6868 7958
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6840 7002 6868 7754
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6932 6458 6960 7142
rect 7116 7002 7144 7278
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7116 6254 7144 6938
rect 7104 6248 7156 6254
rect 6564 6174 6684 6202
rect 7104 6190 7156 6196
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6564 5846 6592 6054
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6564 5681 6592 5782
rect 6550 5672 6606 5681
rect 6550 5607 6606 5616
rect 6550 4176 6606 4185
rect 6550 4111 6552 4120
rect 6604 4111 6606 4120
rect 6552 4082 6604 4088
rect 6420 3488 6500 3516
rect 6368 3470 6420 3476
rect 6182 3360 6238 3369
rect 6182 3295 6238 3304
rect 6472 3194 6500 3488
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6276 3120 6328 3126
rect 6274 3088 6276 3097
rect 6328 3088 6330 3097
rect 6000 3052 6052 3058
rect 6564 3058 6592 4082
rect 6274 3023 6330 3032
rect 6552 3052 6604 3058
rect 6000 2994 6052 3000
rect 6552 2994 6604 3000
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 6656 2904 6684 6174
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5778 6960 6054
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5098 6960 5510
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 7208 4758 7236 13790
rect 7300 11762 7328 15846
rect 7392 12889 7420 17002
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7378 12880 7434 12889
rect 7378 12815 7434 12824
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7300 11354 7328 11698
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7300 9722 7328 11018
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7300 9178 7328 9454
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7300 7449 7328 8026
rect 7392 7993 7420 11834
rect 7378 7984 7434 7993
rect 7378 7919 7434 7928
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7300 6118 7328 6734
rect 7392 6458 7420 6802
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5302 7328 6054
rect 7288 5296 7340 5302
rect 7286 5264 7288 5273
rect 7340 5264 7342 5273
rect 7286 5199 7342 5208
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6932 3670 6960 4558
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6288 2876 6684 2904
rect 6288 2666 6316 2876
rect 6196 2638 6316 2666
rect 6366 2680 6422 2689
rect 6840 2650 6868 3538
rect 6932 3505 6960 3606
rect 6918 3496 6974 3505
rect 6918 3431 6974 3440
rect 7300 3398 7328 4694
rect 7484 4128 7512 16934
rect 7562 15056 7618 15065
rect 7562 14991 7618 15000
rect 7576 5914 7604 14991
rect 7668 13394 7696 18022
rect 8128 16046 8156 18294
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7852 14822 7880 15506
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7746 13968 7802 13977
rect 7746 13903 7802 13912
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7668 12782 7696 13330
rect 7760 12850 7788 13903
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7668 12374 7696 12718
rect 7852 12442 7880 14758
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7656 12368 7708 12374
rect 7944 12322 7972 15846
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 8036 14618 8064 15370
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8128 13433 8156 15846
rect 8114 13424 8170 13433
rect 8114 13359 8170 13368
rect 8114 13152 8170 13161
rect 8114 13087 8170 13096
rect 8128 12889 8156 13087
rect 8114 12880 8170 12889
rect 8024 12844 8076 12850
rect 8114 12815 8170 12824
rect 8024 12786 8076 12792
rect 7656 12310 7708 12316
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7852 12294 7972 12322
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7668 10538 7696 12174
rect 7760 11506 7788 12242
rect 7852 11694 7880 12294
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7840 11552 7892 11558
rect 7760 11500 7840 11506
rect 7760 11494 7892 11500
rect 7760 11478 7880 11494
rect 7746 10976 7802 10985
rect 7746 10911 7802 10920
rect 7760 10742 7788 10911
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7852 10606 7880 11478
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7668 9625 7696 10202
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7760 9874 7788 10066
rect 7852 10033 7880 10406
rect 7838 10024 7894 10033
rect 7838 9959 7894 9968
rect 7838 9888 7894 9897
rect 7760 9846 7838 9874
rect 7838 9823 7894 9832
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7654 9616 7710 9625
rect 7654 9551 7710 9560
rect 7654 9480 7710 9489
rect 7654 9415 7710 9424
rect 7668 5914 7696 9415
rect 7760 7410 7788 9658
rect 7852 9382 7880 9823
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 9081 7880 9318
rect 7838 9072 7894 9081
rect 7838 9007 7894 9016
rect 7944 8537 7972 12174
rect 7930 8528 7986 8537
rect 7930 8463 7986 8472
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7944 7750 7972 8366
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 8036 7562 8064 12786
rect 8114 11792 8170 11801
rect 8114 11727 8170 11736
rect 8128 11286 8156 11727
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8220 11150 8248 16662
rect 8312 15065 8340 17478
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8298 15056 8354 15065
rect 8298 14991 8354 15000
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8312 14074 8340 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8312 13462 8340 14010
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8312 12986 8340 13398
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8404 11370 8432 16934
rect 8482 16824 8538 16833
rect 8482 16759 8538 16768
rect 8496 16658 8524 16759
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16250 8524 16594
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8496 14074 8524 14418
rect 8588 14396 8616 18226
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 12162 17776 12218 17785
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 9956 17740 10008 17746
rect 12162 17711 12218 17720
rect 9956 17682 10008 17688
rect 8956 16998 8984 17682
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9034 17096 9090 17105
rect 9034 17031 9036 17040
rect 9088 17031 9090 17040
rect 9036 17002 9088 17008
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 9126 16960 9182 16969
rect 8666 15736 8722 15745
rect 8666 15671 8722 15680
rect 8680 14550 8708 15671
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8588 14368 8708 14396
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8574 13968 8630 13977
rect 8574 13903 8630 13912
rect 8588 13870 8616 13903
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8680 13569 8708 14368
rect 8758 13696 8814 13705
rect 8758 13631 8814 13640
rect 8666 13560 8722 13569
rect 8666 13495 8722 13504
rect 8576 12640 8628 12646
rect 8574 12608 8576 12617
rect 8628 12608 8630 12617
rect 8574 12543 8630 12552
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8496 11830 8524 12242
rect 8680 12170 8708 13495
rect 8772 12782 8800 13631
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8312 11342 8432 11370
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8220 10554 8248 10610
rect 8312 10554 8340 11342
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8220 10526 8340 10554
rect 8220 10130 8248 10526
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10124 8260 10130
rect 8128 10084 8208 10112
rect 8128 9722 8156 10084
rect 8208 10066 8260 10072
rect 8312 9738 8340 10406
rect 8404 10266 8432 11222
rect 8496 11082 8524 11766
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8680 9761 8708 10542
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8220 9710 8340 9738
rect 8666 9752 8722 9761
rect 8114 9480 8170 9489
rect 8114 9415 8170 9424
rect 8128 7886 8156 9415
rect 8220 8974 8248 9710
rect 8666 9687 8722 9696
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8206 8664 8262 8673
rect 8206 8599 8262 8608
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7944 7534 8064 7562
rect 8128 7546 8156 7822
rect 8116 7540 8168 7546
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7852 6322 7880 6734
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7576 5234 7604 5850
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7564 4140 7616 4146
rect 7484 4100 7564 4128
rect 7840 4140 7892 4146
rect 7616 4100 7788 4128
rect 7564 4082 7616 4088
rect 7760 4010 7788 4100
rect 7840 4082 7892 4088
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7378 3632 7434 3641
rect 7378 3567 7380 3576
rect 7432 3567 7434 3576
rect 7380 3538 7432 3544
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7116 2990 7144 3334
rect 7852 3126 7880 4082
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6196 480 6224 2638
rect 6366 2615 6368 2624
rect 6420 2615 6422 2624
rect 6828 2644 6880 2650
rect 6368 2586 6420 2592
rect 6828 2586 6880 2592
rect 7944 610 7972 7534
rect 8116 7482 8168 7488
rect 8220 5846 8248 8599
rect 8312 7546 8340 9386
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8312 7342 8340 7482
rect 8864 7342 8892 7890
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8496 7041 8524 7142
rect 8482 7032 8538 7041
rect 8482 6967 8538 6976
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8680 6118 8708 6326
rect 8772 6254 8800 6598
rect 8760 6248 8812 6254
rect 8758 6216 8760 6225
rect 8812 6216 8814 6225
rect 8758 6151 8814 6160
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5704 8168 5710
rect 8114 5672 8116 5681
rect 8168 5672 8170 5681
rect 8114 5607 8170 5616
rect 8220 5370 8248 5782
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8496 4826 8524 5034
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8680 3670 8708 6054
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8128 3194 8156 3606
rect 8300 3528 8352 3534
rect 8220 3505 8300 3516
rect 8206 3496 8300 3505
rect 8262 3488 8300 3496
rect 8300 3470 8352 3476
rect 8206 3431 8262 3440
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8022 2952 8078 2961
rect 8022 2887 8078 2896
rect 8036 1034 8064 2887
rect 8220 2582 8248 3431
rect 8772 2650 8800 4490
rect 8956 3602 8984 16934
rect 9126 16895 9182 16904
rect 9140 16046 9168 16895
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9600 16114 9628 16594
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9140 15706 9168 15982
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9128 15700 9180 15706
rect 9048 15660 9128 15688
rect 9048 13002 9076 15660
rect 9128 15642 9180 15648
rect 9126 15056 9182 15065
rect 9126 14991 9182 15000
rect 9140 13138 9168 14991
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9140 13110 9260 13138
rect 9048 12974 9168 13002
rect 9140 12306 9168 12974
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 4026 9076 11494
rect 9232 9654 9260 13110
rect 9324 12238 9352 14350
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9416 11218 9444 15846
rect 9600 15026 9628 16050
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9508 12442 9536 14826
rect 9600 14618 9628 14962
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9692 14482 9720 15438
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9784 13938 9812 16730
rect 9772 13932 9824 13938
rect 9692 13892 9772 13920
rect 9692 13546 9720 13892
rect 9772 13874 9824 13880
rect 9600 13530 9720 13546
rect 9588 13524 9720 13530
rect 9640 13518 9720 13524
rect 9770 13560 9826 13569
rect 9770 13495 9826 13504
rect 9588 13466 9640 13472
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9508 11762 9536 12378
rect 9692 12322 9720 13398
rect 9784 13297 9812 13495
rect 9770 13288 9826 13297
rect 9770 13223 9826 13232
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12442 9812 13126
rect 9876 12442 9904 17478
rect 9968 16998 9996 17682
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9692 12294 9904 12322
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 11354 9536 11494
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9416 10266 9444 11154
rect 9508 10810 9536 11290
rect 9600 11098 9628 11562
rect 9772 11144 9824 11150
rect 9600 11070 9720 11098
rect 9772 11086 9824 11092
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9508 9568 9536 10746
rect 9692 10674 9720 11070
rect 9784 10742 9812 11086
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9508 9540 9720 9568
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9496 9376 9548 9382
rect 9494 9344 9496 9353
rect 9548 9344 9550 9353
rect 9494 9279 9550 9288
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9324 8634 9352 9046
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9416 7546 9444 8366
rect 9508 8090 9536 8910
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9600 8072 9628 9386
rect 9692 9110 9720 9540
rect 9784 9178 9812 9998
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9680 8968 9732 8974
rect 9678 8936 9680 8945
rect 9732 8936 9734 8945
rect 9678 8871 9734 8880
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8344 9720 8774
rect 9770 8528 9826 8537
rect 9770 8463 9772 8472
rect 9824 8463 9826 8472
rect 9772 8434 9824 8440
rect 9772 8356 9824 8362
rect 9692 8316 9772 8344
rect 9772 8298 9824 8304
rect 9680 8084 9732 8090
rect 9600 8044 9680 8072
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9324 5914 9352 6734
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9140 5234 9168 5510
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9416 5098 9444 7482
rect 9600 6866 9628 8044
rect 9680 8026 9732 8032
rect 9784 7970 9812 8298
rect 9692 7942 9812 7970
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9692 5914 9720 7942
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9784 7002 9812 7686
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9876 6440 9904 12294
rect 9784 6412 9904 6440
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9678 5672 9734 5681
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9508 4554 9536 5646
rect 9678 5607 9734 5616
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4146 9168 4422
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9048 3998 9168 4026
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 3058 8892 3334
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8312 2446 8340 2518
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8864 1873 8892 2994
rect 8956 2961 8984 3538
rect 8942 2952 8998 2961
rect 8942 2887 8998 2896
rect 8850 1864 8906 1873
rect 8850 1799 8906 1808
rect 8036 1006 8156 1034
rect 7196 604 7248 610
rect 7196 546 7248 552
rect 7932 604 7984 610
rect 7932 546 7984 552
rect 7208 480 7236 546
rect 8128 480 8156 1006
rect 9140 480 9168 3998
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9232 3194 9260 3946
rect 9402 3496 9458 3505
rect 9402 3431 9458 3440
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9416 2650 9444 3431
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9508 2514 9536 4082
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9600 3670 9628 3946
rect 9692 3738 9720 5607
rect 9784 4146 9812 6412
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 5098 9904 6054
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9876 4826 9904 5034
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9600 2689 9628 3130
rect 9968 3074 9996 16934
rect 10060 13462 10088 17070
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10152 16250 10180 16594
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10152 15745 10180 16186
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10138 15736 10194 15745
rect 10289 15728 10585 15748
rect 10888 15745 10916 17002
rect 10874 15736 10930 15745
rect 10138 15671 10194 15680
rect 10874 15671 10930 15680
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 10152 14346 10180 15370
rect 10244 15201 10272 15574
rect 10230 15192 10286 15201
rect 10230 15127 10232 15136
rect 10284 15127 10286 15136
rect 10690 15192 10746 15201
rect 10690 15127 10746 15136
rect 10232 15098 10284 15104
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10232 14544 10284 14550
rect 10704 14498 10732 15127
rect 10232 14486 10284 14492
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 10152 12986 10180 14282
rect 10244 13802 10272 14486
rect 10612 14470 10732 14498
rect 10876 14476 10928 14482
rect 10612 14006 10640 14470
rect 10876 14418 10928 14424
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13462 10732 14214
rect 10888 14006 10916 14418
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10232 13456 10284 13462
rect 10230 13424 10232 13433
rect 10692 13456 10744 13462
rect 10284 13424 10286 13433
rect 10692 13398 10744 13404
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 10230 13359 10286 13368
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10046 12880 10102 12889
rect 10244 12866 10272 13359
rect 10888 12918 10916 13398
rect 10876 12912 10928 12918
rect 10046 12815 10102 12824
rect 10152 12838 10272 12866
rect 10874 12880 10876 12889
rect 10928 12880 10930 12889
rect 10060 7018 10088 12815
rect 10152 12238 10180 12838
rect 10874 12815 10930 12824
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10612 11898 10640 12106
rect 10704 12102 10732 12650
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10324 11824 10376 11830
rect 10322 11792 10324 11801
rect 10376 11792 10378 11801
rect 10322 11727 10378 11736
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 10810 10732 12038
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 10266 10180 10610
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10416 10192 10468 10198
rect 10796 10180 10824 12310
rect 10416 10134 10468 10140
rect 10750 10152 10824 10180
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10336 9654 10364 9930
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10336 9432 10364 9590
rect 10428 9518 10456 10134
rect 10750 10112 10778 10152
rect 10750 10084 10824 10112
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10152 9404 10364 9432
rect 10152 7886 10180 9404
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 8974 10732 9930
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10598 8664 10654 8673
rect 10598 8599 10600 8608
rect 10652 8599 10654 8608
rect 10600 8570 10652 8576
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10152 7410 10180 7822
rect 10244 7546 10272 7958
rect 10704 7750 10732 8774
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10428 7274 10456 7686
rect 10796 7528 10824 10084
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9654 10916 9998
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10888 8634 10916 9386
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10874 7848 10930 7857
rect 10874 7783 10930 7792
rect 10704 7500 10824 7528
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10060 6990 10180 7018
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 5234 10088 5646
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10152 4826 10180 6990
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10244 5370 10272 5782
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10600 4072 10652 4078
rect 10598 4040 10600 4049
rect 10652 4040 10654 4049
rect 10598 3975 10654 3984
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3738 10732 7500
rect 10888 7478 10916 7783
rect 10876 7472 10928 7478
rect 10796 7432 10876 7460
rect 10796 5234 10824 7432
rect 10876 7414 10928 7420
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 6390 10916 6598
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10060 3194 10088 3538
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10520 3194 10548 3334
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 9968 3046 10088 3074
rect 10704 3058 10732 3674
rect 10796 3398 10824 4694
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10060 2802 10088 3046
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10796 2922 10824 3334
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10060 2774 10133 2802
rect 9586 2680 9642 2689
rect 10105 2666 10133 2774
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10690 2680 10746 2689
rect 9586 2615 9642 2624
rect 10060 2638 10133 2666
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9220 2440 9272 2446
rect 9218 2408 9220 2417
rect 9272 2408 9274 2417
rect 9218 2343 9274 2352
rect 10060 480 10088 2638
rect 10690 2615 10692 2624
rect 10744 2615 10746 2624
rect 10692 2586 10744 2592
rect 10980 2446 11008 17614
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 14890 11100 15370
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 11072 13326 11100 14826
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12646 11100 13126
rect 11164 12986 11192 17070
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 15144 11284 16934
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11348 15366 11376 15982
rect 11428 15972 11480 15978
rect 11428 15914 11480 15920
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11256 15116 11376 15144
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11256 14278 11284 14962
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 14074 11284 14214
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11164 12782 11192 12922
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12442 11100 12582
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11164 11937 11192 12718
rect 11150 11928 11206 11937
rect 11150 11863 11206 11872
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10470 11100 10950
rect 11164 10713 11192 11863
rect 11150 10704 11206 10713
rect 11150 10639 11206 10648
rect 11060 10464 11112 10470
rect 11058 10432 11060 10441
rect 11112 10432 11114 10441
rect 11058 10367 11114 10376
rect 11348 9994 11376 15116
rect 11440 14482 11468 15914
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11440 14074 11468 14418
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11440 12306 11468 13670
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11532 10266 11560 15982
rect 11900 15910 11928 16594
rect 12176 16572 12204 17711
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12256 16584 12308 16590
rect 12176 16544 12256 16572
rect 12176 16250 12204 16544
rect 12256 16526 12308 16532
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12176 16046 12204 16186
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11532 9897 11560 10202
rect 11518 9888 11574 9897
rect 11518 9823 11574 9832
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11072 8430 11100 9454
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11072 5914 11100 6190
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11164 5522 11192 8910
rect 11242 8392 11298 8401
rect 11242 8327 11298 8336
rect 11256 6322 11284 8327
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11440 7546 11468 7890
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11440 5914 11468 7482
rect 11716 6186 11744 11494
rect 11808 11218 11836 15642
rect 11900 15570 11928 15846
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 11900 14822 11928 15506
rect 12268 15162 12296 15506
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 11888 14816 11940 14822
rect 12268 14793 12296 14826
rect 11888 14758 11940 14764
rect 12254 14784 12310 14793
rect 11900 12753 11928 14758
rect 12254 14719 12310 14728
rect 12268 14618 12296 14719
rect 12360 14634 12388 16594
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16114 12480 16390
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12452 15570 12480 16050
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12714 15872 12770 15881
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12256 14612 12308 14618
rect 12360 14606 12480 14634
rect 12256 14554 12308 14560
rect 12452 13938 12480 14606
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12070 13016 12126 13025
rect 12070 12951 12126 12960
rect 12084 12753 12112 12951
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 11886 12744 11942 12753
rect 11886 12679 11942 12688
rect 12070 12744 12126 12753
rect 12360 12714 12388 12786
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12070 12679 12126 12688
rect 12348 12708 12400 12714
rect 11900 11529 11928 12679
rect 12348 12650 12400 12656
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12176 11540 12204 12242
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12256 11552 12308 11558
rect 11886 11520 11942 11529
rect 12176 11512 12256 11540
rect 12256 11494 12308 11500
rect 11886 11455 11942 11464
rect 12268 11286 12296 11494
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11808 10810 11836 11154
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 12268 10470 12296 11222
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 11794 10296 11850 10305
rect 11794 10231 11850 10240
rect 11808 9654 11836 10231
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 12084 9382 12112 10066
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9450 12204 9862
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11978 9072 12034 9081
rect 11978 9007 11980 9016
rect 12032 9007 12034 9016
rect 11980 8978 12032 8984
rect 11992 8090 12020 8978
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12084 6361 12112 9318
rect 12268 9110 12296 10406
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12268 8498 12296 9046
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7818 12204 8230
rect 12360 8090 12388 11766
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 6866 12204 7754
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12268 7206 12296 7482
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12176 6458 12204 6802
rect 12268 6730 12296 7142
rect 12360 6798 12388 7822
rect 12452 7546 12480 12718
rect 12544 12646 12572 13330
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12544 11354 12572 12310
rect 12636 11762 12664 15846
rect 12714 15807 12770 15816
rect 12728 15609 12756 15807
rect 12714 15600 12770 15609
rect 12714 15535 12770 15544
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12728 15026 12756 15302
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12728 14278 12756 14826
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12728 14074 12756 14214
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12636 11286 12664 11698
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12622 10840 12678 10849
rect 12622 10775 12678 10784
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12544 8498 12572 9114
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12544 7342 12572 8026
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6866 12480 7142
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12452 6662 12480 6802
rect 12636 6798 12664 10775
rect 12728 10577 12756 12582
rect 12714 10568 12770 10577
rect 12714 10503 12770 10512
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12728 8022 12756 9046
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12820 7546 12848 16934
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 13938 13032 14214
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13004 9654 13032 9930
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8022 12940 8774
rect 13004 8498 13032 9590
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 13004 7886 13032 8434
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12898 7304 12954 7313
rect 12898 7239 12954 7248
rect 12912 7206 12940 7239
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12070 6352 12126 6361
rect 12070 6287 12126 6296
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11992 5778 12020 6122
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11072 5494 11192 5522
rect 11072 3534 11100 5494
rect 11888 5296 11940 5302
rect 11886 5264 11888 5273
rect 11940 5264 11942 5273
rect 11886 5199 11942 5208
rect 11992 5030 12020 5714
rect 12268 5166 12296 6054
rect 12360 5914 12388 6190
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12452 5234 12480 6598
rect 12544 6254 12572 6666
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12544 5642 12572 6190
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11060 3528 11112 3534
rect 11058 3496 11060 3505
rect 11112 3496 11114 3505
rect 11058 3431 11114 3440
rect 11058 3360 11114 3369
rect 11058 3295 11114 3304
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 1737 10272 2246
rect 10230 1728 10286 1737
rect 10230 1663 10286 1672
rect 11072 480 11100 3295
rect 11164 2582 11192 3606
rect 11532 3398 11560 3878
rect 11624 3505 11652 4558
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 3670 11744 4422
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11610 3496 11666 3505
rect 11610 3431 11666 3440
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11624 2582 11652 3431
rect 11716 3058 11744 3606
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11716 2650 11744 2790
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 11992 480 12020 4966
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12544 4146 12572 4762
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12084 3738 12112 4014
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12636 3670 12664 4422
rect 12820 4282 12848 4626
rect 12912 4593 12940 6054
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12898 4584 12954 4593
rect 12898 4519 12954 4528
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12820 4078 12848 4218
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12624 3664 12676 3670
rect 12544 3624 12624 3652
rect 12544 3194 12572 3624
rect 12624 3606 12676 3612
rect 12624 3528 12676 3534
rect 12622 3496 12624 3505
rect 12676 3496 12678 3505
rect 12622 3431 12678 3440
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12728 2514 12756 3334
rect 12820 2922 12848 4014
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 13004 480 13032 5102
rect 13096 3534 13124 17070
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13280 14482 13308 16730
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 14006 13308 14418
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13280 12617 13308 13262
rect 13266 12608 13322 12617
rect 13266 12543 13322 12552
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11286 13308 11494
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13280 10810 13308 11222
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13372 10266 13400 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 23492 21593 23520 23462
rect 23570 23216 23626 23225
rect 23570 23151 23626 23160
rect 16486 21584 16542 21593
rect 16486 21519 16542 21528
rect 23478 21584 23534 21593
rect 23478 21519 23534 21528
rect 13450 21448 13506 21457
rect 13450 21383 13452 21392
rect 13504 21383 13506 21392
rect 13452 21354 13504 21360
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13556 16946 13584 21286
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14094 19952 14150 19961
rect 14094 19887 14150 19896
rect 14002 18184 14058 18193
rect 14002 18119 14058 18128
rect 13464 16918 13584 16946
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13188 9110 13216 10066
rect 13372 9586 13400 10202
rect 13464 10062 13492 16918
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13648 15434 13676 16594
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13832 15638 13860 15914
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13728 15496 13780 15502
rect 13726 15464 13728 15473
rect 13780 15464 13782 15473
rect 13636 15428 13688 15434
rect 13726 15399 13782 15408
rect 13636 15370 13688 15376
rect 13634 15192 13690 15201
rect 13832 15178 13860 15574
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13690 15150 13860 15178
rect 13634 15127 13636 15136
rect 13688 15127 13690 15136
rect 13636 15098 13688 15104
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13556 13802 13584 14486
rect 13924 13977 13952 15370
rect 13910 13968 13966 13977
rect 13910 13903 13966 13912
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13726 13560 13782 13569
rect 13726 13495 13782 13504
rect 13740 13326 13768 13495
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13556 12345 13584 12922
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13542 12336 13598 12345
rect 13542 12271 13598 12280
rect 13556 11801 13584 12271
rect 13542 11792 13598 11801
rect 13542 11727 13598 11736
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13556 9489 13584 9522
rect 13542 9480 13598 9489
rect 13542 9415 13598 9424
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13648 8090 13676 12650
rect 13740 12442 13768 13262
rect 13832 12986 13860 13398
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13924 12866 13952 13262
rect 13832 12838 13952 12866
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13728 11144 13780 11150
rect 13832 11132 13860 12838
rect 13780 11104 13860 11132
rect 13728 11086 13780 11092
rect 13832 11014 13860 11104
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10674 13860 10950
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13832 10266 13860 10610
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13924 10441 13952 10474
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13820 10124 13872 10130
rect 13924 10112 13952 10367
rect 13872 10084 13952 10112
rect 13820 10066 13872 10072
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9194 13860 9862
rect 13740 9178 13860 9194
rect 13728 9172 13860 9178
rect 13780 9166 13860 9172
rect 13728 9114 13780 9120
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13188 7002 13216 7958
rect 13360 7880 13412 7886
rect 13358 7848 13360 7857
rect 13412 7848 13414 7857
rect 13832 7834 13860 8502
rect 13358 7783 13414 7792
rect 13648 7806 13860 7834
rect 13648 7546 13676 7806
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13096 3126 13124 3470
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13280 2417 13308 7482
rect 13740 7449 13768 7686
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13542 6760 13598 6769
rect 13542 6695 13598 6704
rect 13556 5914 13584 6695
rect 13832 6254 13860 7142
rect 13924 6458 13952 8910
rect 14016 8498 14044 18119
rect 14108 10130 14136 19887
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 16210 18728 16266 18737
rect 16210 18663 16266 18672
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 16046 14412 16390
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14292 15910 14320 15982
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14384 15552 14412 15982
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14200 15524 14412 15552
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14108 9722 14136 10066
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9081 14136 9318
rect 14200 9178 14228 15524
rect 14476 14929 14504 15846
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 15026 14596 15302
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14462 14920 14518 14929
rect 14372 14884 14424 14890
rect 14462 14855 14518 14864
rect 14372 14826 14424 14832
rect 14384 14618 14412 14826
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14384 12714 14412 12815
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14292 12442 14320 12650
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 11694 14320 12242
rect 14384 11801 14412 12310
rect 14370 11792 14426 11801
rect 14370 11727 14426 11736
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14384 11286 14412 11727
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14370 9616 14426 9625
rect 14370 9551 14426 9560
rect 14384 9450 14412 9551
rect 14476 9518 14504 14855
rect 14568 12850 14596 14962
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14660 11762 14688 16050
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14554 11520 14610 11529
rect 14554 11455 14610 11464
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14094 9072 14150 9081
rect 14094 9007 14150 9016
rect 14278 9072 14334 9081
rect 14278 9007 14280 9016
rect 14332 9007 14334 9016
rect 14280 8978 14332 8984
rect 14292 8634 14320 8978
rect 14384 8974 14412 9386
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14476 8566 14504 9046
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14108 7478 14136 8026
rect 14384 8022 14412 8366
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14096 7472 14148 7478
rect 14148 7432 14320 7460
rect 14096 7414 14148 7420
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 7002 14044 7278
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14200 6497 14228 6802
rect 14186 6488 14242 6497
rect 13912 6452 13964 6458
rect 14186 6423 14242 6432
rect 13912 6394 13964 6400
rect 13924 6254 13952 6394
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 14094 6216 14150 6225
rect 14094 6151 14150 6160
rect 14108 6118 14136 6151
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13820 5772 13872 5778
rect 13648 5732 13820 5760
rect 13648 5409 13676 5732
rect 13820 5714 13872 5720
rect 13740 5642 13952 5658
rect 13728 5636 13952 5642
rect 13780 5630 13952 5636
rect 13728 5578 13780 5584
rect 13634 5400 13690 5409
rect 13634 5335 13636 5344
rect 13688 5335 13690 5344
rect 13636 5306 13688 5312
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13832 4622 13860 5102
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13740 3398 13768 4422
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13450 3224 13506 3233
rect 13450 3159 13452 3168
rect 13504 3159 13506 3168
rect 13452 3130 13504 3136
rect 13832 3126 13860 4558
rect 13820 3120 13872 3126
rect 13818 3088 13820 3097
rect 13872 3088 13874 3097
rect 13818 3023 13874 3032
rect 13634 2816 13690 2825
rect 13634 2751 13690 2760
rect 13648 2650 13676 2751
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13266 2408 13322 2417
rect 13266 2343 13322 2352
rect 13924 480 13952 5630
rect 14016 4690 14044 5850
rect 14186 5672 14242 5681
rect 14186 5607 14242 5616
rect 14200 5273 14228 5607
rect 14186 5264 14242 5273
rect 14186 5199 14242 5208
rect 14292 5137 14320 7432
rect 14476 7206 14504 7890
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14568 6254 14596 11455
rect 14646 10568 14702 10577
rect 14646 10503 14702 10512
rect 14660 7410 14688 10503
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14568 5914 14596 6190
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14556 5704 14608 5710
rect 14370 5672 14426 5681
rect 14556 5646 14608 5652
rect 14370 5607 14426 5616
rect 14094 5128 14150 5137
rect 14094 5063 14096 5072
rect 14148 5063 14150 5072
rect 14278 5128 14334 5137
rect 14278 5063 14334 5072
rect 14096 5034 14148 5040
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4282 14044 4422
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14016 3670 14044 4218
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14108 2650 14136 2926
rect 14200 2689 14228 4966
rect 14278 4584 14334 4593
rect 14278 4519 14280 4528
rect 14332 4519 14334 4528
rect 14280 4490 14332 4496
rect 14384 3602 14412 5607
rect 14568 5166 14596 5646
rect 14646 5264 14702 5273
rect 14646 5199 14702 5208
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14278 3496 14334 3505
rect 14278 3431 14280 3440
rect 14332 3431 14334 3440
rect 14280 3402 14332 3408
rect 14568 2990 14596 5102
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14186 2680 14242 2689
rect 14096 2644 14148 2650
rect 14186 2615 14242 2624
rect 14096 2586 14148 2592
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14292 2417 14320 2450
rect 14278 2408 14334 2417
rect 14278 2343 14334 2352
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 2009 14504 2246
rect 14462 2000 14518 2009
rect 14462 1935 14518 1944
rect 14660 762 14688 5199
rect 14752 3058 14780 17070
rect 16224 16794 16252 18663
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 15910 15332 16594
rect 15292 15904 15344 15910
rect 15752 15904 15804 15910
rect 15292 15846 15344 15852
rect 15474 15872 15530 15881
rect 15752 15846 15804 15852
rect 15474 15807 15530 15816
rect 15290 15464 15346 15473
rect 15290 15399 15346 15408
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 15162 15332 15399
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14385 14872 14826
rect 15304 14618 15332 15098
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 14830 14376 14886 14385
rect 14830 14311 14886 14320
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14830 13968 14886 13977
rect 14830 13903 14886 13912
rect 14844 12170 14872 13903
rect 15396 13870 15424 14758
rect 15488 14482 15516 15807
rect 15658 15736 15714 15745
rect 15658 15671 15714 15680
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15488 14249 15516 14418
rect 15474 14240 15530 14249
rect 15474 14175 15530 14184
rect 15488 14074 15516 14175
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15474 13968 15530 13977
rect 15474 13903 15476 13912
rect 15528 13903 15530 13912
rect 15476 13874 15528 13880
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 13190 15424 13670
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 14832 12164 14884 12170
rect 14832 12106 14884 12112
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 9586 14872 11630
rect 15028 11354 15056 11698
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10554 15332 12582
rect 15396 11626 15424 13126
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15488 11286 15516 13398
rect 15476 11280 15528 11286
rect 15382 11248 15438 11257
rect 15476 11222 15528 11228
rect 15382 11183 15438 11192
rect 15396 11150 15424 11183
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15396 10674 15424 11086
rect 15488 10810 15516 11222
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15672 10690 15700 15671
rect 15764 12617 15792 15846
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15856 15366 15884 15574
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15856 14890 15884 15302
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15856 14793 15884 14826
rect 15842 14784 15898 14793
rect 15842 14719 15898 14728
rect 15948 13870 15976 16730
rect 16120 16720 16172 16726
rect 16026 16688 16082 16697
rect 16120 16662 16172 16668
rect 16026 16623 16082 16632
rect 16040 15337 16068 16623
rect 16026 15328 16082 15337
rect 16026 15263 16082 15272
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 16028 13320 16080 13326
rect 16026 13288 16028 13297
rect 16080 13288 16082 13297
rect 16026 13223 16082 13232
rect 16040 12986 16068 13223
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15750 12608 15806 12617
rect 15750 12543 15806 12552
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15488 10662 15700 10690
rect 15120 10538 15332 10554
rect 15108 10532 15332 10538
rect 15160 10526 15332 10532
rect 15108 10474 15160 10480
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 10066
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15212 8906 15240 9318
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14844 7478 14872 8366
rect 15304 8362 15332 9454
rect 15396 8945 15424 10202
rect 15382 8936 15438 8945
rect 15382 8871 15438 8880
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 15304 7410 15332 7890
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6780 15240 7142
rect 15304 6934 15332 7346
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 15212 6752 15332 6780
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6186 15332 6752
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 4758 15332 5714
rect 15396 5681 15424 8774
rect 15488 6610 15516 10662
rect 15764 10554 15792 12543
rect 15934 12200 15990 12209
rect 15934 12135 15990 12144
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15856 10810 15884 11562
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15672 10526 15792 10554
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15580 8974 15608 10066
rect 15672 9110 15700 10526
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 9178 15792 10406
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15580 8838 15608 8910
rect 15568 8832 15620 8838
rect 15566 8800 15568 8809
rect 15620 8800 15622 8809
rect 15566 8735 15622 8744
rect 15672 7818 15700 9046
rect 15750 7984 15806 7993
rect 15750 7919 15806 7928
rect 15764 7886 15792 7919
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15672 6798 15700 7754
rect 15856 7750 15884 9454
rect 15948 9382 15976 12135
rect 16040 12102 16068 12786
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15934 9208 15990 9217
rect 15934 9143 15990 9152
rect 15948 9042 15976 9143
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15948 8430 15976 8978
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15948 7954 15976 8366
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 6866 15884 7686
rect 15948 7546 15976 7890
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15488 6582 15608 6610
rect 15382 5672 15438 5681
rect 15382 5607 15438 5616
rect 15580 4865 15608 6582
rect 15672 5778 15700 6734
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 6118 15792 6190
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15856 5914 15884 6802
rect 16040 6066 16068 12038
rect 15948 6038 16068 6066
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15660 5296 15712 5302
rect 15658 5264 15660 5273
rect 15712 5264 15714 5273
rect 15658 5199 15714 5208
rect 15566 4856 15622 4865
rect 15566 4791 15622 4800
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15198 4040 15254 4049
rect 15120 3738 15148 4014
rect 15198 3975 15254 3984
rect 15212 3942 15240 3975
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15120 3602 15148 3674
rect 15396 3641 15424 3674
rect 15382 3632 15438 3641
rect 15108 3596 15160 3602
rect 15382 3567 15438 3576
rect 15108 3538 15160 3544
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14844 3074 14872 3334
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 14922 3088 14978 3097
rect 14740 3052 14792 3058
rect 14844 3046 14922 3074
rect 14922 3023 14978 3032
rect 14740 2994 14792 3000
rect 14936 2650 14964 3023
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15304 2446 15332 3130
rect 15580 2514 15608 4791
rect 15764 4690 15792 5510
rect 15948 5386 15976 6038
rect 16132 5574 16160 16662
rect 16224 16114 16252 16730
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 14618 16252 15438
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16316 13954 16344 16934
rect 16500 15502 16528 21519
rect 23584 21457 23612 23151
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23570 21448 23626 21457
rect 23570 21383 23626 21392
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 23480 20800 23532 20806
rect 17590 20768 17646 20777
rect 17590 20703 17646 20712
rect 23478 20768 23480 20777
rect 23532 20768 23534 20777
rect 23478 20703 23534 20712
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16868 15502 16896 15914
rect 16960 15910 16988 16594
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16500 14074 16528 14486
rect 16868 14414 16896 15438
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16578 14104 16634 14113
rect 16488 14068 16540 14074
rect 16578 14039 16634 14048
rect 16488 14010 16540 14016
rect 16592 14006 16620 14039
rect 16580 14000 16632 14006
rect 16316 13926 16528 13954
rect 16580 13942 16632 13948
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12850 16344 13262
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16316 12481 16344 12786
rect 16302 12472 16358 12481
rect 16302 12407 16358 12416
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16224 11898 16252 12310
rect 16316 12238 16344 12407
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 6497 16252 11494
rect 16316 11354 16344 12174
rect 16408 11558 16436 13806
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16500 11234 16528 13926
rect 16868 13530 16896 14350
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16776 12986 16804 13398
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16960 12424 16988 15846
rect 17406 14920 17462 14929
rect 17406 14855 17462 14864
rect 17420 14482 17448 14855
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17040 14408 17092 14414
rect 17038 14376 17040 14385
rect 17092 14376 17094 14385
rect 17038 14311 17094 14320
rect 17420 14074 17448 14418
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 16960 12396 17080 12424
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11937 16804 12174
rect 16762 11928 16818 11937
rect 16762 11863 16818 11872
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16316 11206 16528 11234
rect 16316 9110 16344 11206
rect 16580 11144 16632 11150
rect 16500 11104 16580 11132
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16408 9654 16436 9862
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16408 9042 16436 9590
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16408 8430 16436 8978
rect 16396 8424 16448 8430
rect 16302 8392 16358 8401
rect 16396 8366 16448 8372
rect 16302 8327 16358 8336
rect 16210 6488 16266 6497
rect 16210 6423 16266 6432
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15948 5358 16068 5386
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15764 4078 15792 4626
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15764 2990 15792 4014
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 15764 2650 15792 2926
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 1601 15332 2382
rect 15752 2304 15804 2310
rect 15750 2272 15752 2281
rect 15804 2272 15806 2281
rect 15750 2207 15806 2216
rect 15290 1592 15346 1601
rect 15290 1527 15346 1536
rect 14660 734 14964 762
rect 14936 480 14964 734
rect 15856 480 15884 4966
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15948 4146 15976 4626
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15934 3632 15990 3641
rect 15934 3567 15936 3576
rect 15988 3567 15990 3576
rect 15936 3538 15988 3544
rect 15948 2990 15976 3538
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15948 2825 15976 2926
rect 15934 2816 15990 2825
rect 15934 2751 15990 2760
rect 16040 2417 16068 5358
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16132 5166 16160 5238
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16224 3602 16252 6326
rect 16316 6322 16344 8327
rect 16408 8090 16436 8366
rect 16500 8294 16528 11104
rect 16580 11086 16632 11092
rect 16776 10577 16804 11630
rect 16948 11552 17000 11558
rect 16946 11520 16948 11529
rect 17000 11520 17002 11529
rect 16946 11455 17002 11464
rect 16762 10568 16818 10577
rect 16762 10503 16818 10512
rect 16948 10464 17000 10470
rect 16946 10432 16948 10441
rect 17000 10432 17002 10441
rect 16946 10367 17002 10376
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16868 9042 16896 9522
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16592 8430 16620 8978
rect 16868 8498 16896 8978
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16592 8022 16620 8366
rect 16580 8016 16632 8022
rect 16632 7976 16712 8004
rect 16580 7958 16632 7964
rect 16578 7440 16634 7449
rect 16578 7375 16634 7384
rect 16592 7342 16620 7375
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16684 6866 16712 7976
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16776 7206 16804 7890
rect 16868 7818 16896 8434
rect 16960 7954 16988 10367
rect 17052 10010 17080 12396
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17144 10810 17172 11562
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17144 10130 17172 10746
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17052 9982 17172 10010
rect 17144 9518 17172 9982
rect 17236 9926 17264 13806
rect 17314 13696 17370 13705
rect 17314 13631 17370 13640
rect 17328 13530 17356 13631
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17328 13326 17356 13466
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17314 10704 17370 10713
rect 17314 10639 17370 10648
rect 17328 10033 17356 10639
rect 17420 10538 17448 11222
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17512 10266 17540 12922
rect 17604 12866 17632 20703
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 23676 18737 23704 22374
rect 23662 18728 23718 18737
rect 23662 18663 23718 18672
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19522 17232 19578 17241
rect 19522 17167 19578 17176
rect 18050 17096 18106 17105
rect 18050 17031 18106 17040
rect 17776 15632 17828 15638
rect 17774 15600 17776 15609
rect 17868 15632 17920 15638
rect 17828 15600 17830 15609
rect 17868 15574 17920 15580
rect 17774 15535 17830 15544
rect 17788 15162 17816 15535
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17880 15026 17908 15574
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17696 12986 17724 13398
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17880 12889 17908 14962
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17972 13977 18000 14554
rect 17958 13968 18014 13977
rect 17958 13903 18014 13912
rect 18064 12918 18092 17031
rect 18512 15904 18564 15910
rect 18788 15904 18840 15910
rect 18564 15864 18644 15892
rect 18512 15846 18564 15852
rect 18328 14816 18380 14822
rect 18512 14816 18564 14822
rect 18380 14776 18460 14804
rect 18328 14758 18380 14764
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18156 14006 18184 14418
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18052 12912 18104 12918
rect 17866 12880 17922 12889
rect 17604 12838 17724 12866
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17314 10024 17370 10033
rect 17314 9959 17370 9968
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 8090 17172 8502
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 17130 7304 17186 7313
rect 17130 7239 17132 7248
rect 17184 7239 17186 7248
rect 17132 7210 17184 7216
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16408 5914 16436 6802
rect 16776 6118 16804 7142
rect 16946 7032 17002 7041
rect 16946 6967 16948 6976
rect 17000 6967 17002 6976
rect 16948 6938 17000 6944
rect 17604 6798 17632 12718
rect 17696 12238 17724 12838
rect 18052 12854 18104 12860
rect 17866 12815 17922 12824
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18052 12640 18104 12646
rect 18156 12617 18184 12718
rect 18052 12582 18104 12588
rect 18142 12608 18198 12617
rect 17958 12472 18014 12481
rect 17958 12407 18014 12416
rect 17776 12368 17828 12374
rect 17774 12336 17776 12345
rect 17828 12336 17830 12345
rect 17774 12271 17830 12280
rect 17972 12238 18000 12407
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17696 11898 17724 12174
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6186 17448 6598
rect 17604 6458 17632 6734
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17500 6248 17552 6254
rect 17696 6236 17724 9862
rect 18064 9217 18092 12582
rect 18142 12543 18198 12552
rect 18156 12442 18184 12543
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11801 18184 12038
rect 18142 11792 18198 11801
rect 18248 11762 18276 13262
rect 18326 13152 18382 13161
rect 18326 13087 18382 13096
rect 18340 12481 18368 13087
rect 18432 12646 18460 14776
rect 18512 14758 18564 14764
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18326 12472 18382 12481
rect 18326 12407 18382 12416
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18142 11727 18144 11736
rect 18196 11727 18198 11736
rect 18236 11756 18288 11762
rect 18144 11698 18196 11704
rect 18236 11698 18288 11704
rect 18248 11150 18276 11698
rect 18432 11354 18460 12310
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18524 11234 18552 14758
rect 18432 11206 18552 11234
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18248 9994 18276 10474
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18340 9926 18368 10542
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18050 9208 18106 9217
rect 18050 9143 18106 9152
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8362 17908 8774
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17880 7750 17908 8298
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17880 7410 17908 7686
rect 18064 7546 18092 8230
rect 18156 7886 18184 9386
rect 18248 9042 18276 9454
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18248 8430 18276 8978
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18248 7954 18276 8366
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17552 6208 17724 6236
rect 17500 6190 17552 6196
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16408 5778 16436 5850
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16224 3194 16252 3538
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16224 2990 16252 3130
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16316 2553 16344 4966
rect 16408 4690 16436 5714
rect 16592 4690 16620 5714
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16684 4826 16712 5646
rect 16776 5522 16804 6054
rect 16856 5704 16908 5710
rect 16854 5672 16856 5681
rect 16908 5672 16910 5681
rect 16854 5607 16910 5616
rect 16776 5494 16896 5522
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16408 4146 16436 4626
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16408 3670 16436 4082
rect 16592 3738 16620 4626
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16592 3097 16620 3674
rect 16684 3602 16712 4014
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16578 3088 16634 3097
rect 16578 3023 16634 3032
rect 16592 2990 16620 3023
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16684 2650 16712 3538
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16302 2544 16358 2553
rect 16302 2479 16358 2488
rect 16026 2408 16082 2417
rect 16026 2343 16082 2352
rect 16776 1873 16804 2790
rect 16762 1864 16818 1873
rect 16762 1799 16818 1808
rect 16868 480 16896 5494
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17236 4078 17264 4762
rect 17420 4214 17448 6122
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17512 3074 17540 6190
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17590 5944 17646 5953
rect 17590 5879 17592 5888
rect 17644 5879 17646 5888
rect 17592 5850 17644 5856
rect 17604 5778 17632 5850
rect 17696 5778 17724 6054
rect 17880 5846 17908 7346
rect 17958 6488 18014 6497
rect 17958 6423 18014 6432
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17972 5778 18000 6423
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17696 5030 17724 5714
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17972 5137 18000 5170
rect 18064 5166 18092 7482
rect 18156 7206 18184 7822
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18052 5160 18104 5166
rect 17958 5128 18014 5137
rect 18052 5102 18104 5108
rect 17958 5063 18014 5072
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17590 4720 17646 4729
rect 17590 4655 17592 4664
rect 17644 4655 17646 4664
rect 17592 4626 17644 4632
rect 17696 3602 17724 4966
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4185 17816 4422
rect 17972 4282 18000 4694
rect 18064 4690 18092 5102
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17774 4176 17830 4185
rect 17774 4111 17830 4120
rect 17972 4026 18000 4218
rect 18156 4146 18184 7142
rect 18248 6866 18276 7890
rect 18340 7002 18368 9658
rect 18432 9586 18460 11206
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18524 9081 18552 10406
rect 18616 10266 18644 15864
rect 18788 15846 18840 15852
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18708 13530 18736 13806
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18708 12782 18736 13466
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18616 9518 18644 10202
rect 18708 9722 18736 12582
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18510 9072 18566 9081
rect 18510 9007 18566 9016
rect 18616 7954 18644 9454
rect 18800 9042 18828 15846
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18878 13560 18934 13569
rect 18878 13495 18880 13504
rect 18932 13495 18934 13504
rect 18880 13466 18932 13472
rect 18984 10112 19012 14758
rect 19076 11898 19104 15846
rect 19536 14482 19564 17167
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20994 16552 21050 16561
rect 20994 16487 21050 16496
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 19982 15056 20038 15065
rect 19982 14991 20038 15000
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 14090 19564 14418
rect 19536 14074 19656 14090
rect 19536 14068 19668 14074
rect 19536 14062 19616 14068
rect 19616 14010 19668 14016
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19168 12646 19196 13330
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19168 12481 19196 12582
rect 19154 12472 19210 12481
rect 19154 12407 19210 12416
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19260 11286 19288 12242
rect 19248 11280 19300 11286
rect 19352 11257 19380 12582
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11898 19472 12038
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19444 11626 19472 11834
rect 19432 11620 19484 11626
rect 19432 11562 19484 11568
rect 19248 11222 19300 11228
rect 19338 11248 19394 11257
rect 19338 11183 19394 11192
rect 19536 10554 19564 13942
rect 19996 13802 20024 14991
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19352 10526 19564 10554
rect 18984 10084 19104 10112
rect 18972 9988 19024 9994
rect 18972 9930 19024 9936
rect 18984 9042 19012 9930
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18800 8566 18828 8978
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18800 8430 18828 8502
rect 18984 8430 19012 8978
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18616 7206 18644 7890
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18616 6866 18644 7142
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18248 6662 18276 6802
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6254 18276 6598
rect 18510 6352 18566 6361
rect 18510 6287 18566 6296
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18432 4078 18460 5646
rect 18524 5234 18552 6287
rect 18616 6254 18644 6802
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18892 6254 18920 6734
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18984 5778 19012 6802
rect 19076 6254 19104 10084
rect 19352 9654 19380 10526
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 9654 19564 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19892 10192 19944 10198
rect 19892 10134 19944 10140
rect 19982 10160 20038 10169
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19260 9518 19288 9590
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 9024 19288 9454
rect 19352 9178 19380 9590
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19340 9036 19392 9042
rect 19260 8996 19340 9024
rect 19340 8978 19392 8984
rect 19338 8800 19394 8809
rect 19338 8735 19394 8744
rect 19352 8634 19380 8735
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19444 8090 19472 9454
rect 19904 9364 19932 10134
rect 19982 10095 19984 10104
rect 20036 10095 20038 10104
rect 19984 10066 20036 10072
rect 19904 9336 20024 9364
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 8430 20024 9336
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19536 7954 19564 8366
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19536 7546 19564 7890
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19168 6848 19196 7278
rect 19444 7041 19472 7278
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19430 7032 19486 7041
rect 19622 7024 19918 7044
rect 19430 6967 19486 6976
rect 19340 6860 19392 6866
rect 19168 6820 19340 6848
rect 19340 6802 19392 6808
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19260 6497 19288 6666
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19246 6488 19302 6497
rect 19246 6423 19302 6432
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19246 6216 19302 6225
rect 19076 5953 19104 6190
rect 19246 6151 19302 6160
rect 19260 6118 19288 6151
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19062 5944 19118 5953
rect 19444 5914 19472 6598
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19062 5879 19118 5888
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18512 4480 18564 4486
rect 18616 4468 18644 5714
rect 18984 5370 19012 5714
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 18972 5364 19024 5370
rect 19260 5352 19288 5646
rect 19340 5364 19392 5370
rect 19260 5324 19340 5352
rect 18972 5306 19024 5312
rect 19340 5306 19392 5312
rect 18880 4820 18932 4826
rect 18984 4808 19012 5306
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 18932 4780 19012 4808
rect 19430 4856 19486 4865
rect 19622 4848 19918 4868
rect 19430 4791 19432 4800
rect 18880 4762 18932 4768
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18564 4440 18644 4468
rect 18512 4422 18564 4428
rect 17880 4010 18000 4026
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 17868 4004 18000 4010
rect 17920 3998 18000 4004
rect 17868 3946 17920 3952
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17696 3194 17724 3538
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 16948 3052 17000 3058
rect 17512 3046 17816 3074
rect 16948 2994 17000 3000
rect 16960 1737 16988 2994
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17420 2145 17448 2382
rect 17406 2136 17462 2145
rect 17406 2071 17462 2080
rect 16946 1728 17002 1737
rect 16946 1663 17002 1672
rect 17788 480 17816 3046
rect 17880 2650 17908 3470
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17972 2582 18000 3998
rect 18064 3194 18092 4014
rect 18432 3670 18460 4014
rect 18420 3664 18472 3670
rect 18418 3632 18420 3641
rect 18472 3632 18474 3641
rect 18524 3602 18552 4422
rect 18708 4010 18736 4558
rect 18984 4146 19012 4780
rect 19484 4791 19486 4800
rect 19432 4762 19484 4768
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18418 3567 18474 3576
rect 18512 3596 18564 3602
rect 18432 3466 18460 3567
rect 18512 3538 18564 3544
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18064 2990 18092 3130
rect 18432 2990 18460 3402
rect 18892 2990 18920 4014
rect 19524 4004 19576 4010
rect 19524 3946 19576 3952
rect 19536 3738 19564 3946
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 19168 3058 19196 3470
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19260 2990 19288 3538
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 18788 2576 18840 2582
rect 19260 2553 19288 2790
rect 19444 2650 19472 2790
rect 19536 2650 19564 3402
rect 19996 3194 20024 3878
rect 20088 3534 20116 15438
rect 20626 15328 20682 15337
rect 20626 15263 20682 15272
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20640 15042 20668 15263
rect 20180 10198 20208 15030
rect 20640 15014 20760 15042
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20168 10192 20220 10198
rect 20168 10134 20220 10140
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20180 9654 20208 9998
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20180 9178 20208 9590
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20272 8514 20300 14758
rect 20350 11656 20406 11665
rect 20350 11591 20352 11600
rect 20404 11591 20406 11600
rect 20352 11562 20404 11568
rect 20364 11286 20392 11562
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 9586 20392 10406
rect 20548 10198 20576 14758
rect 20640 12986 20668 15014
rect 20732 14958 20760 15014
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20720 14272 20772 14278
rect 20916 14249 20944 14418
rect 20720 14214 20772 14220
rect 20902 14240 20958 14249
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20640 12481 20668 12922
rect 20626 12472 20682 12481
rect 20626 12407 20682 12416
rect 20732 12186 20760 14214
rect 20902 14175 20958 14184
rect 20916 14074 20944 14175
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20812 12776 20864 12782
rect 20810 12744 20812 12753
rect 20864 12744 20866 12753
rect 20810 12679 20866 12688
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20640 12158 20760 12186
rect 20536 10192 20588 10198
rect 20536 10134 20588 10140
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20456 9518 20484 9862
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20272 8486 20484 8514
rect 20258 8392 20314 8401
rect 20258 8327 20260 8336
rect 20312 8327 20314 8336
rect 20260 8298 20312 8304
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20180 7342 20208 7686
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 6118 20300 7142
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20364 5846 20392 6190
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20456 5778 20484 8486
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20548 5250 20576 9998
rect 20456 5222 20576 5250
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20364 4758 20392 5034
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20180 3466 20208 3878
rect 20456 3618 20484 5222
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20548 4554 20576 5102
rect 20640 5012 20668 12158
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11801 20760 12038
rect 20718 11792 20774 11801
rect 20718 11727 20774 11736
rect 20824 11558 20852 12242
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20824 10577 20852 11494
rect 20810 10568 20866 10577
rect 20810 10503 20866 10512
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20824 9450 20852 9522
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20824 8294 20852 9386
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20824 7274 20852 8230
rect 20916 8129 20944 13670
rect 21008 13394 21036 16487
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23492 15609 23520 15846
rect 23478 15600 23534 15609
rect 23478 15535 23534 15544
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 21008 12986 21036 13330
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 21008 10810 21036 12582
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 20902 8120 20958 8129
rect 20902 8055 20958 8064
rect 20996 8016 21048 8022
rect 20916 7976 20996 8004
rect 20916 7274 20944 7976
rect 20996 7958 21048 7964
rect 21100 7886 21128 13126
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 20996 7472 21048 7478
rect 20994 7440 20996 7449
rect 21048 7440 21050 7449
rect 20994 7375 21050 7384
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20904 7268 20956 7274
rect 20904 7210 20956 7216
rect 20916 6866 20944 7210
rect 21008 7206 21036 7375
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21100 7002 21128 7822
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20916 6458 20944 6802
rect 21192 6746 21220 13806
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21284 11354 21312 11630
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21284 10742 21312 11290
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21284 10470 21312 10678
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10266 21312 10406
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21376 10146 21404 14010
rect 21100 6718 21220 6746
rect 21284 10118 21404 10146
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20720 5160 20772 5166
rect 20718 5128 20720 5137
rect 20772 5128 20774 5137
rect 20718 5063 20774 5072
rect 20916 5030 20944 6054
rect 20904 5024 20956 5030
rect 20640 4984 20760 5012
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20548 4010 20576 4490
rect 20640 4146 20668 4984
rect 20732 4826 20760 4984
rect 20904 4966 20956 4972
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20548 3738 20576 3946
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20456 3590 20760 3618
rect 20732 3466 20760 3590
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20916 2922 20944 4966
rect 21100 4706 21128 6718
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21192 5817 21220 6598
rect 21284 6254 21312 10118
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21376 9178 21404 9998
rect 21468 9761 21496 14758
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21454 9752 21510 9761
rect 21454 9687 21510 9696
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21560 7274 21588 14214
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21652 11286 21680 11494
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21652 10810 21680 11222
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21652 9466 21680 10202
rect 21744 9704 21772 15438
rect 23860 15042 23888 25327
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24674 24304 24730 24313
rect 24674 24239 24730 24248
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 24239
rect 24780 23866 24808 27367
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24780 23662 24808 23802
rect 24768 23656 24820 23662
rect 24768 23598 24820 23604
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24688 22574 24716 22714
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24674 22264 24730 22273
rect 24674 22199 24730 22208
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21010 24716 22199
rect 24766 21176 24822 21185
rect 24766 21111 24822 21120
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 20946
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24674 19136 24730 19145
rect 24674 19071 24730 19080
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24214 18048 24270 18057
rect 24214 17983 24270 17992
rect 23860 15014 24072 15042
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22006 14512 22062 14521
rect 22006 14447 22008 14456
rect 22060 14447 22062 14456
rect 22008 14418 22060 14424
rect 22020 14362 22048 14418
rect 21928 14334 22048 14362
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 21928 14074 21956 14334
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21824 11008 21876 11014
rect 21824 10950 21876 10956
rect 21836 10674 21864 10950
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21836 10062 21864 10610
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21824 9716 21876 9722
rect 21744 9676 21824 9704
rect 21824 9658 21876 9664
rect 21928 9654 21956 10134
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21652 9438 21864 9466
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 21652 7002 21680 8774
rect 21744 8362 21772 9046
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21744 6497 21772 6802
rect 21730 6488 21786 6497
rect 21730 6423 21732 6432
rect 21784 6423 21786 6432
rect 21732 6394 21784 6400
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21178 5808 21234 5817
rect 21178 5743 21234 5752
rect 21454 5672 21510 5681
rect 21454 5607 21456 5616
rect 21508 5607 21510 5616
rect 21456 5578 21508 5584
rect 21468 5234 21496 5578
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21008 4678 21128 4706
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21008 4622 21036 4678
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 21100 4146 21128 4558
rect 21376 4282 21404 4694
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21088 4140 21140 4146
rect 21140 4100 21312 4128
rect 21088 4082 21140 4088
rect 21088 3664 21140 3670
rect 21088 3606 21140 3612
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 21008 2650 21036 3470
rect 21100 3194 21128 3606
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 21284 2689 21312 4100
rect 21456 3460 21508 3466
rect 21456 3402 21508 3408
rect 21270 2680 21326 2689
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20996 2644 21048 2650
rect 21270 2615 21326 2624
rect 20996 2586 21048 2592
rect 18788 2518 18840 2524
rect 19246 2544 19302 2553
rect 18800 480 18828 2518
rect 19246 2479 19302 2488
rect 19260 2446 19288 2479
rect 21284 2446 21312 2615
rect 21468 2446 21496 3402
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 20718 2272 20774 2281
rect 20718 2207 20774 2216
rect 19706 2000 19762 2009
rect 19706 1935 19762 1944
rect 19720 480 19748 1935
rect 20732 480 20760 2207
rect 21560 2145 21588 3130
rect 21546 2136 21602 2145
rect 21546 2071 21602 2080
rect 21652 480 21680 5510
rect 21836 4593 21864 9438
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21928 8090 21956 8910
rect 22020 8378 22048 14214
rect 22098 12200 22154 12209
rect 22098 12135 22100 12144
rect 22152 12135 22154 12144
rect 22100 12106 22152 12112
rect 22098 12064 22154 12073
rect 22098 11999 22154 12008
rect 22112 11150 22140 11999
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22112 10810 22140 11086
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22020 8350 22140 8378
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22112 7954 22140 8350
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 22020 7478 22048 7754
rect 22008 7472 22060 7478
rect 21928 7432 22008 7460
rect 21822 4584 21878 4593
rect 21822 4519 21878 4528
rect 21928 3670 21956 7432
rect 22008 7414 22060 7420
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22112 7274 22140 7346
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22020 7002 22048 7210
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22204 6610 22232 14350
rect 22296 12442 22324 14758
rect 23952 14634 23980 14894
rect 23860 14606 23980 14634
rect 23570 14376 23626 14385
rect 23570 14311 23626 14320
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22296 11898 22324 12242
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22112 6582 22232 6610
rect 22112 4146 22140 6582
rect 22190 6216 22246 6225
rect 22190 6151 22246 6160
rect 22204 5778 22232 6151
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22204 5370 22232 5714
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22296 4842 22324 11834
rect 22480 9738 22508 12378
rect 22572 10266 22600 13670
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22664 10985 22692 12718
rect 22650 10976 22706 10985
rect 22650 10911 22706 10920
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22480 9710 22600 9738
rect 22572 8106 22600 9710
rect 22572 8078 22784 8106
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22572 7206 22600 7958
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22376 6112 22428 6118
rect 22480 6100 22508 6870
rect 22428 6072 22508 6100
rect 22376 6054 22428 6060
rect 22388 5846 22416 6054
rect 22376 5840 22428 5846
rect 22376 5782 22428 5788
rect 22388 5098 22416 5782
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22296 4814 22416 4842
rect 22284 4616 22336 4622
rect 22282 4584 22284 4593
rect 22336 4584 22338 4593
rect 22388 4554 22416 4814
rect 22664 4758 22692 4966
rect 22652 4752 22704 4758
rect 22652 4694 22704 4700
rect 22282 4519 22338 4528
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 22388 4146 22416 4490
rect 22664 4282 22692 4694
rect 22756 4570 22784 8078
rect 22848 6769 22876 13126
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 22834 6760 22890 6769
rect 22834 6695 22890 6704
rect 22756 4542 22876 4570
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22558 4176 22614 4185
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22376 4140 22428 4146
rect 22558 4111 22614 4120
rect 22376 4082 22428 4088
rect 22112 3738 22140 4082
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 21916 3664 21968 3670
rect 21916 3606 21968 3612
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22480 2650 22508 2926
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22192 2576 22244 2582
rect 22190 2544 22192 2553
rect 22244 2544 22246 2553
rect 22190 2479 22246 2488
rect 22572 1442 22600 4111
rect 22744 3664 22796 3670
rect 22744 3606 22796 3612
rect 22756 2922 22784 3606
rect 22848 2990 22876 4542
rect 22940 3058 22968 12038
rect 23018 11928 23074 11937
rect 23018 11863 23074 11872
rect 23032 11014 23060 11863
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 23032 10810 23060 10950
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23124 10554 23152 13806
rect 23032 10526 23152 10554
rect 23032 3534 23060 10526
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 23124 7857 23152 10406
rect 23216 9654 23244 14214
rect 23584 13394 23612 14311
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23400 12986 23428 13330
rect 23478 13288 23534 13297
rect 23478 13223 23480 13232
rect 23532 13223 23534 13232
rect 23480 13194 23532 13200
rect 23584 12986 23612 13330
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23400 12730 23428 12922
rect 23308 12702 23428 12730
rect 23478 12744 23534 12753
rect 23308 9994 23336 12702
rect 23478 12679 23534 12688
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23400 10266 23428 12582
rect 23492 11801 23520 12679
rect 23768 12073 23796 13874
rect 23754 12064 23810 12073
rect 23754 11999 23810 12008
rect 23478 11792 23534 11801
rect 23478 11727 23534 11736
rect 23480 11688 23532 11694
rect 23860 11642 23888 14606
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23952 13870 23980 14418
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23952 11762 23980 13806
rect 24044 13394 24072 15014
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24136 12594 24164 14758
rect 24228 14006 24256 17983
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14056 24716 19071
rect 24780 16250 24808 21111
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24780 16046 24808 16186
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 14074 24900 14418
rect 24860 14068 24912 14074
rect 24688 14028 24860 14056
rect 24860 14010 24912 14016
rect 24216 14000 24268 14006
rect 24216 13942 24268 13948
rect 24766 13968 24822 13977
rect 24766 13903 24822 13912
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24228 12986 24256 13126
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24044 12566 24164 12594
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23480 11630 23532 11636
rect 23492 10470 23520 11630
rect 23584 11614 23888 11642
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23480 10192 23532 10198
rect 23478 10160 23480 10169
rect 23532 10160 23534 10169
rect 23478 10095 23534 10104
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 23296 9716 23348 9722
rect 23400 9704 23428 9998
rect 23492 9722 23520 10095
rect 23348 9676 23428 9704
rect 23480 9716 23532 9722
rect 23296 9658 23348 9664
rect 23480 9658 23532 9664
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23478 9616 23534 9625
rect 23478 9551 23534 9560
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 23216 9178 23244 9454
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23308 7970 23336 9318
rect 23308 7942 23428 7970
rect 23296 7880 23348 7886
rect 23110 7848 23166 7857
rect 23296 7822 23348 7828
rect 23110 7783 23166 7792
rect 23204 7812 23256 7818
rect 23204 7754 23256 7760
rect 23216 4826 23244 7754
rect 23308 7002 23336 7822
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23400 6610 23428 7942
rect 23492 7410 23520 9551
rect 23584 8634 23612 11614
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23584 8362 23612 8570
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23570 7440 23626 7449
rect 23480 7404 23532 7410
rect 23570 7375 23626 7384
rect 23480 7346 23532 7352
rect 23478 7304 23534 7313
rect 23478 7239 23480 7248
rect 23532 7239 23534 7248
rect 23480 7210 23532 7216
rect 23308 6582 23428 6610
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23216 4622 23244 4762
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23032 3058 23060 3470
rect 23308 3097 23336 6582
rect 23388 6452 23440 6458
rect 23584 6440 23612 7375
rect 23440 6412 23612 6440
rect 23388 6394 23440 6400
rect 23570 3496 23626 3505
rect 23570 3431 23626 3440
rect 23294 3088 23350 3097
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 23020 3052 23072 3058
rect 23294 3023 23350 3032
rect 23020 2994 23072 3000
rect 22836 2984 22888 2990
rect 22836 2926 22888 2932
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22652 2848 22704 2854
rect 22650 2816 22652 2825
rect 23388 2848 23440 2854
rect 22704 2816 22706 2825
rect 23388 2790 23440 2796
rect 22650 2751 22706 2760
rect 23400 2530 23428 2790
rect 23400 2514 23520 2530
rect 23400 2508 23532 2514
rect 23400 2502 23480 2508
rect 23480 2450 23532 2456
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23032 1465 23060 2246
rect 23018 1456 23074 1465
rect 22572 1414 22692 1442
rect 22664 480 22692 1414
rect 23018 1391 23074 1400
rect 23584 480 23612 3431
rect 23676 2582 23704 11494
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23768 9586 23796 10202
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23860 9450 23888 10542
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 7750 23796 9318
rect 23860 9178 23888 9386
rect 23952 9330 23980 11086
rect 24044 9450 24072 12566
rect 24214 12472 24270 12481
rect 24214 12407 24270 12416
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24136 11694 24164 12242
rect 24124 11688 24176 11694
rect 24122 11656 24124 11665
rect 24176 11656 24178 11665
rect 24122 11591 24178 11600
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 9722 24164 11494
rect 24228 11218 24256 12407
rect 24780 12306 24808 13903
rect 24964 13433 24992 14758
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 24950 13424 25006 13433
rect 24950 13359 25006 13368
rect 25136 13388 25188 13394
rect 24964 12889 24992 13359
rect 25136 13330 25188 13336
rect 25148 12986 25176 13330
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 24950 12880 25006 12889
rect 24950 12815 25006 12824
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24780 11898 24808 12242
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24320 10996 24348 11630
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24412 11150 24440 11494
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24228 10968 24348 10996
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 23952 9302 24072 9330
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 23952 8566 23980 9114
rect 24044 8838 24072 9302
rect 24136 9110 24164 9522
rect 24124 9104 24176 9110
rect 24124 9046 24176 9052
rect 24228 8974 24256 10968
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11154
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24308 9648 24360 9654
rect 24308 9590 24360 9596
rect 24216 8968 24268 8974
rect 24320 8945 24348 9590
rect 24216 8910 24268 8916
rect 24306 8936 24362 8945
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23940 8560 23992 8566
rect 23940 8502 23992 8508
rect 23952 8430 23980 8502
rect 24228 8498 24256 8910
rect 24306 8871 24362 8880
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 23940 8424 23992 8430
rect 23846 8392 23902 8401
rect 23940 8366 23992 8372
rect 23846 8327 23902 8336
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23768 7002 23796 7346
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23860 5098 23888 8327
rect 23952 7954 23980 8366
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24044 8022 24072 8230
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 23952 7546 23980 7890
rect 24032 7812 24084 7818
rect 24032 7754 24084 7760
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24044 7410 24072 7754
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24136 6798 24164 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24216 6928 24268 6934
rect 24216 6870 24268 6876
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 24136 6458 24164 6734
rect 24228 6662 24256 6870
rect 24216 6656 24268 6662
rect 24216 6598 24268 6604
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 23848 5092 23900 5098
rect 23848 5034 23900 5040
rect 24044 3670 24072 6054
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24136 5234 24164 5850
rect 24228 5574 24256 6598
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 5681 24716 10610
rect 24780 8809 24808 10950
rect 24872 10606 24900 11018
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24964 10198 24992 12038
rect 25056 10849 25084 12650
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25042 10840 25098 10849
rect 25042 10775 25098 10784
rect 25148 10674 25176 12582
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 25226 10568 25282 10577
rect 25044 10532 25096 10538
rect 25226 10503 25282 10512
rect 25044 10474 25096 10480
rect 25056 10198 25084 10474
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 25044 10192 25096 10198
rect 25044 10134 25096 10140
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24766 8800 24822 8809
rect 24766 8735 24822 8744
rect 24674 5672 24730 5681
rect 24674 5607 24730 5616
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24676 5568 24728 5574
rect 24872 5522 24900 9318
rect 24964 9178 24992 10134
rect 25056 9722 25084 10134
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 25148 9586 25176 9998
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 24950 8936 25006 8945
rect 24950 8871 25006 8880
rect 24964 5846 24992 8871
rect 25148 8634 25176 9522
rect 25240 9518 25268 10503
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25226 8120 25282 8129
rect 25226 8055 25282 8064
rect 25240 7342 25268 8055
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 25056 6186 25084 6734
rect 25332 6458 25360 14214
rect 25596 13728 25648 13734
rect 25596 13670 25648 13676
rect 25502 12336 25558 12345
rect 25502 12271 25558 12280
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25424 9761 25452 10406
rect 25410 9752 25466 9761
rect 25410 9687 25466 9696
rect 25412 7200 25464 7206
rect 25412 7142 25464 7148
rect 25424 6633 25452 7142
rect 25410 6624 25466 6633
rect 25410 6559 25466 6568
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25044 6180 25096 6186
rect 25044 6122 25096 6128
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24676 5510 24728 5516
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24136 4690 24164 5170
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24228 4826 24256 4966
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 24136 4282 24164 4626
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24032 3664 24084 3670
rect 24032 3606 24084 3612
rect 24688 3602 24716 5510
rect 24780 5494 24900 5522
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3194 24716 3538
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 24674 3088 24730 3097
rect 23860 2922 23888 3062
rect 24674 3023 24730 3032
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 23848 2916 23900 2922
rect 23848 2858 23900 2864
rect 23768 2650 23796 2858
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23860 2582 23888 2858
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 23676 2009 23704 2518
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23662 2000 23718 2009
rect 23662 1935 23718 1944
rect 24688 1170 24716 3023
rect 24780 2553 24808 5494
rect 24964 5302 24992 5782
rect 25056 5710 25084 6122
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 25056 4826 25084 5646
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25410 4584 25466 4593
rect 25410 4519 25466 4528
rect 25424 3942 25452 4519
rect 25516 4146 25544 12271
rect 25608 8401 25636 13670
rect 25686 10024 25742 10033
rect 25686 9959 25742 9968
rect 25594 8392 25650 8401
rect 25594 8327 25650 8336
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 25502 4040 25558 4049
rect 25502 3975 25558 3984
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25410 3496 25466 3505
rect 25410 3431 25466 3440
rect 25424 3194 25452 3431
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 25410 2680 25466 2689
rect 25410 2615 25412 2624
rect 25464 2615 25466 2624
rect 25412 2586 25464 2592
rect 24766 2544 24822 2553
rect 24766 2479 24822 2488
rect 24858 2408 24914 2417
rect 24858 2343 24860 2352
rect 24912 2343 24914 2352
rect 24860 2314 24912 2320
rect 24596 1142 24716 1170
rect 24596 480 24624 1142
rect 25516 480 25544 3975
rect 25700 2990 25728 9959
rect 26514 5808 26570 5817
rect 26514 5743 26570 5752
rect 25688 2984 25740 2990
rect 25688 2926 25740 2932
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 26160 2310 26188 2450
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 26160 513 26188 2246
rect 26436 2009 26464 2246
rect 26422 2000 26478 2009
rect 26422 1935 26478 1944
rect 26146 504 26202 513
rect 2778 439 2834 448
rect 3330 0 3386 480
rect 4250 0 4306 480
rect 5262 0 5318 480
rect 6182 0 6238 480
rect 7194 0 7250 480
rect 8114 0 8170 480
rect 9126 0 9182 480
rect 10046 0 10102 480
rect 11058 0 11114 480
rect 11978 0 12034 480
rect 12990 0 13046 480
rect 13910 0 13966 480
rect 14922 0 14978 480
rect 15842 0 15898 480
rect 16854 0 16910 480
rect 17774 0 17830 480
rect 18786 0 18842 480
rect 19706 0 19762 480
rect 20718 0 20774 480
rect 21638 0 21694 480
rect 22650 0 22706 480
rect 23570 0 23626 480
rect 24582 0 24638 480
rect 25502 0 25558 480
rect 26528 480 26556 5743
rect 27434 2816 27490 2825
rect 27434 2751 27490 2760
rect 27448 480 27476 2751
rect 26146 439 26202 448
rect 26514 0 26570 480
rect 27434 0 27490 480
<< via2 >>
rect 1582 27376 1638 27432
rect 24766 27376 24822 27432
rect 1398 25336 1454 25392
rect 1214 23160 1270 23216
rect 386 18264 442 18320
rect 1398 21120 1454 21176
rect 2594 26288 2650 26344
rect 23478 26288 23534 26344
rect 1214 12416 1270 12472
rect 1398 17992 1454 18048
rect 1490 12416 1546 12472
rect 570 9696 626 9752
rect 1674 10920 1730 10976
rect 1582 7656 1638 7712
rect 1582 5616 1638 5672
rect 1582 4528 1638 4584
rect 2134 20868 2190 20904
rect 2134 20848 2136 20868
rect 2136 20848 2188 20868
rect 2188 20848 2190 20868
rect 1858 19352 1914 19408
rect 1950 17740 2006 17776
rect 1950 17720 1952 17740
rect 1952 17720 2004 17740
rect 2004 17720 2006 17740
rect 2134 19236 2190 19272
rect 2134 19216 2136 19236
rect 2136 19216 2188 19236
rect 2188 19216 2190 19236
rect 2134 16496 2190 16552
rect 1950 12688 2006 12744
rect 1950 12552 2006 12608
rect 2318 16088 2374 16144
rect 2318 14456 2374 14512
rect 2134 12416 2190 12472
rect 2226 12280 2282 12336
rect 1858 9968 1914 10024
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 2962 24248 3018 24304
rect 2686 21936 2742 21992
rect 2778 20032 2834 20088
rect 2594 18264 2650 18320
rect 2134 9832 2190 9888
rect 2226 9016 2282 9072
rect 1582 3440 1638 3496
rect 2042 3188 2098 3224
rect 2042 3168 2044 3188
rect 2044 3168 2096 3188
rect 2096 3168 2098 3188
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 23846 25336 23902 25392
rect 13542 23724 13598 23760
rect 13542 23704 13544 23724
rect 13544 23704 13596 23724
rect 13596 23704 13598 23724
rect 23478 23704 23534 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 7102 20848 7158 20904
rect 2962 16904 3018 16960
rect 2686 14456 2742 14512
rect 2686 12416 2742 12472
rect 2778 11192 2834 11248
rect 2778 4664 2834 4720
rect 2686 4528 2742 4584
rect 2594 4120 2650 4176
rect 2962 13912 3018 13968
rect 3330 16768 3386 16824
rect 3054 7112 3110 7168
rect 1582 1400 1638 1456
rect 2778 448 2834 504
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 3882 14864 3938 14920
rect 3882 13232 3938 13288
rect 3514 9580 3570 9616
rect 3514 9560 3516 9580
rect 3516 9560 3568 9580
rect 3568 9560 3570 9580
rect 3514 5616 3570 5672
rect 4342 17040 4398 17096
rect 4250 16088 4306 16144
rect 4250 14492 4252 14512
rect 4252 14492 4304 14512
rect 4304 14492 4306 14512
rect 4250 14456 4306 14492
rect 4066 13776 4122 13832
rect 4158 11228 4160 11248
rect 4160 11228 4212 11248
rect 4212 11228 4214 11248
rect 4158 11192 4214 11228
rect 4066 8744 4122 8800
rect 4434 14864 4490 14920
rect 3974 7248 4030 7304
rect 4158 7148 4160 7168
rect 4160 7148 4212 7168
rect 4212 7148 4214 7168
rect 4158 7112 4214 7148
rect 4066 6160 4122 6216
rect 4250 6568 4306 6624
rect 4066 4936 4122 4992
rect 3882 3168 3938 3224
rect 4342 5208 4398 5264
rect 4250 4664 4306 4720
rect 3882 2488 3938 2544
rect 4802 16496 4858 16552
rect 4802 15816 4858 15872
rect 4618 9968 4674 10024
rect 4802 12280 4858 12336
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5078 17176 5134 17232
rect 5170 15816 5226 15872
rect 5078 13640 5134 13696
rect 4986 10920 5042 10976
rect 4986 10104 5042 10160
rect 4894 7404 4950 7440
rect 4894 7384 4896 7404
rect 4896 7384 4948 7404
rect 4948 7384 4950 7404
rect 4986 6296 5042 6352
rect 4618 5072 4674 5128
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5630 13640 5686 13696
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6090 11600 6146 11656
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5722 6976 5778 7032
rect 5998 6976 6054 7032
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5722 6160 5778 6216
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6366 13912 6422 13968
rect 6274 12688 6330 12744
rect 6366 10784 6422 10840
rect 6366 9968 6422 10024
rect 6274 8356 6330 8392
rect 6274 8336 6276 8356
rect 6276 8336 6328 8356
rect 6328 8336 6330 8356
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5170 3052 5226 3088
rect 5170 3032 5172 3052
rect 5172 3032 5224 3052
rect 5224 3032 5226 3052
rect 4802 2508 4858 2544
rect 4802 2488 4804 2508
rect 4804 2488 4856 2508
rect 4856 2488 4858 2508
rect 4434 1536 4490 1592
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6550 14456 6606 14512
rect 6550 12280 6606 12336
rect 6550 10104 6606 10160
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 7470 18148 7526 18184
rect 7470 18128 7472 18148
rect 7472 18128 7524 18148
rect 7524 18128 7526 18148
rect 7010 12724 7012 12744
rect 7012 12724 7064 12744
rect 7064 12724 7066 12744
rect 7010 12688 7066 12724
rect 7102 9696 7158 9752
rect 6826 9288 6882 9344
rect 6550 5616 6606 5672
rect 6550 4140 6606 4176
rect 6550 4120 6552 4140
rect 6552 4120 6604 4140
rect 6604 4120 6606 4140
rect 6182 3304 6238 3360
rect 6274 3068 6276 3088
rect 6276 3068 6328 3088
rect 6328 3068 6330 3088
rect 6274 3032 6330 3068
rect 7378 12824 7434 12880
rect 7378 7928 7434 7984
rect 7286 7384 7342 7440
rect 7286 5244 7288 5264
rect 7288 5244 7340 5264
rect 7340 5244 7342 5264
rect 7286 5208 7342 5244
rect 6366 2644 6422 2680
rect 6918 3440 6974 3496
rect 7562 15000 7618 15056
rect 7746 13912 7802 13968
rect 8114 13368 8170 13424
rect 8114 13096 8170 13152
rect 8114 12824 8170 12880
rect 7746 10920 7802 10976
rect 7838 9968 7894 10024
rect 7838 9832 7894 9888
rect 7654 9560 7710 9616
rect 7654 9424 7710 9480
rect 7838 9016 7894 9072
rect 7930 8472 7986 8528
rect 8114 11736 8170 11792
rect 8298 15000 8354 15056
rect 8482 16768 8538 16824
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 12162 17720 12218 17776
rect 9034 17060 9090 17096
rect 9034 17040 9036 17060
rect 9036 17040 9088 17060
rect 9088 17040 9090 17060
rect 8666 15680 8722 15736
rect 8574 13912 8630 13968
rect 8758 13640 8814 13696
rect 8666 13504 8722 13560
rect 8574 12588 8576 12608
rect 8576 12588 8628 12608
rect 8628 12588 8630 12608
rect 8574 12552 8630 12588
rect 8114 9424 8170 9480
rect 8666 9696 8722 9752
rect 8206 8608 8262 8664
rect 7378 3596 7434 3632
rect 7378 3576 7380 3596
rect 7380 3576 7432 3596
rect 7432 3576 7434 3596
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6366 2624 6368 2644
rect 6368 2624 6420 2644
rect 6420 2624 6422 2644
rect 8482 6976 8538 7032
rect 8758 6196 8760 6216
rect 8760 6196 8812 6216
rect 8812 6196 8814 6216
rect 8758 6160 8814 6196
rect 8114 5652 8116 5672
rect 8116 5652 8168 5672
rect 8168 5652 8170 5672
rect 8114 5616 8170 5652
rect 8206 3440 8262 3496
rect 8022 2896 8078 2952
rect 9126 16904 9182 16960
rect 9126 15000 9182 15056
rect 9770 13504 9826 13560
rect 9770 13232 9826 13288
rect 9494 9324 9496 9344
rect 9496 9324 9548 9344
rect 9548 9324 9550 9344
rect 9494 9288 9550 9324
rect 9678 8916 9680 8936
rect 9680 8916 9732 8936
rect 9732 8916 9734 8936
rect 9678 8880 9734 8916
rect 9770 8492 9826 8528
rect 9770 8472 9772 8492
rect 9772 8472 9824 8492
rect 9824 8472 9826 8492
rect 9678 5616 9734 5672
rect 8942 2896 8998 2952
rect 8850 1808 8906 1864
rect 9402 3440 9458 3496
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10138 15680 10194 15736
rect 10874 15680 10930 15736
rect 10230 15156 10286 15192
rect 10230 15136 10232 15156
rect 10232 15136 10284 15156
rect 10284 15136 10286 15156
rect 10690 15136 10746 15192
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10230 13404 10232 13424
rect 10232 13404 10284 13424
rect 10284 13404 10286 13424
rect 10230 13368 10286 13404
rect 10046 12824 10102 12880
rect 10874 12860 10876 12880
rect 10876 12860 10928 12880
rect 10928 12860 10930 12880
rect 10874 12824 10930 12860
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10322 11772 10324 11792
rect 10324 11772 10376 11792
rect 10376 11772 10378 11792
rect 10322 11736 10378 11772
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10598 8628 10654 8664
rect 10598 8608 10600 8628
rect 10600 8608 10652 8628
rect 10652 8608 10654 8628
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10874 7792 10930 7848
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10598 4020 10600 4040
rect 10600 4020 10652 4040
rect 10652 4020 10654 4040
rect 10598 3984 10654 4020
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 9586 2624 9642 2680
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10690 2644 10746 2680
rect 9218 2388 9220 2408
rect 9220 2388 9272 2408
rect 9272 2388 9274 2408
rect 9218 2352 9274 2388
rect 10690 2624 10692 2644
rect 10692 2624 10744 2644
rect 10744 2624 10746 2644
rect 11150 11872 11206 11928
rect 11150 10648 11206 10704
rect 11058 10412 11060 10432
rect 11060 10412 11112 10432
rect 11112 10412 11114 10432
rect 11058 10376 11114 10412
rect 11518 9832 11574 9888
rect 11242 8336 11298 8392
rect 12254 14728 12310 14784
rect 12070 12960 12126 13016
rect 11886 12688 11942 12744
rect 12070 12688 12126 12744
rect 11886 11464 11942 11520
rect 11794 10240 11850 10296
rect 11978 9036 12034 9072
rect 11978 9016 11980 9036
rect 11980 9016 12032 9036
rect 12032 9016 12034 9036
rect 12714 15816 12770 15872
rect 12714 15544 12770 15600
rect 12622 10784 12678 10840
rect 12714 10512 12770 10568
rect 12898 7248 12954 7304
rect 12070 6296 12126 6352
rect 11886 5244 11888 5264
rect 11888 5244 11940 5264
rect 11940 5244 11942 5264
rect 11886 5208 11942 5244
rect 11058 3476 11060 3496
rect 11060 3476 11112 3496
rect 11112 3476 11114 3496
rect 11058 3440 11114 3476
rect 11058 3304 11114 3360
rect 10230 1672 10286 1728
rect 11610 3440 11666 3496
rect 12898 4528 12954 4584
rect 12622 3476 12624 3496
rect 12624 3476 12676 3496
rect 12676 3476 12678 3496
rect 12622 3440 12678 3476
rect 13266 12552 13322 12608
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 23570 23160 23626 23216
rect 16486 21528 16542 21584
rect 23478 21528 23534 21584
rect 13450 21412 13506 21448
rect 13450 21392 13452 21412
rect 13452 21392 13504 21412
rect 13504 21392 13506 21412
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14094 19896 14150 19952
rect 14002 18128 14058 18184
rect 13726 15444 13728 15464
rect 13728 15444 13780 15464
rect 13780 15444 13782 15464
rect 13726 15408 13782 15444
rect 13634 15156 13690 15192
rect 13634 15136 13636 15156
rect 13636 15136 13688 15156
rect 13688 15136 13690 15156
rect 13910 13912 13966 13968
rect 13726 13504 13782 13560
rect 13542 12280 13598 12336
rect 13542 11736 13598 11792
rect 13542 9424 13598 9480
rect 13910 10376 13966 10432
rect 13358 7828 13360 7848
rect 13360 7828 13412 7848
rect 13412 7828 13414 7848
rect 13358 7792 13414 7828
rect 13726 7384 13782 7440
rect 13542 6704 13598 6760
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 16210 18672 16266 18728
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14462 14864 14518 14920
rect 14370 12824 14426 12880
rect 14370 11736 14426 11792
rect 14370 9560 14426 9616
rect 14554 11464 14610 11520
rect 14094 9016 14150 9072
rect 14278 9036 14334 9072
rect 14278 9016 14280 9036
rect 14280 9016 14332 9036
rect 14332 9016 14334 9036
rect 14186 6432 14242 6488
rect 14094 6160 14150 6216
rect 13634 5364 13690 5400
rect 13634 5344 13636 5364
rect 13636 5344 13688 5364
rect 13688 5344 13690 5364
rect 13450 3188 13506 3224
rect 13450 3168 13452 3188
rect 13452 3168 13504 3188
rect 13504 3168 13506 3188
rect 13818 3068 13820 3088
rect 13820 3068 13872 3088
rect 13872 3068 13874 3088
rect 13818 3032 13874 3068
rect 13634 2760 13690 2816
rect 13266 2352 13322 2408
rect 14186 5616 14242 5672
rect 14186 5208 14242 5264
rect 14646 10512 14702 10568
rect 14370 5616 14426 5672
rect 14094 5092 14150 5128
rect 14094 5072 14096 5092
rect 14096 5072 14148 5092
rect 14148 5072 14150 5092
rect 14278 5072 14334 5128
rect 14278 4548 14334 4584
rect 14278 4528 14280 4548
rect 14280 4528 14332 4548
rect 14332 4528 14334 4548
rect 14646 5208 14702 5264
rect 14278 3460 14334 3496
rect 14278 3440 14280 3460
rect 14280 3440 14332 3460
rect 14332 3440 14334 3460
rect 14186 2624 14242 2680
rect 14278 2352 14334 2408
rect 14462 1944 14518 2000
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15474 15816 15530 15872
rect 15290 15408 15346 15464
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14830 14320 14886 14376
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14830 13912 14886 13968
rect 15658 15680 15714 15736
rect 15474 14184 15530 14240
rect 15474 13932 15530 13968
rect 15474 13912 15476 13932
rect 15476 13912 15528 13932
rect 15528 13912 15530 13932
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15382 11192 15438 11248
rect 15842 14728 15898 14784
rect 16026 16632 16082 16688
rect 16026 15272 16082 15328
rect 16026 13268 16028 13288
rect 16028 13268 16080 13288
rect 16080 13268 16082 13288
rect 16026 13232 16082 13268
rect 15750 12552 15806 12608
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15382 8880 15438 8936
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15934 12144 15990 12200
rect 15566 8780 15568 8800
rect 15568 8780 15620 8800
rect 15620 8780 15622 8800
rect 15566 8744 15622 8780
rect 15750 7928 15806 7984
rect 15934 9152 15990 9208
rect 15382 5616 15438 5672
rect 15658 5244 15660 5264
rect 15660 5244 15712 5264
rect 15712 5244 15714 5264
rect 15658 5208 15714 5244
rect 15566 4800 15622 4856
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15198 3984 15254 4040
rect 15382 3576 15438 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14922 3032 14978 3088
rect 23570 21392 23626 21448
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 17590 20712 17646 20768
rect 23478 20748 23480 20768
rect 23480 20748 23532 20768
rect 23532 20748 23534 20768
rect 23478 20712 23534 20748
rect 16578 14048 16634 14104
rect 16302 12416 16358 12472
rect 17406 14864 17462 14920
rect 17038 14356 17040 14376
rect 17040 14356 17092 14376
rect 17092 14356 17094 14376
rect 17038 14320 17094 14356
rect 16762 11872 16818 11928
rect 16302 8336 16358 8392
rect 16210 6432 16266 6488
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15750 2252 15752 2272
rect 15752 2252 15804 2272
rect 15804 2252 15806 2272
rect 15750 2216 15806 2252
rect 15290 1536 15346 1592
rect 15934 3596 15990 3632
rect 15934 3576 15936 3596
rect 15936 3576 15988 3596
rect 15988 3576 15990 3596
rect 15934 2760 15990 2816
rect 16946 11500 16948 11520
rect 16948 11500 17000 11520
rect 17000 11500 17002 11520
rect 16946 11464 17002 11500
rect 16762 10512 16818 10568
rect 16946 10412 16948 10432
rect 16948 10412 17000 10432
rect 17000 10412 17002 10432
rect 16946 10376 17002 10412
rect 16578 7384 16634 7440
rect 17314 13640 17370 13696
rect 17314 10648 17370 10704
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 23662 18672 23718 18728
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19522 17176 19578 17232
rect 18050 17040 18106 17096
rect 17774 15580 17776 15600
rect 17776 15580 17828 15600
rect 17828 15580 17830 15600
rect 17774 15544 17830 15580
rect 17958 13912 18014 13968
rect 17314 9968 17370 10024
rect 17130 7268 17186 7304
rect 17130 7248 17132 7268
rect 17132 7248 17184 7268
rect 17184 7248 17186 7268
rect 16946 6996 17002 7032
rect 16946 6976 16948 6996
rect 16948 6976 17000 6996
rect 17000 6976 17002 6996
rect 17866 12824 17922 12880
rect 17958 12416 18014 12472
rect 17774 12316 17776 12336
rect 17776 12316 17828 12336
rect 17828 12316 17830 12336
rect 17774 12280 17830 12316
rect 18142 12552 18198 12608
rect 18142 11756 18198 11792
rect 18326 13096 18382 13152
rect 18326 12416 18382 12472
rect 18142 11736 18144 11756
rect 18144 11736 18196 11756
rect 18196 11736 18198 11756
rect 18050 9152 18106 9208
rect 16854 5652 16856 5672
rect 16856 5652 16908 5672
rect 16908 5652 16910 5672
rect 16854 5616 16910 5652
rect 16578 3032 16634 3088
rect 16302 2488 16358 2544
rect 16026 2352 16082 2408
rect 16762 1808 16818 1864
rect 17590 5908 17646 5944
rect 17590 5888 17592 5908
rect 17592 5888 17644 5908
rect 17644 5888 17646 5908
rect 17958 6432 18014 6488
rect 17958 5072 18014 5128
rect 17590 4684 17646 4720
rect 17590 4664 17592 4684
rect 17592 4664 17644 4684
rect 17644 4664 17646 4684
rect 17774 4120 17830 4176
rect 18510 9016 18566 9072
rect 18878 13524 18934 13560
rect 18878 13504 18880 13524
rect 18880 13504 18932 13524
rect 18932 13504 18934 13524
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20994 16496 21050 16552
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19982 15000 20038 15056
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19154 12416 19210 12472
rect 19338 11192 19394 11248
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 18510 6296 18566 6352
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19338 8744 19394 8800
rect 19982 10124 20038 10160
rect 19982 10104 19984 10124
rect 19984 10104 20036 10124
rect 20036 10104 20038 10124
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19430 6976 19486 7032
rect 19246 6432 19302 6488
rect 19246 6160 19302 6216
rect 19062 5888 19118 5944
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19430 4820 19486 4856
rect 19430 4800 19432 4820
rect 19432 4800 19484 4820
rect 19484 4800 19486 4820
rect 17406 2080 17462 2136
rect 16946 1672 17002 1728
rect 18418 3612 18420 3632
rect 18420 3612 18472 3632
rect 18472 3612 18474 3632
rect 18418 3576 18474 3612
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20626 15272 20682 15328
rect 20350 11620 20406 11656
rect 20350 11600 20352 11620
rect 20352 11600 20404 11620
rect 20404 11600 20406 11620
rect 20626 12416 20682 12472
rect 20902 14184 20958 14240
rect 20810 12724 20812 12744
rect 20812 12724 20864 12744
rect 20864 12724 20866 12744
rect 20810 12688 20866 12724
rect 20258 8356 20314 8392
rect 20258 8336 20260 8356
rect 20260 8336 20312 8356
rect 20312 8336 20314 8356
rect 20718 11736 20774 11792
rect 20810 10512 20866 10568
rect 23478 15544 23534 15600
rect 20902 8064 20958 8120
rect 20994 7420 20996 7440
rect 20996 7420 21048 7440
rect 21048 7420 21050 7440
rect 20994 7384 21050 7420
rect 20718 5108 20720 5128
rect 20720 5108 20772 5128
rect 20772 5108 20774 5128
rect 20718 5072 20774 5108
rect 21454 9696 21510 9752
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24248 24730 24304
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24674 22208 24730 22264
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 21120 24822 21176
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24674 19080 24730 19136
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24214 17992 24270 18048
rect 22006 14476 22062 14512
rect 22006 14456 22008 14476
rect 22008 14456 22060 14476
rect 22060 14456 22062 14476
rect 21730 6452 21786 6488
rect 21730 6432 21732 6452
rect 21732 6432 21784 6452
rect 21784 6432 21786 6452
rect 21178 5752 21234 5808
rect 21454 5636 21510 5672
rect 21454 5616 21456 5636
rect 21456 5616 21508 5636
rect 21508 5616 21510 5636
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 21270 2624 21326 2680
rect 19246 2488 19302 2544
rect 20718 2216 20774 2272
rect 19706 1944 19762 2000
rect 21546 2080 21602 2136
rect 22098 12164 22154 12200
rect 22098 12144 22100 12164
rect 22100 12144 22152 12164
rect 22152 12144 22154 12164
rect 22098 12008 22154 12064
rect 21822 4528 21878 4584
rect 23570 14320 23626 14376
rect 22190 6160 22246 6216
rect 22650 10920 22706 10976
rect 22282 4564 22284 4584
rect 22284 4564 22336 4584
rect 22336 4564 22338 4584
rect 22282 4528 22338 4564
rect 22834 6704 22890 6760
rect 22558 4120 22614 4176
rect 22190 2524 22192 2544
rect 22192 2524 22244 2544
rect 22244 2524 22246 2544
rect 22190 2488 22246 2524
rect 23018 11872 23074 11928
rect 23478 13252 23534 13288
rect 23478 13232 23480 13252
rect 23480 13232 23532 13252
rect 23532 13232 23534 13252
rect 23478 12688 23534 12744
rect 23754 12008 23810 12064
rect 23478 11736 23534 11792
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13912 24822 13968
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 23478 10140 23480 10160
rect 23480 10140 23532 10160
rect 23532 10140 23534 10160
rect 23478 10104 23534 10140
rect 23478 9560 23534 9616
rect 23110 7792 23166 7848
rect 23570 7384 23626 7440
rect 23478 7268 23534 7304
rect 23478 7248 23480 7268
rect 23480 7248 23532 7268
rect 23532 7248 23534 7268
rect 23570 3440 23626 3496
rect 23294 3032 23350 3088
rect 22650 2796 22652 2816
rect 22652 2796 22704 2816
rect 22704 2796 22706 2816
rect 22650 2760 22706 2796
rect 23018 1400 23074 1456
rect 24214 12416 24270 12472
rect 24122 11636 24124 11656
rect 24124 11636 24176 11656
rect 24176 11636 24178 11656
rect 24122 11600 24178 11636
rect 24950 13368 25006 13424
rect 24950 12824 25006 12880
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24306 8880 24362 8936
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 23846 8336 23902 8392
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25042 10784 25098 10840
rect 25226 10512 25282 10568
rect 24766 8744 24822 8800
rect 24674 5616 24730 5672
rect 24950 8880 25006 8936
rect 25226 8064 25282 8120
rect 25502 12280 25558 12336
rect 25410 9696 25466 9752
rect 25410 6568 25466 6624
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24674 3032 24730 3088
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23662 1944 23718 2000
rect 25410 4528 25466 4584
rect 25686 9968 25742 10024
rect 25594 8336 25650 8392
rect 25502 3984 25558 4040
rect 25410 3440 25466 3496
rect 25410 2644 25466 2680
rect 25410 2624 25412 2644
rect 25412 2624 25464 2644
rect 25464 2624 25466 2644
rect 24766 2488 24822 2544
rect 24858 2372 24914 2408
rect 24858 2352 24860 2372
rect 24860 2352 24912 2372
rect 24912 2352 24914 2372
rect 26514 5752 26570 5808
rect 26422 1944 26478 2000
rect 26146 448 26202 504
rect 27434 2760 27490 2816
<< metal3 >>
rect 0 27434 480 27464
rect 1577 27434 1643 27437
rect 0 27432 1643 27434
rect 0 27376 1582 27432
rect 1638 27376 1643 27432
rect 0 27374 1643 27376
rect 0 27344 480 27374
rect 1577 27371 1643 27374
rect 24761 27434 24827 27437
rect 27520 27434 28000 27464
rect 24761 27432 28000 27434
rect 24761 27376 24766 27432
rect 24822 27376 28000 27432
rect 24761 27374 28000 27376
rect 24761 27371 24827 27374
rect 27520 27344 28000 27374
rect 0 26346 480 26376
rect 2589 26346 2655 26349
rect 0 26344 2655 26346
rect 0 26288 2594 26344
rect 2650 26288 2655 26344
rect 0 26286 2655 26288
rect 0 26256 480 26286
rect 2589 26283 2655 26286
rect 23473 26346 23539 26349
rect 27520 26346 28000 26376
rect 23473 26344 28000 26346
rect 23473 26288 23478 26344
rect 23534 26288 28000 26344
rect 23473 26286 28000 26288
rect 23473 26283 23539 26286
rect 27520 26256 28000 26286
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 1393 25394 1459 25397
rect 0 25392 1459 25394
rect 0 25336 1398 25392
rect 1454 25336 1459 25392
rect 0 25334 1459 25336
rect 0 25304 480 25334
rect 1393 25331 1459 25334
rect 23841 25394 23907 25397
rect 27520 25394 28000 25424
rect 23841 25392 28000 25394
rect 23841 25336 23846 25392
rect 23902 25336 28000 25392
rect 23841 25334 28000 25336
rect 23841 25331 23907 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24306 480 24336
rect 2957 24306 3023 24309
rect 0 24304 3023 24306
rect 0 24248 2962 24304
rect 3018 24248 3023 24304
rect 0 24246 3023 24248
rect 0 24216 480 24246
rect 2957 24243 3023 24246
rect 24669 24306 24735 24309
rect 27520 24306 28000 24336
rect 24669 24304 28000 24306
rect 24669 24248 24674 24304
rect 24730 24248 28000 24304
rect 24669 24246 28000 24248
rect 24669 24243 24735 24246
rect 27520 24216 28000 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 13537 23762 13603 23765
rect 23473 23762 23539 23765
rect 13537 23760 23539 23762
rect 13537 23704 13542 23760
rect 13598 23704 23478 23760
rect 23534 23704 23539 23760
rect 13537 23702 23539 23704
rect 13537 23699 13603 23702
rect 23473 23699 23539 23702
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23218 480 23248
rect 1209 23218 1275 23221
rect 0 23216 1275 23218
rect 0 23160 1214 23216
rect 1270 23160 1275 23216
rect 0 23158 1275 23160
rect 0 23128 480 23158
rect 1209 23155 1275 23158
rect 23565 23218 23631 23221
rect 27520 23218 28000 23248
rect 23565 23216 28000 23218
rect 23565 23160 23570 23216
rect 23626 23160 28000 23216
rect 23565 23158 28000 23160
rect 23565 23155 23631 23158
rect 27520 23128 28000 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 24669 22266 24735 22269
rect 27520 22266 28000 22296
rect 0 22206 2146 22266
rect 0 22176 480 22206
rect 2086 21994 2146 22206
rect 24669 22264 28000 22266
rect 24669 22208 24674 22264
rect 24730 22208 28000 22264
rect 24669 22206 28000 22208
rect 24669 22203 24735 22206
rect 27520 22176 28000 22206
rect 2681 21994 2747 21997
rect 2086 21992 2747 21994
rect 2086 21936 2686 21992
rect 2742 21936 2747 21992
rect 2086 21934 2747 21936
rect 2681 21931 2747 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 16481 21586 16547 21589
rect 23473 21586 23539 21589
rect 16481 21584 23539 21586
rect 16481 21528 16486 21584
rect 16542 21528 23478 21584
rect 23534 21528 23539 21584
rect 16481 21526 23539 21528
rect 16481 21523 16547 21526
rect 23473 21523 23539 21526
rect 13445 21450 13511 21453
rect 23565 21450 23631 21453
rect 13445 21448 23631 21450
rect 13445 21392 13450 21448
rect 13506 21392 23570 21448
rect 23626 21392 23631 21448
rect 13445 21390 23631 21392
rect 13445 21387 13511 21390
rect 23565 21387 23631 21390
rect 10277 21248 10597 21249
rect 0 21178 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 480 21118
rect 1393 21115 1459 21118
rect 24761 21178 24827 21181
rect 27520 21178 28000 21208
rect 24761 21176 28000 21178
rect 24761 21120 24766 21176
rect 24822 21120 28000 21176
rect 24761 21118 28000 21120
rect 24761 21115 24827 21118
rect 27520 21088 28000 21118
rect 2129 20906 2195 20909
rect 7097 20906 7163 20909
rect 2129 20904 7163 20906
rect 2129 20848 2134 20904
rect 2190 20848 7102 20904
rect 7158 20848 7163 20904
rect 2129 20846 7163 20848
rect 2129 20843 2195 20846
rect 7097 20843 7163 20846
rect 17585 20770 17651 20773
rect 23473 20770 23539 20773
rect 17585 20768 23539 20770
rect 17585 20712 17590 20768
rect 17646 20712 23478 20768
rect 23534 20712 23539 20768
rect 17585 20710 23539 20712
rect 17585 20707 17651 20710
rect 23473 20707 23539 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 2773 20090 2839 20093
rect 27520 20090 28000 20120
rect 0 20088 2839 20090
rect 0 20032 2778 20088
rect 2834 20032 2839 20088
rect 0 20030 2839 20032
rect 0 20000 480 20030
rect 2773 20027 2839 20030
rect 24902 20030 28000 20090
rect 14089 19954 14155 19957
rect 24902 19954 24962 20030
rect 27520 20000 28000 20030
rect 14089 19952 24962 19954
rect 14089 19896 14094 19952
rect 14150 19896 24962 19952
rect 14089 19894 24962 19896
rect 14089 19891 14155 19894
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 1853 19410 1919 19413
rect 1534 19408 1919 19410
rect 1534 19352 1858 19408
rect 1914 19352 1919 19408
rect 1534 19350 1919 19352
rect 0 19138 480 19168
rect 1534 19138 1594 19350
rect 1853 19347 1919 19350
rect 2129 19274 2195 19277
rect 9806 19274 9812 19276
rect 2129 19272 9812 19274
rect 2129 19216 2134 19272
rect 2190 19216 9812 19272
rect 2129 19214 9812 19216
rect 2129 19211 2195 19214
rect 9806 19212 9812 19214
rect 9876 19212 9882 19276
rect 0 19078 1594 19138
rect 24669 19138 24735 19141
rect 27520 19138 28000 19168
rect 24669 19136 28000 19138
rect 24669 19080 24674 19136
rect 24730 19080 28000 19136
rect 24669 19078 28000 19080
rect 0 19048 480 19078
rect 24669 19075 24735 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 16205 18730 16271 18733
rect 23657 18730 23723 18733
rect 16205 18728 23723 18730
rect 16205 18672 16210 18728
rect 16266 18672 23662 18728
rect 23718 18672 23723 18728
rect 16205 18670 23723 18672
rect 16205 18667 16271 18670
rect 23657 18667 23723 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 381 18322 447 18325
rect 2589 18322 2655 18325
rect 381 18320 2655 18322
rect 381 18264 386 18320
rect 442 18264 2594 18320
rect 2650 18264 2655 18320
rect 381 18262 2655 18264
rect 381 18259 447 18262
rect 2589 18259 2655 18262
rect 7465 18186 7531 18189
rect 13997 18186 14063 18189
rect 7465 18184 14063 18186
rect 7465 18128 7470 18184
rect 7526 18128 14002 18184
rect 14058 18128 14063 18184
rect 7465 18126 14063 18128
rect 7465 18123 7531 18126
rect 13997 18123 14063 18126
rect 0 18050 480 18080
rect 1393 18050 1459 18053
rect 0 18048 1459 18050
rect 0 17992 1398 18048
rect 1454 17992 1459 18048
rect 0 17990 1459 17992
rect 0 17960 480 17990
rect 1393 17987 1459 17990
rect 24209 18050 24275 18053
rect 27520 18050 28000 18080
rect 24209 18048 28000 18050
rect 24209 17992 24214 18048
rect 24270 17992 28000 18048
rect 24209 17990 28000 17992
rect 24209 17987 24275 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 1945 17778 2011 17781
rect 12157 17778 12223 17781
rect 1945 17776 12223 17778
rect 1945 17720 1950 17776
rect 2006 17720 12162 17776
rect 12218 17720 12223 17776
rect 1945 17718 12223 17720
rect 1945 17715 2011 17718
rect 12157 17715 12223 17718
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 5073 17234 5139 17237
rect 19517 17234 19583 17237
rect 5073 17232 24962 17234
rect 5073 17176 5078 17232
rect 5134 17176 19522 17232
rect 19578 17176 24962 17232
rect 5073 17174 24962 17176
rect 5073 17171 5139 17174
rect 19517 17171 19583 17174
rect 0 17098 480 17128
rect 4337 17098 4403 17101
rect 4470 17098 4476 17100
rect 0 17038 2882 17098
rect 0 17008 480 17038
rect 2822 16690 2882 17038
rect 4337 17096 4476 17098
rect 4337 17040 4342 17096
rect 4398 17040 4476 17096
rect 4337 17038 4476 17040
rect 4337 17035 4403 17038
rect 4470 17036 4476 17038
rect 4540 17036 4546 17100
rect 9029 17098 9095 17101
rect 18045 17098 18111 17101
rect 9029 17096 18111 17098
rect 9029 17040 9034 17096
rect 9090 17040 18050 17096
rect 18106 17040 18111 17096
rect 9029 17038 18111 17040
rect 24902 17098 24962 17174
rect 27520 17098 28000 17128
rect 24902 17038 28000 17098
rect 9029 17035 9095 17038
rect 18045 17035 18111 17038
rect 27520 17008 28000 17038
rect 2957 16962 3023 16965
rect 9121 16962 9187 16965
rect 2957 16960 9187 16962
rect 2957 16904 2962 16960
rect 3018 16904 9126 16960
rect 9182 16904 9187 16960
rect 2957 16902 9187 16904
rect 2957 16899 3023 16902
rect 9121 16899 9187 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 3325 16826 3391 16829
rect 8477 16826 8543 16829
rect 3325 16824 8543 16826
rect 3325 16768 3330 16824
rect 3386 16768 8482 16824
rect 8538 16768 8543 16824
rect 3325 16766 8543 16768
rect 3325 16763 3391 16766
rect 8477 16763 8543 16766
rect 16021 16690 16087 16693
rect 2822 16688 16087 16690
rect 2822 16632 16026 16688
rect 16082 16632 16087 16688
rect 2822 16630 16087 16632
rect 16021 16627 16087 16630
rect 2129 16554 2195 16557
rect 4797 16554 4863 16557
rect 20989 16554 21055 16557
rect 2129 16552 24962 16554
rect 2129 16496 2134 16552
rect 2190 16496 4802 16552
rect 4858 16496 20994 16552
rect 21050 16496 24962 16552
rect 2129 16494 24962 16496
rect 2129 16491 2195 16494
rect 4797 16491 4863 16494
rect 20989 16491 21055 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 2313 16146 2379 16149
rect 4245 16146 4311 16149
rect 2313 16144 4311 16146
rect 2313 16088 2318 16144
rect 2374 16088 4250 16144
rect 4306 16088 4311 16144
rect 2313 16086 4311 16088
rect 2313 16083 2379 16086
rect 4245 16083 4311 16086
rect 0 16010 480 16040
rect 24902 16010 24962 16494
rect 27520 16010 28000 16040
rect 0 15950 7666 16010
rect 24902 15950 28000 16010
rect 0 15920 480 15950
rect 4797 15874 4863 15877
rect 5165 15874 5231 15877
rect 4797 15872 5231 15874
rect 4797 15816 4802 15872
rect 4858 15816 5170 15872
rect 5226 15816 5231 15872
rect 4797 15814 5231 15816
rect 4797 15811 4863 15814
rect 5165 15811 5231 15814
rect 7606 15602 7666 15950
rect 27520 15920 28000 15950
rect 12709 15874 12775 15877
rect 15469 15874 15535 15877
rect 12709 15872 15535 15874
rect 12709 15816 12714 15872
rect 12770 15816 15474 15872
rect 15530 15816 15535 15872
rect 12709 15814 15535 15816
rect 12709 15811 12775 15814
rect 15469 15811 15535 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 8661 15738 8727 15741
rect 10133 15738 10199 15741
rect 8661 15736 10199 15738
rect 8661 15680 8666 15736
rect 8722 15680 10138 15736
rect 10194 15680 10199 15736
rect 8661 15678 10199 15680
rect 8661 15675 8727 15678
rect 10133 15675 10199 15678
rect 10869 15738 10935 15741
rect 15653 15738 15719 15741
rect 10869 15736 15719 15738
rect 10869 15680 10874 15736
rect 10930 15680 15658 15736
rect 15714 15680 15719 15736
rect 10869 15678 15719 15680
rect 10869 15675 10935 15678
rect 15653 15675 15719 15678
rect 12709 15602 12775 15605
rect 7606 15600 12775 15602
rect 7606 15544 12714 15600
rect 12770 15544 12775 15600
rect 7606 15542 12775 15544
rect 12709 15539 12775 15542
rect 17769 15602 17835 15605
rect 23473 15602 23539 15605
rect 17769 15600 23539 15602
rect 17769 15544 17774 15600
rect 17830 15544 23478 15600
rect 23534 15544 23539 15600
rect 17769 15542 23539 15544
rect 17769 15539 17835 15542
rect 23473 15539 23539 15542
rect 13721 15466 13787 15469
rect 15285 15466 15351 15469
rect 13721 15464 15351 15466
rect 13721 15408 13726 15464
rect 13782 15408 15290 15464
rect 15346 15408 15351 15464
rect 13721 15406 15351 15408
rect 13721 15403 13787 15406
rect 15285 15403 15351 15406
rect 16021 15330 16087 15333
rect 20621 15330 20687 15333
rect 16021 15328 20687 15330
rect 16021 15272 16026 15328
rect 16082 15272 20626 15328
rect 20682 15272 20687 15328
rect 16021 15270 20687 15272
rect 16021 15267 16087 15270
rect 20621 15267 20687 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10225 15194 10291 15197
rect 10685 15194 10751 15197
rect 13629 15194 13695 15197
rect 10225 15192 13695 15194
rect 10225 15136 10230 15192
rect 10286 15136 10690 15192
rect 10746 15136 13634 15192
rect 13690 15136 13695 15192
rect 10225 15134 13695 15136
rect 10225 15131 10291 15134
rect 10685 15131 10751 15134
rect 13629 15131 13695 15134
rect 7557 15058 7623 15061
rect 8293 15058 8359 15061
rect 9121 15058 9187 15061
rect 19977 15058 20043 15061
rect 7557 15056 8359 15058
rect 7557 15000 7562 15056
rect 7618 15000 8298 15056
rect 8354 15000 8359 15056
rect 7557 14998 8359 15000
rect 7557 14995 7623 14998
rect 8293 14995 8359 14998
rect 8480 15056 20043 15058
rect 8480 15000 9126 15056
rect 9182 15000 19982 15056
rect 20038 15000 20043 15056
rect 8480 14998 20043 15000
rect 0 14922 480 14952
rect 3877 14922 3943 14925
rect 4429 14922 4495 14925
rect 0 14862 3802 14922
rect 0 14832 480 14862
rect 3742 14786 3802 14862
rect 3877 14920 4495 14922
rect 3877 14864 3882 14920
rect 3938 14864 4434 14920
rect 4490 14864 4495 14920
rect 3877 14862 4495 14864
rect 3877 14859 3943 14862
rect 4429 14859 4495 14862
rect 8480 14786 8540 14998
rect 9121 14995 9187 14998
rect 19977 14995 20043 14998
rect 14457 14922 14523 14925
rect 17401 14922 17467 14925
rect 27520 14922 28000 14952
rect 14457 14920 17467 14922
rect 14457 14864 14462 14920
rect 14518 14864 17406 14920
rect 17462 14864 17467 14920
rect 14457 14862 17467 14864
rect 14457 14859 14523 14862
rect 17401 14859 17467 14862
rect 24902 14862 28000 14922
rect 3742 14726 8540 14786
rect 12249 14786 12315 14789
rect 15837 14786 15903 14789
rect 12249 14784 15903 14786
rect 12249 14728 12254 14784
rect 12310 14728 15842 14784
rect 15898 14728 15903 14784
rect 12249 14726 15903 14728
rect 12249 14723 12315 14726
rect 15837 14723 15903 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 2313 14514 2379 14517
rect 2681 14514 2747 14517
rect 4245 14514 4311 14517
rect 2313 14512 4311 14514
rect 2313 14456 2318 14512
rect 2374 14456 2686 14512
rect 2742 14456 4250 14512
rect 4306 14456 4311 14512
rect 2313 14454 4311 14456
rect 2313 14451 2379 14454
rect 2681 14451 2747 14454
rect 4245 14451 4311 14454
rect 6545 14514 6611 14517
rect 22001 14514 22067 14517
rect 24902 14514 24962 14862
rect 27520 14832 28000 14862
rect 6545 14512 24962 14514
rect 6545 14456 6550 14512
rect 6606 14456 22006 14512
rect 22062 14456 24962 14512
rect 6545 14454 24962 14456
rect 6545 14451 6611 14454
rect 22001 14451 22067 14454
rect 14825 14378 14891 14381
rect 17033 14378 17099 14381
rect 23565 14378 23631 14381
rect 14825 14376 23631 14378
rect 14825 14320 14830 14376
rect 14886 14320 17038 14376
rect 17094 14320 23570 14376
rect 23626 14320 23631 14376
rect 14825 14318 23631 14320
rect 14825 14315 14891 14318
rect 17033 14315 17099 14318
rect 23565 14315 23631 14318
rect 15469 14242 15535 14245
rect 20897 14242 20963 14245
rect 15469 14240 20963 14242
rect 15469 14184 15474 14240
rect 15530 14184 20902 14240
rect 20958 14184 20963 14240
rect 15469 14182 20963 14184
rect 15469 14179 15535 14182
rect 20897 14179 20963 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 16573 14106 16639 14109
rect 15334 14104 16639 14106
rect 15334 14048 16578 14104
rect 16634 14048 16639 14104
rect 15334 14046 16639 14048
rect 0 13970 480 14000
rect 2957 13970 3023 13973
rect 0 13968 3023 13970
rect 0 13912 2962 13968
rect 3018 13912 3023 13968
rect 0 13910 3023 13912
rect 0 13880 480 13910
rect 2957 13907 3023 13910
rect 6361 13970 6427 13973
rect 7741 13970 7807 13973
rect 8569 13970 8635 13973
rect 6361 13968 8635 13970
rect 6361 13912 6366 13968
rect 6422 13912 7746 13968
rect 7802 13912 8574 13968
rect 8630 13912 8635 13968
rect 6361 13910 8635 13912
rect 6361 13907 6427 13910
rect 7741 13907 7807 13910
rect 8569 13907 8635 13910
rect 13905 13970 13971 13973
rect 14825 13970 14891 13973
rect 15334 13970 15394 14046
rect 16573 14043 16639 14046
rect 13905 13968 15394 13970
rect 13905 13912 13910 13968
rect 13966 13912 14830 13968
rect 14886 13912 15394 13968
rect 13905 13910 15394 13912
rect 15469 13970 15535 13973
rect 17953 13970 18019 13973
rect 15469 13968 18019 13970
rect 15469 13912 15474 13968
rect 15530 13912 17958 13968
rect 18014 13912 18019 13968
rect 15469 13910 18019 13912
rect 13905 13907 13971 13910
rect 14825 13907 14891 13910
rect 15469 13907 15535 13910
rect 17953 13907 18019 13910
rect 24761 13970 24827 13973
rect 27520 13970 28000 14000
rect 24761 13968 28000 13970
rect 24761 13912 24766 13968
rect 24822 13912 28000 13968
rect 24761 13910 28000 13912
rect 24761 13907 24827 13910
rect 27520 13880 28000 13910
rect 4061 13834 4127 13837
rect 4061 13832 15026 13834
rect 4061 13776 4066 13832
rect 4122 13776 15026 13832
rect 4061 13774 15026 13776
rect 4061 13771 4127 13774
rect 5073 13698 5139 13701
rect 5625 13698 5691 13701
rect 8753 13698 8819 13701
rect 5073 13696 8819 13698
rect 5073 13640 5078 13696
rect 5134 13640 5630 13696
rect 5686 13640 8758 13696
rect 8814 13640 8819 13696
rect 5073 13638 8819 13640
rect 14966 13698 15026 13774
rect 17309 13698 17375 13701
rect 14966 13696 17375 13698
rect 14966 13640 17314 13696
rect 17370 13640 17375 13696
rect 14966 13638 17375 13640
rect 5073 13635 5139 13638
rect 5625 13635 5691 13638
rect 8753 13635 8819 13638
rect 17309 13635 17375 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 8661 13562 8727 13565
rect 9765 13562 9831 13565
rect 8661 13560 9831 13562
rect 8661 13504 8666 13560
rect 8722 13504 9770 13560
rect 9826 13504 9831 13560
rect 8661 13502 9831 13504
rect 8661 13499 8727 13502
rect 9765 13499 9831 13502
rect 13721 13562 13787 13565
rect 18873 13562 18939 13565
rect 13721 13560 18939 13562
rect 13721 13504 13726 13560
rect 13782 13504 18878 13560
rect 18934 13504 18939 13560
rect 13721 13502 18939 13504
rect 13721 13499 13787 13502
rect 18873 13499 18939 13502
rect 8109 13426 8175 13429
rect 10225 13426 10291 13429
rect 24945 13426 25011 13429
rect 8109 13424 10291 13426
rect 8109 13368 8114 13424
rect 8170 13368 10230 13424
rect 10286 13368 10291 13424
rect 8109 13366 10291 13368
rect 8109 13363 8175 13366
rect 10225 13363 10291 13366
rect 10366 13424 25011 13426
rect 10366 13368 24950 13424
rect 25006 13368 25011 13424
rect 10366 13366 25011 13368
rect 3877 13290 3943 13293
rect 9765 13290 9831 13293
rect 10366 13290 10426 13366
rect 24945 13363 25011 13366
rect 16021 13290 16087 13293
rect 23473 13290 23539 13293
rect 3877 13288 6194 13290
rect 3877 13232 3882 13288
rect 3938 13232 6194 13288
rect 3877 13230 6194 13232
rect 3877 13227 3943 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 6134 13018 6194 13230
rect 9765 13288 10426 13290
rect 9765 13232 9770 13288
rect 9826 13232 10426 13288
rect 9765 13230 10426 13232
rect 14782 13230 15946 13290
rect 9765 13227 9831 13230
rect 8109 13154 8175 13157
rect 14782 13154 14842 13230
rect 8109 13152 14842 13154
rect 8109 13096 8114 13152
rect 8170 13096 14842 13152
rect 8109 13094 14842 13096
rect 15886 13154 15946 13230
rect 16021 13288 23539 13290
rect 16021 13232 16026 13288
rect 16082 13232 23478 13288
rect 23534 13232 23539 13288
rect 16021 13230 23539 13232
rect 16021 13227 16087 13230
rect 23473 13227 23539 13230
rect 18321 13154 18387 13157
rect 15886 13152 18387 13154
rect 15886 13096 18326 13152
rect 18382 13096 18387 13152
rect 15886 13094 18387 13096
rect 8109 13091 8175 13094
rect 18321 13091 18387 13094
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 12065 13018 12131 13021
rect 6134 13016 12131 13018
rect 6134 12960 12070 13016
rect 12126 12960 12131 13016
rect 6134 12958 12131 12960
rect 12065 12955 12131 12958
rect 0 12882 480 12912
rect 7373 12882 7439 12885
rect 8109 12882 8175 12885
rect 0 12880 8175 12882
rect 0 12824 7378 12880
rect 7434 12824 8114 12880
rect 8170 12824 8175 12880
rect 0 12822 8175 12824
rect 0 12792 480 12822
rect 7373 12819 7439 12822
rect 8109 12819 8175 12822
rect 9806 12820 9812 12884
rect 9876 12882 9882 12884
rect 10041 12882 10107 12885
rect 9876 12880 10107 12882
rect 9876 12824 10046 12880
rect 10102 12824 10107 12880
rect 9876 12822 10107 12824
rect 9876 12820 9882 12822
rect 10041 12819 10107 12822
rect 10869 12882 10935 12885
rect 14365 12882 14431 12885
rect 17861 12882 17927 12885
rect 10869 12880 17927 12882
rect 10869 12824 10874 12880
rect 10930 12824 14370 12880
rect 14426 12824 17866 12880
rect 17922 12824 17927 12880
rect 10869 12822 17927 12824
rect 10869 12819 10935 12822
rect 14365 12819 14431 12822
rect 17861 12819 17927 12822
rect 24945 12882 25011 12885
rect 27520 12882 28000 12912
rect 24945 12880 28000 12882
rect 24945 12824 24950 12880
rect 25006 12824 28000 12880
rect 24945 12822 28000 12824
rect 24945 12819 25011 12822
rect 27520 12792 28000 12822
rect 1945 12746 2011 12749
rect 6269 12746 6335 12749
rect 1945 12744 6335 12746
rect 1945 12688 1950 12744
rect 2006 12688 6274 12744
rect 6330 12688 6335 12744
rect 1945 12686 6335 12688
rect 1945 12683 2011 12686
rect 6269 12683 6335 12686
rect 7005 12746 7071 12749
rect 11881 12746 11947 12749
rect 7005 12744 11947 12746
rect 7005 12688 7010 12744
rect 7066 12688 11886 12744
rect 11942 12688 11947 12744
rect 7005 12686 11947 12688
rect 7005 12683 7071 12686
rect 11881 12683 11947 12686
rect 12065 12746 12131 12749
rect 20805 12746 20871 12749
rect 23473 12746 23539 12749
rect 12065 12744 23539 12746
rect 12065 12688 12070 12744
rect 12126 12688 20810 12744
rect 20866 12688 23478 12744
rect 23534 12688 23539 12744
rect 12065 12686 23539 12688
rect 12065 12683 12131 12686
rect 20805 12683 20871 12686
rect 23473 12683 23539 12686
rect 1945 12610 2011 12613
rect 8569 12610 8635 12613
rect 1945 12608 8635 12610
rect 1945 12552 1950 12608
rect 2006 12552 8574 12608
rect 8630 12552 8635 12608
rect 1945 12550 8635 12552
rect 1945 12547 2011 12550
rect 8569 12547 8635 12550
rect 13261 12610 13327 12613
rect 15745 12610 15811 12613
rect 18137 12610 18203 12613
rect 13261 12608 18203 12610
rect 13261 12552 13266 12608
rect 13322 12552 15750 12608
rect 15806 12552 18142 12608
rect 18198 12552 18203 12608
rect 13261 12550 18203 12552
rect 13261 12547 13327 12550
rect 15745 12547 15811 12550
rect 18137 12547 18203 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 1209 12474 1275 12477
rect 1485 12474 1551 12477
rect 1209 12472 1551 12474
rect 1209 12416 1214 12472
rect 1270 12416 1490 12472
rect 1546 12416 1551 12472
rect 1209 12414 1551 12416
rect 1209 12411 1275 12414
rect 1485 12411 1551 12414
rect 2129 12474 2195 12477
rect 2681 12474 2747 12477
rect 2129 12472 2747 12474
rect 2129 12416 2134 12472
rect 2190 12416 2686 12472
rect 2742 12416 2747 12472
rect 2129 12414 2747 12416
rect 2129 12411 2195 12414
rect 2681 12411 2747 12414
rect 16297 12474 16363 12477
rect 17953 12474 18019 12477
rect 16297 12472 18019 12474
rect 16297 12416 16302 12472
rect 16358 12416 17958 12472
rect 18014 12416 18019 12472
rect 16297 12414 18019 12416
rect 16297 12411 16363 12414
rect 17953 12411 18019 12414
rect 18321 12474 18387 12477
rect 19149 12474 19215 12477
rect 20621 12474 20687 12477
rect 24209 12474 24275 12477
rect 18321 12472 19442 12474
rect 18321 12416 18326 12472
rect 18382 12416 19154 12472
rect 19210 12416 19442 12472
rect 18321 12414 19442 12416
rect 18321 12411 18387 12414
rect 19149 12411 19215 12414
rect 2221 12338 2287 12341
rect 4797 12338 4863 12341
rect 6545 12338 6611 12341
rect 2221 12336 6611 12338
rect 2221 12280 2226 12336
rect 2282 12280 4802 12336
rect 4858 12280 6550 12336
rect 6606 12280 6611 12336
rect 2221 12278 6611 12280
rect 2221 12275 2287 12278
rect 4797 12275 4863 12278
rect 6545 12275 6611 12278
rect 13537 12338 13603 12341
rect 17769 12338 17835 12341
rect 13537 12336 17835 12338
rect 13537 12280 13542 12336
rect 13598 12280 17774 12336
rect 17830 12280 17835 12336
rect 13537 12278 17835 12280
rect 19382 12338 19442 12414
rect 20621 12472 24275 12474
rect 20621 12416 20626 12472
rect 20682 12416 24214 12472
rect 24270 12416 24275 12472
rect 20621 12414 24275 12416
rect 20621 12411 20687 12414
rect 24209 12411 24275 12414
rect 25497 12338 25563 12341
rect 19382 12336 25563 12338
rect 19382 12280 25502 12336
rect 25558 12280 25563 12336
rect 19382 12278 25563 12280
rect 13537 12275 13603 12278
rect 17769 12275 17835 12278
rect 25497 12275 25563 12278
rect 15929 12202 15995 12205
rect 22093 12202 22159 12205
rect 15929 12200 22159 12202
rect 15929 12144 15934 12200
rect 15990 12144 22098 12200
rect 22154 12144 22159 12200
rect 15929 12142 22159 12144
rect 15929 12139 15995 12142
rect 22093 12139 22159 12142
rect 22093 12066 22159 12069
rect 23749 12066 23815 12069
rect 22093 12064 23815 12066
rect 22093 12008 22098 12064
rect 22154 12008 23754 12064
rect 23810 12008 23815 12064
rect 22093 12006 23815 12008
rect 22093 12003 22159 12006
rect 23749 12003 23815 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 11145 11930 11211 11933
rect 16757 11930 16823 11933
rect 23013 11930 23079 11933
rect 7974 11928 11211 11930
rect 7974 11872 11150 11928
rect 11206 11872 11211 11928
rect 7974 11870 11211 11872
rect 0 11794 480 11824
rect 7974 11794 8034 11870
rect 11145 11867 11211 11870
rect 15334 11928 23079 11930
rect 15334 11872 16762 11928
rect 16818 11872 23018 11928
rect 23074 11872 23079 11928
rect 15334 11870 23079 11872
rect 0 11734 8034 11794
rect 8109 11794 8175 11797
rect 10317 11794 10383 11797
rect 13537 11794 13603 11797
rect 8109 11792 13603 11794
rect 8109 11736 8114 11792
rect 8170 11736 10322 11792
rect 10378 11736 13542 11792
rect 13598 11736 13603 11792
rect 8109 11734 13603 11736
rect 0 11704 480 11734
rect 8109 11731 8175 11734
rect 10317 11731 10383 11734
rect 13537 11731 13603 11734
rect 14365 11794 14431 11797
rect 15334 11794 15394 11870
rect 16757 11867 16823 11870
rect 23013 11867 23079 11870
rect 14365 11792 15394 11794
rect 14365 11736 14370 11792
rect 14426 11736 15394 11792
rect 14365 11734 15394 11736
rect 18137 11794 18203 11797
rect 20713 11794 20779 11797
rect 18137 11792 20779 11794
rect 18137 11736 18142 11792
rect 18198 11736 20718 11792
rect 20774 11736 20779 11792
rect 18137 11734 20779 11736
rect 14365 11731 14431 11734
rect 18137 11731 18203 11734
rect 20713 11731 20779 11734
rect 23473 11794 23539 11797
rect 27520 11794 28000 11824
rect 23473 11792 28000 11794
rect 23473 11736 23478 11792
rect 23534 11736 28000 11792
rect 23473 11734 28000 11736
rect 23473 11731 23539 11734
rect 27520 11704 28000 11734
rect 4470 11596 4476 11660
rect 4540 11658 4546 11660
rect 6085 11658 6151 11661
rect 4540 11656 6151 11658
rect 4540 11600 6090 11656
rect 6146 11600 6151 11656
rect 4540 11598 6151 11600
rect 4540 11596 4546 11598
rect 6085 11595 6151 11598
rect 20345 11658 20411 11661
rect 24117 11658 24183 11661
rect 20345 11656 24183 11658
rect 20345 11600 20350 11656
rect 20406 11600 24122 11656
rect 24178 11600 24183 11656
rect 20345 11598 24183 11600
rect 20345 11595 20411 11598
rect 24117 11595 24183 11598
rect 11881 11522 11947 11525
rect 14549 11522 14615 11525
rect 16941 11522 17007 11525
rect 11881 11520 17007 11522
rect 11881 11464 11886 11520
rect 11942 11464 14554 11520
rect 14610 11464 16946 11520
rect 17002 11464 17007 11520
rect 11881 11462 17007 11464
rect 11881 11459 11947 11462
rect 14549 11459 14615 11462
rect 16941 11459 17007 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2773 11250 2839 11253
rect 4153 11250 4219 11253
rect 2773 11248 4219 11250
rect 2773 11192 2778 11248
rect 2834 11192 4158 11248
rect 4214 11192 4219 11248
rect 2773 11190 4219 11192
rect 2773 11187 2839 11190
rect 4153 11187 4219 11190
rect 15377 11250 15443 11253
rect 19333 11250 19399 11253
rect 15377 11248 19399 11250
rect 15377 11192 15382 11248
rect 15438 11192 19338 11248
rect 19394 11192 19399 11248
rect 15377 11190 19399 11192
rect 15377 11187 15443 11190
rect 19333 11187 19399 11190
rect 14782 11054 15394 11114
rect 1669 10978 1735 10981
rect 4981 10978 5047 10981
rect 1669 10976 5047 10978
rect 1669 10920 1674 10976
rect 1730 10920 4986 10976
rect 5042 10920 5047 10976
rect 1669 10918 5047 10920
rect 1669 10915 1735 10918
rect 4981 10915 5047 10918
rect 7741 10978 7807 10981
rect 14782 10978 14842 11054
rect 7741 10976 14842 10978
rect 7741 10920 7746 10976
rect 7802 10920 14842 10976
rect 7741 10918 14842 10920
rect 15334 10978 15394 11054
rect 22645 10978 22711 10981
rect 15334 10976 22711 10978
rect 15334 10920 22650 10976
rect 22706 10920 22711 10976
rect 15334 10918 22711 10920
rect 7741 10915 7807 10918
rect 22645 10915 22711 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 6361 10842 6427 10845
rect 12617 10842 12683 10845
rect 0 10782 4906 10842
rect 0 10752 480 10782
rect 4846 10570 4906 10782
rect 6361 10840 12683 10842
rect 6361 10784 6366 10840
rect 6422 10784 12622 10840
rect 12678 10784 12683 10840
rect 6361 10782 12683 10784
rect 6361 10779 6427 10782
rect 12617 10779 12683 10782
rect 25037 10842 25103 10845
rect 27520 10842 28000 10872
rect 25037 10840 28000 10842
rect 25037 10784 25042 10840
rect 25098 10784 28000 10840
rect 25037 10782 28000 10784
rect 25037 10779 25103 10782
rect 27520 10752 28000 10782
rect 11145 10706 11211 10709
rect 17309 10706 17375 10709
rect 11145 10704 17375 10706
rect 11145 10648 11150 10704
rect 11206 10648 17314 10704
rect 17370 10648 17375 10704
rect 11145 10646 17375 10648
rect 11145 10643 11211 10646
rect 17309 10643 17375 10646
rect 12709 10570 12775 10573
rect 14641 10570 14707 10573
rect 16757 10570 16823 10573
rect 20805 10570 20871 10573
rect 25221 10570 25287 10573
rect 4846 10510 10748 10570
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 10688 10298 10748 10510
rect 12709 10568 14474 10570
rect 12709 10512 12714 10568
rect 12770 10512 14474 10568
rect 12709 10510 14474 10512
rect 12709 10507 12775 10510
rect 11053 10434 11119 10437
rect 13905 10434 13971 10437
rect 11053 10432 13971 10434
rect 11053 10376 11058 10432
rect 11114 10376 13910 10432
rect 13966 10376 13971 10432
rect 11053 10374 13971 10376
rect 14414 10434 14474 10510
rect 14641 10568 16823 10570
rect 14641 10512 14646 10568
rect 14702 10512 16762 10568
rect 16818 10512 16823 10568
rect 14641 10510 16823 10512
rect 14641 10507 14707 10510
rect 16757 10507 16823 10510
rect 19014 10568 25287 10570
rect 19014 10512 20810 10568
rect 20866 10512 25226 10568
rect 25282 10512 25287 10568
rect 19014 10510 25287 10512
rect 16941 10434 17007 10437
rect 14414 10432 17007 10434
rect 14414 10376 16946 10432
rect 17002 10376 17007 10432
rect 14414 10374 17007 10376
rect 11053 10371 11119 10374
rect 13905 10371 13971 10374
rect 16941 10371 17007 10374
rect 11789 10298 11855 10301
rect 19014 10298 19074 10510
rect 20805 10507 20871 10510
rect 25221 10507 25287 10510
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 10688 10296 19074 10298
rect 10688 10240 11794 10296
rect 11850 10240 19074 10296
rect 10688 10238 19074 10240
rect 11789 10235 11855 10238
rect 4981 10162 5047 10165
rect 6545 10162 6611 10165
rect 4981 10160 6611 10162
rect 4981 10104 4986 10160
rect 5042 10104 6550 10160
rect 6606 10104 6611 10160
rect 4981 10102 6611 10104
rect 4981 10099 5047 10102
rect 6545 10099 6611 10102
rect 19977 10162 20043 10165
rect 23473 10162 23539 10165
rect 19977 10160 23539 10162
rect 19977 10104 19982 10160
rect 20038 10104 23478 10160
rect 23534 10104 23539 10160
rect 19977 10102 23539 10104
rect 19977 10099 20043 10102
rect 23473 10099 23539 10102
rect 1853 10026 1919 10029
rect 4613 10026 4679 10029
rect 6361 10026 6427 10029
rect 7833 10026 7899 10029
rect 1853 10024 4679 10026
rect 1853 9968 1858 10024
rect 1914 9968 4618 10024
rect 4674 9968 4679 10024
rect 1853 9966 4679 9968
rect 1853 9963 1919 9966
rect 4613 9963 4679 9966
rect 5398 10024 7899 10026
rect 5398 9968 6366 10024
rect 6422 9968 7838 10024
rect 7894 9968 7899 10024
rect 5398 9966 7899 9968
rect 2129 9890 2195 9893
rect 5398 9890 5458 9966
rect 6361 9963 6427 9966
rect 7833 9963 7899 9966
rect 17309 10026 17375 10029
rect 25681 10026 25747 10029
rect 17309 10024 25747 10026
rect 17309 9968 17314 10024
rect 17370 9968 25686 10024
rect 25742 9968 25747 10024
rect 17309 9966 25747 9968
rect 17309 9963 17375 9966
rect 25681 9963 25747 9966
rect 2129 9888 5458 9890
rect 2129 9832 2134 9888
rect 2190 9832 5458 9888
rect 2129 9830 5458 9832
rect 7833 9890 7899 9893
rect 11513 9890 11579 9893
rect 7833 9888 11579 9890
rect 7833 9832 7838 9888
rect 7894 9832 11518 9888
rect 11574 9832 11579 9888
rect 7833 9830 11579 9832
rect 2129 9827 2195 9830
rect 7833 9827 7899 9830
rect 11513 9827 11579 9830
rect 5610 9824 5930 9825
rect 0 9754 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 565 9754 631 9757
rect 0 9752 631 9754
rect 0 9696 570 9752
rect 626 9696 631 9752
rect 0 9694 631 9696
rect 0 9664 480 9694
rect 565 9691 631 9694
rect 7097 9754 7163 9757
rect 8661 9754 8727 9757
rect 21449 9754 21515 9757
rect 25405 9754 25471 9757
rect 27520 9754 28000 9784
rect 7097 9752 7850 9754
rect 7097 9696 7102 9752
rect 7158 9696 7850 9752
rect 7097 9694 7850 9696
rect 7097 9691 7163 9694
rect 3509 9618 3575 9621
rect 7649 9618 7715 9621
rect 3509 9616 7715 9618
rect 3509 9560 3514 9616
rect 3570 9560 7654 9616
rect 7710 9560 7715 9616
rect 3509 9558 7715 9560
rect 3509 9555 3575 9558
rect 7649 9555 7715 9558
rect 7649 9482 7715 9485
rect 7790 9482 7850 9694
rect 8661 9752 9690 9754
rect 8661 9696 8666 9752
rect 8722 9696 9690 9752
rect 8661 9694 9690 9696
rect 8661 9691 8727 9694
rect 9630 9618 9690 9694
rect 21449 9752 23536 9754
rect 21449 9696 21454 9752
rect 21510 9696 23536 9752
rect 21449 9694 23536 9696
rect 21449 9691 21515 9694
rect 23476 9621 23536 9694
rect 25405 9752 28000 9754
rect 25405 9696 25410 9752
rect 25466 9696 28000 9752
rect 25405 9694 28000 9696
rect 25405 9691 25471 9694
rect 27520 9664 28000 9694
rect 14365 9618 14431 9621
rect 9630 9616 14431 9618
rect 9630 9560 14370 9616
rect 14426 9560 14431 9616
rect 9630 9558 14431 9560
rect 14365 9555 14431 9558
rect 23473 9616 23539 9621
rect 23473 9560 23478 9616
rect 23534 9560 23539 9616
rect 23473 9555 23539 9560
rect 7649 9480 7850 9482
rect 7649 9424 7654 9480
rect 7710 9424 7850 9480
rect 7649 9422 7850 9424
rect 8109 9482 8175 9485
rect 13537 9482 13603 9485
rect 8109 9480 13603 9482
rect 8109 9424 8114 9480
rect 8170 9424 13542 9480
rect 13598 9424 13603 9480
rect 8109 9422 13603 9424
rect 7649 9419 7715 9422
rect 8109 9419 8175 9422
rect 13537 9419 13603 9422
rect 6821 9346 6887 9349
rect 9489 9346 9555 9349
rect 6821 9344 9555 9346
rect 6821 9288 6826 9344
rect 6882 9288 9494 9344
rect 9550 9288 9555 9344
rect 6821 9286 9555 9288
rect 6821 9283 6887 9286
rect 9489 9283 9555 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 15929 9210 15995 9213
rect 18045 9210 18111 9213
rect 15929 9208 18111 9210
rect 15929 9152 15934 9208
rect 15990 9152 18050 9208
rect 18106 9152 18111 9208
rect 15929 9150 18111 9152
rect 15929 9147 15995 9150
rect 18045 9147 18111 9150
rect 2221 9074 2287 9077
rect 7833 9074 7899 9077
rect 2221 9072 7899 9074
rect 2221 9016 2226 9072
rect 2282 9016 7838 9072
rect 7894 9016 7899 9072
rect 2221 9014 7899 9016
rect 2221 9011 2287 9014
rect 7833 9011 7899 9014
rect 11973 9074 12039 9077
rect 14089 9074 14155 9077
rect 11973 9072 14155 9074
rect 11973 9016 11978 9072
rect 12034 9016 14094 9072
rect 14150 9016 14155 9072
rect 11973 9014 14155 9016
rect 11973 9011 12039 9014
rect 14089 9011 14155 9014
rect 14273 9074 14339 9077
rect 18505 9074 18571 9077
rect 14273 9072 18571 9074
rect 14273 9016 14278 9072
rect 14334 9016 18510 9072
rect 18566 9016 18571 9072
rect 14273 9014 18571 9016
rect 14273 9011 14339 9014
rect 18505 9011 18571 9014
rect 9673 8938 9739 8941
rect 15377 8938 15443 8941
rect 9673 8936 15443 8938
rect 9673 8880 9678 8936
rect 9734 8880 15382 8936
rect 15438 8880 15443 8936
rect 9673 8878 15443 8880
rect 9673 8875 9739 8878
rect 15377 8875 15443 8878
rect 24301 8938 24367 8941
rect 24945 8938 25011 8941
rect 24301 8936 25011 8938
rect 24301 8880 24306 8936
rect 24362 8880 24950 8936
rect 25006 8880 25011 8936
rect 24301 8878 25011 8880
rect 24301 8875 24367 8878
rect 24945 8875 25011 8878
rect 0 8802 480 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 0 8712 480 8742
rect 4061 8739 4127 8742
rect 15561 8802 15627 8805
rect 19333 8802 19399 8805
rect 15561 8800 19399 8802
rect 15561 8744 15566 8800
rect 15622 8744 19338 8800
rect 19394 8744 19399 8800
rect 15561 8742 19399 8744
rect 15561 8739 15627 8742
rect 19333 8739 19399 8742
rect 24761 8802 24827 8805
rect 27520 8802 28000 8832
rect 24761 8800 28000 8802
rect 24761 8744 24766 8800
rect 24822 8744 28000 8800
rect 24761 8742 28000 8744
rect 24761 8739 24827 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8742
rect 24277 8671 24597 8672
rect 8201 8666 8267 8669
rect 10593 8666 10659 8669
rect 8201 8664 10659 8666
rect 8201 8608 8206 8664
rect 8262 8608 10598 8664
rect 10654 8608 10659 8664
rect 8201 8606 10659 8608
rect 8201 8603 8267 8606
rect 10593 8603 10659 8606
rect 7925 8530 7991 8533
rect 9765 8530 9831 8533
rect 7925 8528 9831 8530
rect 7925 8472 7930 8528
rect 7986 8472 9770 8528
rect 9826 8472 9831 8528
rect 7925 8470 9831 8472
rect 7925 8467 7991 8470
rect 9765 8467 9831 8470
rect 6269 8394 6335 8397
rect 11237 8394 11303 8397
rect 6269 8392 11303 8394
rect 6269 8336 6274 8392
rect 6330 8336 11242 8392
rect 11298 8336 11303 8392
rect 6269 8334 11303 8336
rect 6269 8331 6335 8334
rect 11237 8331 11303 8334
rect 16297 8394 16363 8397
rect 20253 8394 20319 8397
rect 16297 8392 20319 8394
rect 16297 8336 16302 8392
rect 16358 8336 20258 8392
rect 20314 8336 20319 8392
rect 16297 8334 20319 8336
rect 16297 8331 16363 8334
rect 20253 8331 20319 8334
rect 23841 8394 23907 8397
rect 25589 8394 25655 8397
rect 23841 8392 25655 8394
rect 23841 8336 23846 8392
rect 23902 8336 25594 8392
rect 25650 8336 25655 8392
rect 23841 8334 25655 8336
rect 23841 8331 23907 8334
rect 25589 8331 25655 8334
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 20897 8122 20963 8125
rect 25221 8122 25287 8125
rect 20897 8120 25287 8122
rect 20897 8064 20902 8120
rect 20958 8064 25226 8120
rect 25282 8064 25287 8120
rect 20897 8062 25287 8064
rect 20897 8059 20963 8062
rect 25221 8059 25287 8062
rect 7373 7986 7439 7989
rect 15745 7986 15811 7989
rect 7373 7984 15811 7986
rect 7373 7928 7378 7984
rect 7434 7928 15750 7984
rect 15806 7928 15811 7984
rect 7373 7926 15811 7928
rect 7373 7923 7439 7926
rect 15745 7923 15811 7926
rect 10869 7850 10935 7853
rect 13353 7850 13419 7853
rect 23105 7850 23171 7853
rect 10869 7848 23171 7850
rect 10869 7792 10874 7848
rect 10930 7792 13358 7848
rect 13414 7792 23110 7848
rect 23166 7792 23171 7848
rect 10869 7790 23171 7792
rect 10869 7787 10935 7790
rect 13353 7787 13419 7790
rect 23105 7787 23171 7790
rect 0 7714 480 7744
rect 1577 7714 1643 7717
rect 27520 7714 28000 7744
rect 0 7712 1643 7714
rect 0 7656 1582 7712
rect 1638 7656 1643 7712
rect 0 7654 1643 7656
rect 0 7624 480 7654
rect 1577 7651 1643 7654
rect 24764 7654 28000 7714
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 4889 7442 4955 7445
rect 7281 7442 7347 7445
rect 4889 7440 7347 7442
rect 4889 7384 4894 7440
rect 4950 7384 7286 7440
rect 7342 7384 7347 7440
rect 4889 7382 7347 7384
rect 4889 7379 4955 7382
rect 7281 7379 7347 7382
rect 13721 7442 13787 7445
rect 16573 7442 16639 7445
rect 20989 7442 21055 7445
rect 13721 7440 21055 7442
rect 13721 7384 13726 7440
rect 13782 7384 16578 7440
rect 16634 7384 20994 7440
rect 21050 7384 21055 7440
rect 13721 7382 21055 7384
rect 13721 7379 13787 7382
rect 16573 7379 16639 7382
rect 20989 7379 21055 7382
rect 23565 7442 23631 7445
rect 24764 7442 24824 7654
rect 27520 7624 28000 7654
rect 23565 7440 24824 7442
rect 23565 7384 23570 7440
rect 23626 7384 24824 7440
rect 23565 7382 24824 7384
rect 23565 7379 23631 7382
rect 3969 7306 4035 7309
rect 12893 7306 12959 7309
rect 3969 7304 12959 7306
rect 3969 7248 3974 7304
rect 4030 7248 12898 7304
rect 12954 7248 12959 7304
rect 3969 7246 12959 7248
rect 3969 7243 4035 7246
rect 12893 7243 12959 7246
rect 17125 7306 17191 7309
rect 23473 7306 23539 7309
rect 17125 7304 23539 7306
rect 17125 7248 17130 7304
rect 17186 7248 23478 7304
rect 23534 7248 23539 7304
rect 17125 7246 23539 7248
rect 17125 7243 17191 7246
rect 23473 7243 23539 7246
rect 3049 7170 3115 7173
rect 4153 7170 4219 7173
rect 3049 7168 4219 7170
rect 3049 7112 3054 7168
rect 3110 7112 4158 7168
rect 4214 7112 4219 7168
rect 3049 7110 4219 7112
rect 3049 7107 3115 7110
rect 4153 7107 4219 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 5717 7034 5783 7037
rect 5993 7034 6059 7037
rect 8477 7034 8543 7037
rect 5717 7032 8543 7034
rect 5717 6976 5722 7032
rect 5778 6976 5998 7032
rect 6054 6976 8482 7032
rect 8538 6976 8543 7032
rect 5717 6974 8543 6976
rect 5717 6971 5783 6974
rect 5993 6971 6059 6974
rect 8477 6971 8543 6974
rect 16941 7034 17007 7037
rect 19425 7034 19491 7037
rect 16941 7032 19491 7034
rect 16941 6976 16946 7032
rect 17002 6976 19430 7032
rect 19486 6976 19491 7032
rect 16941 6974 19491 6976
rect 16941 6971 17007 6974
rect 19425 6971 19491 6974
rect 13537 6762 13603 6765
rect 22829 6762 22895 6765
rect 13537 6760 22895 6762
rect 13537 6704 13542 6760
rect 13598 6704 22834 6760
rect 22890 6704 22895 6760
rect 13537 6702 22895 6704
rect 13537 6699 13603 6702
rect 22829 6699 22895 6702
rect 0 6626 480 6656
rect 4245 6626 4311 6629
rect 0 6624 4311 6626
rect 0 6568 4250 6624
rect 4306 6568 4311 6624
rect 0 6566 4311 6568
rect 0 6536 480 6566
rect 4245 6563 4311 6566
rect 25405 6626 25471 6629
rect 27520 6626 28000 6656
rect 25405 6624 28000 6626
rect 25405 6568 25410 6624
rect 25466 6568 28000 6624
rect 25405 6566 28000 6568
rect 25405 6563 25471 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 14181 6490 14247 6493
rect 6134 6488 14247 6490
rect 6134 6432 14186 6488
rect 14242 6432 14247 6488
rect 6134 6430 14247 6432
rect 4981 6354 5047 6357
rect 6134 6354 6194 6430
rect 14181 6427 14247 6430
rect 16205 6490 16271 6493
rect 17953 6490 18019 6493
rect 16205 6488 18019 6490
rect 16205 6432 16210 6488
rect 16266 6432 17958 6488
rect 18014 6432 18019 6488
rect 16205 6430 18019 6432
rect 16205 6427 16271 6430
rect 17953 6427 18019 6430
rect 19241 6490 19307 6493
rect 21725 6490 21791 6493
rect 19241 6488 21791 6490
rect 19241 6432 19246 6488
rect 19302 6432 21730 6488
rect 21786 6432 21791 6488
rect 19241 6430 21791 6432
rect 19241 6427 19307 6430
rect 21725 6427 21791 6430
rect 4981 6352 6194 6354
rect 4981 6296 4986 6352
rect 5042 6296 6194 6352
rect 4981 6294 6194 6296
rect 12065 6354 12131 6357
rect 18505 6354 18571 6357
rect 12065 6352 18571 6354
rect 12065 6296 12070 6352
rect 12126 6296 18510 6352
rect 18566 6296 18571 6352
rect 12065 6294 18571 6296
rect 4981 6291 5047 6294
rect 12065 6291 12131 6294
rect 18505 6291 18571 6294
rect 4061 6218 4127 6221
rect 5717 6218 5783 6221
rect 4061 6216 5783 6218
rect 4061 6160 4066 6216
rect 4122 6160 5722 6216
rect 5778 6160 5783 6216
rect 4061 6158 5783 6160
rect 4061 6155 4127 6158
rect 5717 6155 5783 6158
rect 8753 6218 8819 6221
rect 14089 6218 14155 6221
rect 8753 6216 14155 6218
rect 8753 6160 8758 6216
rect 8814 6160 14094 6216
rect 14150 6160 14155 6216
rect 8753 6158 14155 6160
rect 8753 6155 8819 6158
rect 14089 6155 14155 6158
rect 19241 6218 19307 6221
rect 22185 6218 22251 6221
rect 19241 6216 22251 6218
rect 19241 6160 19246 6216
rect 19302 6160 22190 6216
rect 22246 6160 22251 6216
rect 19241 6158 22251 6160
rect 19241 6155 19307 6158
rect 22185 6155 22251 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 17585 5946 17651 5949
rect 19057 5946 19123 5949
rect 17585 5944 19123 5946
rect 17585 5888 17590 5944
rect 17646 5888 19062 5944
rect 19118 5888 19123 5944
rect 17585 5886 19123 5888
rect 17585 5883 17651 5886
rect 19057 5883 19123 5886
rect 21173 5810 21239 5813
rect 26509 5810 26575 5813
rect 21173 5808 26575 5810
rect 21173 5752 21178 5808
rect 21234 5752 26514 5808
rect 26570 5752 26575 5808
rect 21173 5750 26575 5752
rect 21173 5747 21239 5750
rect 26509 5747 26575 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 3509 5674 3575 5677
rect 6545 5674 6611 5677
rect 3509 5672 6611 5674
rect 3509 5616 3514 5672
rect 3570 5616 6550 5672
rect 6606 5616 6611 5672
rect 3509 5614 6611 5616
rect 3509 5611 3575 5614
rect 6545 5611 6611 5614
rect 8109 5674 8175 5677
rect 9673 5674 9739 5677
rect 8109 5672 9739 5674
rect 8109 5616 8114 5672
rect 8170 5616 9678 5672
rect 9734 5616 9739 5672
rect 8109 5614 9739 5616
rect 8109 5611 8175 5614
rect 9673 5611 9739 5614
rect 14181 5674 14247 5677
rect 14365 5674 14431 5677
rect 15377 5674 15443 5677
rect 14181 5672 15443 5674
rect 14181 5616 14186 5672
rect 14242 5616 14370 5672
rect 14426 5616 15382 5672
rect 15438 5616 15443 5672
rect 14181 5614 15443 5616
rect 14181 5611 14247 5614
rect 14365 5611 14431 5614
rect 15377 5611 15443 5614
rect 16849 5674 16915 5677
rect 21449 5674 21515 5677
rect 16849 5672 21515 5674
rect 16849 5616 16854 5672
rect 16910 5616 21454 5672
rect 21510 5616 21515 5672
rect 16849 5614 21515 5616
rect 16849 5611 16915 5614
rect 21449 5611 21515 5614
rect 24669 5674 24735 5677
rect 27520 5674 28000 5704
rect 24669 5672 28000 5674
rect 24669 5616 24674 5672
rect 24730 5616 28000 5672
rect 24669 5614 28000 5616
rect 24669 5611 24735 5614
rect 27520 5584 28000 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 13629 5402 13695 5405
rect 7422 5400 14474 5402
rect 7422 5344 13634 5400
rect 13690 5344 14474 5400
rect 7422 5342 14474 5344
rect 4337 5266 4403 5269
rect 7281 5266 7347 5269
rect 4337 5264 7347 5266
rect 4337 5208 4342 5264
rect 4398 5208 7286 5264
rect 7342 5208 7347 5264
rect 4337 5206 7347 5208
rect 4337 5203 4403 5206
rect 7281 5203 7347 5206
rect 4613 5130 4679 5133
rect 7422 5130 7482 5342
rect 13629 5339 13695 5342
rect 11881 5266 11947 5269
rect 14181 5266 14247 5269
rect 11881 5264 14247 5266
rect 11881 5208 11886 5264
rect 11942 5208 14186 5264
rect 14242 5208 14247 5264
rect 11881 5206 14247 5208
rect 14414 5266 14474 5342
rect 14641 5266 14707 5269
rect 15653 5266 15719 5269
rect 14414 5264 15719 5266
rect 14414 5208 14646 5264
rect 14702 5208 15658 5264
rect 15714 5208 15719 5264
rect 14414 5206 15719 5208
rect 11881 5203 11947 5206
rect 14181 5203 14247 5206
rect 14641 5203 14707 5206
rect 15653 5203 15719 5206
rect 14089 5130 14155 5133
rect 4613 5128 7482 5130
rect 4613 5072 4618 5128
rect 4674 5072 7482 5128
rect 4613 5070 7482 5072
rect 7606 5128 14155 5130
rect 7606 5072 14094 5128
rect 14150 5072 14155 5128
rect 7606 5070 14155 5072
rect 4613 5067 4679 5070
rect 4061 4994 4127 4997
rect 7606 4994 7666 5070
rect 14089 5067 14155 5070
rect 14273 5130 14339 5133
rect 17953 5130 18019 5133
rect 20713 5130 20779 5133
rect 14273 5128 20779 5130
rect 14273 5072 14278 5128
rect 14334 5072 17958 5128
rect 18014 5072 20718 5128
rect 20774 5072 20779 5128
rect 14273 5070 20779 5072
rect 14273 5067 14339 5070
rect 17953 5067 18019 5070
rect 20713 5067 20779 5070
rect 4061 4992 7666 4994
rect 4061 4936 4066 4992
rect 4122 4936 7666 4992
rect 4061 4934 7666 4936
rect 4061 4931 4127 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 15561 4858 15627 4861
rect 19425 4858 19491 4861
rect 15561 4856 19491 4858
rect 15561 4800 15566 4856
rect 15622 4800 19430 4856
rect 19486 4800 19491 4856
rect 15561 4798 19491 4800
rect 15561 4795 15627 4798
rect 19425 4795 19491 4798
rect 2773 4722 2839 4725
rect 4245 4722 4311 4725
rect 2773 4720 4311 4722
rect 2773 4664 2778 4720
rect 2834 4664 4250 4720
rect 4306 4664 4311 4720
rect 2773 4662 4311 4664
rect 2773 4659 2839 4662
rect 4245 4659 4311 4662
rect 17585 4722 17651 4725
rect 17585 4720 18338 4722
rect 17585 4664 17590 4720
rect 17646 4664 18338 4720
rect 17585 4662 18338 4664
rect 17585 4659 17651 4662
rect 0 4586 480 4616
rect 1577 4586 1643 4589
rect 0 4584 1643 4586
rect 0 4528 1582 4584
rect 1638 4528 1643 4584
rect 0 4526 1643 4528
rect 0 4496 480 4526
rect 1577 4523 1643 4526
rect 2681 4586 2747 4589
rect 12893 4586 12959 4589
rect 2681 4584 12959 4586
rect 2681 4528 2686 4584
rect 2742 4528 12898 4584
rect 12954 4528 12959 4584
rect 2681 4526 12959 4528
rect 2681 4523 2747 4526
rect 12893 4523 12959 4526
rect 14273 4586 14339 4589
rect 18278 4586 18338 4662
rect 21817 4586 21883 4589
rect 22277 4586 22343 4589
rect 14273 4584 18200 4586
rect 14273 4528 14278 4584
rect 14334 4528 18200 4584
rect 14273 4526 18200 4528
rect 18278 4584 22343 4586
rect 18278 4528 21822 4584
rect 21878 4528 22282 4584
rect 22338 4528 22343 4584
rect 18278 4526 22343 4528
rect 14273 4523 14339 4526
rect 18140 4450 18200 4526
rect 21817 4523 21883 4526
rect 22277 4523 22343 4526
rect 25405 4586 25471 4589
rect 27520 4586 28000 4616
rect 25405 4584 28000 4586
rect 25405 4528 25410 4584
rect 25466 4528 28000 4584
rect 25405 4526 28000 4528
rect 25405 4523 25471 4526
rect 27520 4496 28000 4526
rect 18140 4390 23858 4450
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 2589 4178 2655 4181
rect 6545 4178 6611 4181
rect 2589 4176 6611 4178
rect 2589 4120 2594 4176
rect 2650 4120 6550 4176
rect 6606 4120 6611 4176
rect 2589 4118 6611 4120
rect 2589 4115 2655 4118
rect 6545 4115 6611 4118
rect 17769 4178 17835 4181
rect 22553 4178 22619 4181
rect 17769 4176 22619 4178
rect 17769 4120 17774 4176
rect 17830 4120 22558 4176
rect 22614 4120 22619 4176
rect 17769 4118 22619 4120
rect 17769 4115 17835 4118
rect 22553 4115 22619 4118
rect 10593 4042 10659 4045
rect 15193 4042 15259 4045
rect 10593 4040 15259 4042
rect 10593 3984 10598 4040
rect 10654 3984 15198 4040
rect 15254 3984 15259 4040
rect 10593 3982 15259 3984
rect 23798 4042 23858 4390
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 25497 4042 25563 4045
rect 23798 4040 25563 4042
rect 23798 3984 25502 4040
rect 25558 3984 25563 4040
rect 23798 3982 25563 3984
rect 10593 3979 10659 3982
rect 15193 3979 15259 3982
rect 25497 3979 25563 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 7373 3634 7439 3637
rect 15377 3634 15443 3637
rect 7373 3632 15443 3634
rect 7373 3576 7378 3632
rect 7434 3576 15382 3632
rect 15438 3576 15443 3632
rect 7373 3574 15443 3576
rect 7373 3571 7439 3574
rect 15377 3571 15443 3574
rect 15929 3634 15995 3637
rect 18413 3634 18479 3637
rect 15929 3632 18479 3634
rect 15929 3576 15934 3632
rect 15990 3576 18418 3632
rect 18474 3576 18479 3632
rect 15929 3574 18479 3576
rect 15929 3571 15995 3574
rect 18413 3571 18479 3574
rect 0 3498 480 3528
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3408 480 3438
rect 1577 3435 1643 3438
rect 6913 3498 6979 3501
rect 8201 3498 8267 3501
rect 6913 3496 8267 3498
rect 6913 3440 6918 3496
rect 6974 3440 8206 3496
rect 8262 3440 8267 3496
rect 6913 3438 8267 3440
rect 6913 3435 6979 3438
rect 8201 3435 8267 3438
rect 9397 3498 9463 3501
rect 11053 3498 11119 3501
rect 9397 3496 11119 3498
rect 9397 3440 9402 3496
rect 9458 3440 11058 3496
rect 11114 3440 11119 3496
rect 9397 3438 11119 3440
rect 9397 3435 9463 3438
rect 11053 3435 11119 3438
rect 11605 3498 11671 3501
rect 12617 3498 12683 3501
rect 11605 3496 12683 3498
rect 11605 3440 11610 3496
rect 11666 3440 12622 3496
rect 12678 3440 12683 3496
rect 11605 3438 12683 3440
rect 11605 3435 11671 3438
rect 12617 3435 12683 3438
rect 14273 3498 14339 3501
rect 23565 3498 23631 3501
rect 14273 3496 23631 3498
rect 14273 3440 14278 3496
rect 14334 3440 23570 3496
rect 23626 3440 23631 3496
rect 14273 3438 23631 3440
rect 14273 3435 14339 3438
rect 23565 3435 23631 3438
rect 25405 3498 25471 3501
rect 27520 3498 28000 3528
rect 25405 3496 28000 3498
rect 25405 3440 25410 3496
rect 25466 3440 28000 3496
rect 25405 3438 28000 3440
rect 25405 3435 25471 3438
rect 27520 3408 28000 3438
rect 6177 3362 6243 3365
rect 11053 3362 11119 3365
rect 6177 3360 11119 3362
rect 6177 3304 6182 3360
rect 6238 3304 11058 3360
rect 11114 3304 11119 3360
rect 6177 3302 11119 3304
rect 6177 3299 6243 3302
rect 11053 3299 11119 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2037 3226 2103 3229
rect 3877 3226 3943 3229
rect 13445 3226 13511 3229
rect 2037 3224 3943 3226
rect 2037 3168 2042 3224
rect 2098 3168 3882 3224
rect 3938 3168 3943 3224
rect 2037 3166 3943 3168
rect 2037 3163 2103 3166
rect 3877 3163 3943 3166
rect 6134 3224 13511 3226
rect 6134 3168 13450 3224
rect 13506 3168 13511 3224
rect 6134 3166 13511 3168
rect 5165 3090 5231 3093
rect 6134 3090 6194 3166
rect 13445 3163 13511 3166
rect 5165 3088 6194 3090
rect 5165 3032 5170 3088
rect 5226 3032 6194 3088
rect 5165 3030 6194 3032
rect 6269 3090 6335 3093
rect 13813 3090 13879 3093
rect 6269 3088 13879 3090
rect 6269 3032 6274 3088
rect 6330 3032 13818 3088
rect 13874 3032 13879 3088
rect 6269 3030 13879 3032
rect 5165 3027 5231 3030
rect 6269 3027 6335 3030
rect 13813 3027 13879 3030
rect 14917 3090 14983 3093
rect 16573 3090 16639 3093
rect 14917 3088 16639 3090
rect 14917 3032 14922 3088
rect 14978 3032 16578 3088
rect 16634 3032 16639 3088
rect 14917 3030 16639 3032
rect 14917 3027 14983 3030
rect 16573 3027 16639 3030
rect 23289 3090 23355 3093
rect 24669 3090 24735 3093
rect 23289 3088 24735 3090
rect 23289 3032 23294 3088
rect 23350 3032 24674 3088
rect 24730 3032 24735 3088
rect 23289 3030 24735 3032
rect 23289 3027 23355 3030
rect 24669 3027 24735 3030
rect 8017 2954 8083 2957
rect 8937 2954 9003 2957
rect 8017 2952 9003 2954
rect 8017 2896 8022 2952
rect 8078 2896 8942 2952
rect 8998 2896 9003 2952
rect 8017 2894 9003 2896
rect 8017 2891 8083 2894
rect 8937 2891 9003 2894
rect 13629 2818 13695 2821
rect 15929 2818 15995 2821
rect 13629 2816 15995 2818
rect 13629 2760 13634 2816
rect 13690 2760 15934 2816
rect 15990 2760 15995 2816
rect 13629 2758 15995 2760
rect 13629 2755 13695 2758
rect 15929 2755 15995 2758
rect 22645 2818 22711 2821
rect 27429 2818 27495 2821
rect 22645 2816 27495 2818
rect 22645 2760 22650 2816
rect 22706 2760 27434 2816
rect 27490 2760 27495 2816
rect 22645 2758 27495 2760
rect 22645 2755 22711 2758
rect 27429 2755 27495 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 6361 2682 6427 2685
rect 9581 2682 9647 2685
rect 6361 2680 9647 2682
rect 6361 2624 6366 2680
rect 6422 2624 9586 2680
rect 9642 2624 9647 2680
rect 6361 2622 9647 2624
rect 6361 2619 6427 2622
rect 9581 2619 9647 2622
rect 10685 2682 10751 2685
rect 14181 2682 14247 2685
rect 10685 2680 14247 2682
rect 10685 2624 10690 2680
rect 10746 2624 14186 2680
rect 14242 2624 14247 2680
rect 10685 2622 14247 2624
rect 10685 2619 10751 2622
rect 14181 2619 14247 2622
rect 21265 2682 21331 2685
rect 25405 2682 25471 2685
rect 21265 2680 25471 2682
rect 21265 2624 21270 2680
rect 21326 2624 25410 2680
rect 25466 2624 25471 2680
rect 21265 2622 25471 2624
rect 21265 2619 21331 2622
rect 25405 2619 25471 2622
rect 0 2546 480 2576
rect 3877 2546 3943 2549
rect 0 2544 3943 2546
rect 0 2488 3882 2544
rect 3938 2488 3943 2544
rect 0 2486 3943 2488
rect 0 2456 480 2486
rect 3877 2483 3943 2486
rect 4797 2546 4863 2549
rect 16297 2546 16363 2549
rect 4797 2544 16363 2546
rect 4797 2488 4802 2544
rect 4858 2488 16302 2544
rect 16358 2488 16363 2544
rect 4797 2486 16363 2488
rect 4797 2483 4863 2486
rect 16297 2483 16363 2486
rect 19241 2546 19307 2549
rect 22185 2546 22251 2549
rect 19241 2544 22251 2546
rect 19241 2488 19246 2544
rect 19302 2488 22190 2544
rect 22246 2488 22251 2544
rect 19241 2486 22251 2488
rect 19241 2483 19307 2486
rect 22185 2483 22251 2486
rect 24761 2546 24827 2549
rect 27520 2546 28000 2576
rect 24761 2544 28000 2546
rect 24761 2488 24766 2544
rect 24822 2488 28000 2544
rect 24761 2486 28000 2488
rect 24761 2483 24827 2486
rect 27520 2456 28000 2486
rect 9213 2410 9279 2413
rect 13261 2410 13327 2413
rect 14273 2410 14339 2413
rect 9213 2408 14339 2410
rect 9213 2352 9218 2408
rect 9274 2352 13266 2408
rect 13322 2352 14278 2408
rect 14334 2352 14339 2408
rect 9213 2350 14339 2352
rect 9213 2347 9279 2350
rect 13261 2347 13327 2350
rect 14273 2347 14339 2350
rect 16021 2410 16087 2413
rect 24853 2410 24919 2413
rect 16021 2408 24919 2410
rect 16021 2352 16026 2408
rect 16082 2352 24858 2408
rect 24914 2352 24919 2408
rect 16021 2350 24919 2352
rect 16021 2347 16087 2350
rect 24853 2347 24919 2350
rect 15745 2274 15811 2277
rect 20713 2274 20779 2277
rect 15745 2272 20779 2274
rect 15745 2216 15750 2272
rect 15806 2216 20718 2272
rect 20774 2216 20779 2272
rect 15745 2214 20779 2216
rect 15745 2211 15811 2214
rect 20713 2211 20779 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 17401 2138 17467 2141
rect 21541 2138 21607 2141
rect 17401 2136 21607 2138
rect 17401 2080 17406 2136
rect 17462 2080 21546 2136
rect 21602 2080 21607 2136
rect 17401 2078 21607 2080
rect 17401 2075 17467 2078
rect 21541 2075 21607 2078
rect 14457 2002 14523 2005
rect 19701 2002 19767 2005
rect 14457 2000 19767 2002
rect 14457 1944 14462 2000
rect 14518 1944 19706 2000
rect 19762 1944 19767 2000
rect 14457 1942 19767 1944
rect 14457 1939 14523 1942
rect 19701 1939 19767 1942
rect 23657 2002 23723 2005
rect 26417 2002 26483 2005
rect 23657 2000 26483 2002
rect 23657 1944 23662 2000
rect 23718 1944 26422 2000
rect 26478 1944 26483 2000
rect 23657 1942 26483 1944
rect 23657 1939 23723 1942
rect 26417 1939 26483 1942
rect 8845 1866 8911 1869
rect 16757 1866 16823 1869
rect 8845 1864 16823 1866
rect 8845 1808 8850 1864
rect 8906 1808 16762 1864
rect 16818 1808 16823 1864
rect 8845 1806 16823 1808
rect 8845 1803 8911 1806
rect 16757 1803 16823 1806
rect 10225 1730 10291 1733
rect 16941 1730 17007 1733
rect 10225 1728 17007 1730
rect 10225 1672 10230 1728
rect 10286 1672 16946 1728
rect 17002 1672 17007 1728
rect 10225 1670 17007 1672
rect 10225 1667 10291 1670
rect 16941 1667 17007 1670
rect 4429 1594 4495 1597
rect 15285 1594 15351 1597
rect 4429 1592 15351 1594
rect 4429 1536 4434 1592
rect 4490 1536 15290 1592
rect 15346 1536 15351 1592
rect 4429 1534 15351 1536
rect 4429 1531 4495 1534
rect 15285 1531 15351 1534
rect 0 1458 480 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 480 1398
rect 1577 1395 1643 1398
rect 23013 1458 23079 1461
rect 27520 1458 28000 1488
rect 23013 1456 28000 1458
rect 23013 1400 23018 1456
rect 23074 1400 28000 1456
rect 23013 1398 28000 1400
rect 23013 1395 23079 1398
rect 27520 1368 28000 1398
rect 0 506 480 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 480 446
rect 2773 443 2839 446
rect 26141 506 26207 509
rect 27520 506 28000 536
rect 26141 504 28000 506
rect 26141 448 26146 504
rect 26202 448 28000 504
rect 26141 446 28000 448
rect 26141 443 26207 446
rect 27520 416 28000 446
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 9812 19212 9876 19276
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 4476 17036 4540 17100
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 9812 12820 9876 12884
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 4476 11596 4540 11660
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9811 19276 9877 19277
rect 9811 19212 9812 19276
rect 9876 19212 9877 19276
rect 9811 19211 9877 19212
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 4475 17100 4541 17101
rect 4475 17036 4476 17100
rect 4540 17036 4541 17100
rect 4475 17035 4541 17036
rect 4478 11661 4538 17035
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 9814 12885 9874 19211
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 9811 12884 9877 12885
rect 9811 12820 9812 12884
rect 9876 12820 9877 12884
rect 9811 12819 9877 12820
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 4475 11660 4541 11661
rect 4475 11596 4476 11660
rect 4540 11596 4541 11660
rect 4475 11595 4541 11596
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _228_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_11
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 130 592
use scs8hd_conb_1  _215_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_1  _106_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_30
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _090_
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_18 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_8  _124_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_68
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_142
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_149
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _246_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _245_
timestamp 1586364061
transform 1 0 15548 0 -1 2720
box -38 -48 406 592
use scs8hd_nor4_4  _170_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 1602 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__D
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_161
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18400 0 -1 2720
box -38 -48 1050 592
use scs8hd_nor4_4  _172_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1602 592
use scs8hd_decap_3  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_201
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_235
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_270 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_13
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_or3_4  _125_
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_79
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_116
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_133
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _171_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_176
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _174_
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_229
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_241
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_245
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _160_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_78
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_82
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_144
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__C
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_169
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _173_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_218
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 314 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_270
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_20
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_24
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_28
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_45 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_53
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_57
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_98
timestamp 1586364061
transform 1 0 10120 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_112
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__D
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__D
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23460 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_262
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_25
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_29
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_48
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 406 592
use scs8hd_inv_8  _098_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 314 592
use scs8hd_or3_4  _089_
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 866 592
use scs8hd_or3_4  _114_
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_233
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_241
timestamp 1586364061
transform 1 0 23276 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_249
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_261
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_9
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_24
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_28
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_or3_4  _108_
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 866 592
use scs8hd_or3_4  _105_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_119
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_nor4_4  _176_
timestamp 1586364061
transform 1 0 15364 0 -1 5984
box -38 -48 1602 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_172
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_176
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__D
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__C
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _175_
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _179_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__C
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_205
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_197
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_219
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  _244_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_230
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_226
timestamp 1586364061
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_223
timestamp 1586364061
transform 1 0 21620 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 21804 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_240
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_249
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_250
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_261
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_265
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_20
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_24
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_28
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 590 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_116
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__D
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _177_
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__D
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _180_
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_203
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 20976 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_220
timestamp 1586364061
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_257
timestamp 1586364061
transform 1 0 24748 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_269
timestamp 1586364061
transform 1 0 25852 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_28
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _102_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _095_
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_161
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__D
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__C
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 314 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_270
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_11
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_58
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_75
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_81
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_85
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 590 592
use scs8hd_buf_1  _085_
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__C
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use scs8hd_or3_4  _153_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _112_
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__C
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _181_
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__184__D
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__C
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_241
timestamp 1586364061
transform 1 0 23276 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _220_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _145_
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_137
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _185_
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__185__D
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _183_
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__D
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_202
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_206
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 590 592
use scs8hd_decap_3  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_259
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_275
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_14
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_12_65
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_69
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_133
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 130 592
use scs8hd_nor4_4  _186_
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__C
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 314 592
use scs8hd_nor4_4  _184_
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_201
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_209
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_240
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_243
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_262
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_24
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _221_
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_114
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_131
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_146
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_or3_4  _116_
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__C
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__C
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__D
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _182_
timestamp 1586364061
transform 1 0 18124 0 1 9248
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_206
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 1050 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_226
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_221
timestamp 1586364061
transform 1 0 21436 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_233
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_254
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_250
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_260
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_270
timestamp 1586364061
transform 1 0 25944 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 1050 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_129
timestamp 1586364061
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_133
timestamp 1586364061
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_146
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_13
timestamp 1586364061
transform 1 0 2300 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_207
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_220
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_231
timestamp 1586364061
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_243
timestamp 1586364061
transform 1 0 23460 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_46
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 406 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 130 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_210
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_227
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_231
timestamp 1586364061
transform 1 0 22356 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_248
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_252
timestamp 1586364061
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_267
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_8
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_104
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_108
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_116
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_1  _117_
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_161
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 590 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_205
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_218
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_226
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_244
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_248
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_8
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 1050 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_39
timestamp 1586364061
transform 1 0 4692 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_58
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_55
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _136_
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_174
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _137_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_204
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_198
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_221
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_21
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_32
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_152
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_167
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _135_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 774 592
use scs8hd_buf_1  _178_
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_215
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_219
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_234
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_242
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_conb_1  _206_
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_250
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_262
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_21
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_25
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_52
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_72
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_127
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_174
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_203
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_218
timestamp 1586364061
transform 1 0 21160 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_229
timestamp 1586364061
transform 1 0 22172 0 -1 14688
box -38 -48 774 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 22908 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_240
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_262
timestamp 1586364061
transform 1 0 25208 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_6
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_14
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_26
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_43
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_133
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 314 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_209
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_213
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 590 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_226
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_233
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_249
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24196 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_253
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_260
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_272
timestamp 1586364061
transform 1 0 26128 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_20
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_24
timestamp 1586364061
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_111
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_114
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_124
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_160
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_172
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_189
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _207_
timestamp 1586364061
transform 1 0 21528 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_221
timestamp 1586364061
transform 1 0 21436 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_225
timestamp 1586364061
transform 1 0 21804 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_237
timestamp 1586364061
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_249
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_261
timestamp 1586364061
transform 1 0 25116 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_273
timestamp 1586364061
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 1472 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_24
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_68
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_150
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_160
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_172
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_176
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use scs8hd_buf_1  _162_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_198
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_222
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_242
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_262
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_8
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_26
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_20
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_37
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_48
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 6532 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_68
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_72
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 590 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_87
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_91
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_106
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 590 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_148
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_151
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _169_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_1  _161_
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_192
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_204
timestamp 1586364061
transform 1 0 19872 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_38
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_50
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 406 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_57
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _205_
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_96
timestamp 1586364061
transform 1 0 9936 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_119
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_21
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_28
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_45
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_60
timestamp 1586364061
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_94
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_17
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_35
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_82
timestamp 1586364061
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_90
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_17
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_28
timestamp 1586364061
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_17
timestamp 1586364061
transform 1 0 2668 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_29
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_35
timestamp 1586364061
transform 1 0 4324 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_17
timestamp 1586364061
transform 1 0 2668 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_21
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_25
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_37
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_49
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_127
timestamp 1586364061
transform 1 0 12788 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_131
timestamp 1586364061
transform 1 0 13156 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_262
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_274
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_46
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_148
timestamp 1586364061
transform 1 0 14720 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_160
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_172
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_180
timestamp 1586364061
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 11978 0 12034 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 12990 0 13046 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 13910 0 13966 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 14922 0 14978 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 15842 0 15898 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 16854 0 16910 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 17774 0 17830 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 478 0 534 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 10046 0 10102 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 0 17960 480 18080 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 6536 480 6656 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 0 7624 480 7744 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 8712 480 8832 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 27520 17008 28000 17128 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 27520 2456 28000 2576 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 27520 5584 28000 5704 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 27520 9664 28000 9784 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal2 s 27434 0 27490 480 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 data_in
port 63 nsew default input
rlabel metal2 s 11058 0 11114 480 6 enable
port 64 nsew default input
rlabel metal3 s 0 416 480 536 6 left_bottom_grid_pin_12_
port 65 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_11_
port 66 nsew default input
rlabel metal3 s 0 26256 480 26376 6 left_top_grid_pin_13_
port 67 nsew default input
rlabel metal3 s 0 27344 480 27464 6 left_top_grid_pin_15_
port 68 nsew default input
rlabel metal3 s 0 20000 480 20120 6 left_top_grid_pin_1_
port 69 nsew default input
rlabel metal3 s 0 21088 480 21208 6 left_top_grid_pin_3_
port 70 nsew default input
rlabel metal3 s 0 22176 480 22296 6 left_top_grid_pin_5_
port 71 nsew default input
rlabel metal3 s 0 23128 480 23248 6 left_top_grid_pin_7_
port 72 nsew default input
rlabel metal3 s 0 24216 480 24336 6 left_top_grid_pin_9_
port 73 nsew default input
rlabel metal3 s 27520 416 28000 536 6 right_bottom_grid_pin_12_
port 74 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_11_
port 75 nsew default input
rlabel metal3 s 27520 26256 28000 26376 6 right_top_grid_pin_13_
port 76 nsew default input
rlabel metal3 s 27520 27344 28000 27464 6 right_top_grid_pin_15_
port 77 nsew default input
rlabel metal3 s 27520 20000 28000 20120 6 right_top_grid_pin_1_
port 78 nsew default input
rlabel metal3 s 27520 21088 28000 21208 6 right_top_grid_pin_3_
port 79 nsew default input
rlabel metal3 s 27520 22176 28000 22296 6 right_top_grid_pin_5_
port 80 nsew default input
rlabel metal3 s 27520 23128 28000 23248 6 right_top_grid_pin_7_
port 81 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 right_top_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27464
<< end >>
