magic
tech sky130A
magscale 1 2
timestamp 1608157631
<< obsli1 >>
rect 1104 2159 21620 20145
<< obsm1 >>
rect 198 280 22618 21820
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 1030 22000 1086 22800
rect 1490 22000 1546 22800
rect 1950 22000 2006 22800
rect 2410 22000 2466 22800
rect 2870 22000 2926 22800
rect 3330 22000 3386 22800
rect 3790 22000 3846 22800
rect 4250 22000 4306 22800
rect 4710 22000 4766 22800
rect 5170 22000 5226 22800
rect 5630 22000 5686 22800
rect 6090 22000 6146 22800
rect 6550 22000 6606 22800
rect 7010 22000 7066 22800
rect 7470 22000 7526 22800
rect 7930 22000 7986 22800
rect 8390 22000 8446 22800
rect 8850 22000 8906 22800
rect 9310 22000 9366 22800
rect 9770 22000 9826 22800
rect 10230 22000 10286 22800
rect 10690 22000 10746 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12438 22000 12494 22800
rect 12898 22000 12954 22800
rect 13358 22000 13414 22800
rect 13818 22000 13874 22800
rect 14278 22000 14334 22800
rect 14738 22000 14794 22800
rect 15198 22000 15254 22800
rect 15658 22000 15714 22800
rect 16118 22000 16174 22800
rect 16578 22000 16634 22800
rect 17038 22000 17094 22800
rect 17498 22000 17554 22800
rect 17958 22000 18014 22800
rect 18418 22000 18474 22800
rect 18878 22000 18934 22800
rect 19338 22000 19394 22800
rect 19798 22000 19854 22800
rect 20258 22000 20314 22800
rect 20718 22000 20774 22800
rect 21178 22000 21234 22800
rect 21638 22000 21694 22800
rect 22098 22000 22154 22800
rect 22558 22000 22614 22800
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22466 0 22522 800
<< obsm2 >>
rect 314 21944 514 22545
rect 682 21944 974 22545
rect 1142 21944 1434 22545
rect 1602 21944 1894 22545
rect 2062 21944 2354 22545
rect 2522 21944 2814 22545
rect 2982 21944 3274 22545
rect 3442 21944 3734 22545
rect 3902 21944 4194 22545
rect 4362 21944 4654 22545
rect 4822 21944 5114 22545
rect 5282 21944 5574 22545
rect 5742 21944 6034 22545
rect 6202 21944 6494 22545
rect 6662 21944 6954 22545
rect 7122 21944 7414 22545
rect 7582 21944 7874 22545
rect 8042 21944 8334 22545
rect 8502 21944 8794 22545
rect 8962 21944 9254 22545
rect 9422 21944 9714 22545
rect 9882 21944 10174 22545
rect 10342 21944 10634 22545
rect 10802 21944 11094 22545
rect 11262 21944 11554 22545
rect 11722 21944 11922 22545
rect 12090 21944 12382 22545
rect 12550 21944 12842 22545
rect 13010 21944 13302 22545
rect 13470 21944 13762 22545
rect 13930 21944 14222 22545
rect 14390 21944 14682 22545
rect 14850 21944 15142 22545
rect 15310 21944 15602 22545
rect 15770 21944 16062 22545
rect 16230 21944 16522 22545
rect 16690 21944 16982 22545
rect 17150 21944 17442 22545
rect 17610 21944 17902 22545
rect 18070 21944 18362 22545
rect 18530 21944 18822 22545
rect 18990 21944 19282 22545
rect 19450 21944 19742 22545
rect 19910 21944 20202 22545
rect 20370 21944 20662 22545
rect 20830 21944 21122 22545
rect 21290 21944 21582 22545
rect 21750 21944 22042 22545
rect 22210 21944 22502 22545
rect 204 856 22612 21944
rect 314 167 606 856
rect 774 167 1066 856
rect 1234 167 1526 856
rect 1694 167 1986 856
rect 2154 167 2446 856
rect 2614 167 2906 856
rect 3074 167 3366 856
rect 3534 167 3826 856
rect 3994 167 4286 856
rect 4454 167 4746 856
rect 4914 167 5206 856
rect 5374 167 5666 856
rect 5834 167 6126 856
rect 6294 167 6586 856
rect 6754 167 7046 856
rect 7214 167 7506 856
rect 7674 167 8058 856
rect 8226 167 8518 856
rect 8686 167 8978 856
rect 9146 167 9438 856
rect 9606 167 9898 856
rect 10066 167 10358 856
rect 10526 167 10818 856
rect 10986 167 11278 856
rect 11446 167 11738 856
rect 11906 167 12198 856
rect 12366 167 12658 856
rect 12826 167 13118 856
rect 13286 167 13578 856
rect 13746 167 14038 856
rect 14206 167 14498 856
rect 14666 167 14958 856
rect 15126 167 15510 856
rect 15678 167 15970 856
rect 16138 167 16430 856
rect 16598 167 16890 856
rect 17058 167 17350 856
rect 17518 167 17810 856
rect 17978 167 18270 856
rect 18438 167 18730 856
rect 18898 167 19190 856
rect 19358 167 19650 856
rect 19818 167 20110 856
rect 20278 167 20570 856
rect 20738 167 21030 856
rect 21198 167 21490 856
rect 21658 167 21950 856
rect 22118 167 22410 856
rect 22578 167 22612 856
<< metal3 >>
rect 0 22448 800 22568
rect 0 22040 800 22160
rect 0 21496 800 21616
rect 0 21088 800 21208
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 0 19592 800 19712
rect 0 19184 800 19304
rect 0 18640 800 18760
rect 0 18232 800 18352
rect 0 17688 800 17808
rect 0 17280 800 17400
rect 22000 17144 22800 17264
rect 0 16736 800 16856
rect 0 16328 800 16448
rect 0 15784 800 15904
rect 0 15376 800 15496
rect 0 14832 800 14952
rect 0 14424 800 14544
rect 0 13880 800 14000
rect 0 13472 800 13592
rect 0 12928 800 13048
rect 0 12520 800 12640
rect 0 11976 800 12096
rect 0 11568 800 11688
rect 0 11024 800 11144
rect 0 10616 800 10736
rect 0 10072 800 10192
rect 0 9664 800 9784
rect 0 9120 800 9240
rect 0 8712 800 8832
rect 0 8168 800 8288
rect 0 7760 800 7880
rect 0 7216 800 7336
rect 0 6808 800 6928
rect 0 6264 800 6384
rect 0 5856 800 5976
rect 22000 5720 22800 5840
rect 0 5312 800 5432
rect 0 4904 800 5024
rect 0 4360 800 4480
rect 0 3952 800 4072
rect 0 3408 800 3528
rect 0 3000 800 3120
rect 0 2456 800 2576
rect 0 2048 800 2168
rect 0 1504 800 1624
rect 0 1096 800 1216
rect 0 552 800 672
rect 0 144 800 264
<< obsm3 >>
rect 880 22368 22000 22541
rect 800 22240 22000 22368
rect 880 21960 22000 22240
rect 800 21696 22000 21960
rect 880 21416 22000 21696
rect 800 21288 22000 21416
rect 880 21008 22000 21288
rect 800 20744 22000 21008
rect 880 20464 22000 20744
rect 800 20336 22000 20464
rect 880 20056 22000 20336
rect 800 19792 22000 20056
rect 880 19512 22000 19792
rect 800 19384 22000 19512
rect 880 19104 22000 19384
rect 800 18840 22000 19104
rect 880 18560 22000 18840
rect 800 18432 22000 18560
rect 880 18152 22000 18432
rect 800 17888 22000 18152
rect 880 17608 22000 17888
rect 800 17480 22000 17608
rect 880 17344 22000 17480
rect 880 17200 21920 17344
rect 800 17064 21920 17200
rect 800 16936 22000 17064
rect 880 16656 22000 16936
rect 800 16528 22000 16656
rect 880 16248 22000 16528
rect 800 15984 22000 16248
rect 880 15704 22000 15984
rect 800 15576 22000 15704
rect 880 15296 22000 15576
rect 800 15032 22000 15296
rect 880 14752 22000 15032
rect 800 14624 22000 14752
rect 880 14344 22000 14624
rect 800 14080 22000 14344
rect 880 13800 22000 14080
rect 800 13672 22000 13800
rect 880 13392 22000 13672
rect 800 13128 22000 13392
rect 880 12848 22000 13128
rect 800 12720 22000 12848
rect 880 12440 22000 12720
rect 800 12176 22000 12440
rect 880 11896 22000 12176
rect 800 11768 22000 11896
rect 880 11488 22000 11768
rect 800 11224 22000 11488
rect 880 10944 22000 11224
rect 800 10816 22000 10944
rect 880 10536 22000 10816
rect 800 10272 22000 10536
rect 880 9992 22000 10272
rect 800 9864 22000 9992
rect 880 9584 22000 9864
rect 800 9320 22000 9584
rect 880 9040 22000 9320
rect 800 8912 22000 9040
rect 880 8632 22000 8912
rect 800 8368 22000 8632
rect 880 8088 22000 8368
rect 800 7960 22000 8088
rect 880 7680 22000 7960
rect 800 7416 22000 7680
rect 880 7136 22000 7416
rect 800 7008 22000 7136
rect 880 6728 22000 7008
rect 800 6464 22000 6728
rect 880 6184 22000 6464
rect 800 6056 22000 6184
rect 880 5920 22000 6056
rect 880 5776 21920 5920
rect 800 5640 21920 5776
rect 800 5512 22000 5640
rect 880 5232 22000 5512
rect 800 5104 22000 5232
rect 880 4824 22000 5104
rect 800 4560 22000 4824
rect 880 4280 22000 4560
rect 800 4152 22000 4280
rect 880 3872 22000 4152
rect 800 3608 22000 3872
rect 880 3328 22000 3608
rect 800 3200 22000 3328
rect 880 2920 22000 3200
rect 800 2656 22000 2920
rect 880 2376 22000 2656
rect 800 2248 22000 2376
rect 880 1968 22000 2248
rect 800 1704 22000 1968
rect 880 1424 22000 1704
rect 800 1296 22000 1424
rect 880 1016 22000 1296
rect 800 752 22000 1016
rect 880 472 22000 752
rect 800 344 22000 472
rect 880 171 22000 344
<< metal4 >>
rect 4376 2128 4696 20176
rect 7808 2128 8128 20176
<< obsm4 >>
rect 4107 2048 4296 20176
rect 4776 2048 7728 20176
rect 8208 2048 18424 20176
rect 4107 1939 18424 2048
<< labels >>
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 1 nsew default input
rlabel metal2 s 662 0 718 800 6 bottom_left_grid_pin_43_
port 2 nsew default input
rlabel metal2 s 1122 0 1178 800 6 bottom_left_grid_pin_44_
port 3 nsew default input
rlabel metal2 s 1582 0 1638 800 6 bottom_left_grid_pin_45_
port 4 nsew default input
rlabel metal2 s 2042 0 2098 800 6 bottom_left_grid_pin_46_
port 5 nsew default input
rlabel metal2 s 2502 0 2558 800 6 bottom_left_grid_pin_47_
port 6 nsew default input
rlabel metal2 s 2962 0 3018 800 6 bottom_left_grid_pin_48_
port 7 nsew default input
rlabel metal2 s 3422 0 3478 800 6 bottom_left_grid_pin_49_
port 8 nsew default input
rlabel metal2 s 22466 0 22522 800 6 bottom_right_grid_pin_1_
port 9 nsew default input
rlabel metal3 s 22000 5720 22800 5840 6 ccff_head
port 10 nsew default input
rlabel metal3 s 22000 17144 22800 17264 6 ccff_tail
port 11 nsew default output
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 4904 800 5024 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 5856 800 5976 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[0]
port 32 nsew default output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[10]
port 33 nsew default output
rlabel metal3 s 0 18640 800 18760 6 chanx_left_out[11]
port 34 nsew default output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[12]
port 35 nsew default output
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[13]
port 36 nsew default output
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[14]
port 37 nsew default output
rlabel metal3 s 0 20544 800 20664 6 chanx_left_out[15]
port 38 nsew default output
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[16]
port 39 nsew default output
rlabel metal3 s 0 21496 800 21616 6 chanx_left_out[17]
port 40 nsew default output
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[18]
port 41 nsew default output
rlabel metal3 s 0 22448 800 22568 6 chanx_left_out[19]
port 42 nsew default output
rlabel metal3 s 0 13880 800 14000 6 chanx_left_out[1]
port 43 nsew default output
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[2]
port 44 nsew default output
rlabel metal3 s 0 14832 800 14952 6 chanx_left_out[3]
port 45 nsew default output
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[4]
port 46 nsew default output
rlabel metal3 s 0 15784 800 15904 6 chanx_left_out[5]
port 47 nsew default output
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[6]
port 48 nsew default output
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[7]
port 49 nsew default output
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[8]
port 50 nsew default output
rlabel metal3 s 0 17688 800 17808 6 chanx_left_out[9]
port 51 nsew default output
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[0]
port 52 nsew default input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[10]
port 53 nsew default input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[11]
port 54 nsew default input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[12]
port 55 nsew default input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[13]
port 56 nsew default input
rlabel metal2 s 10414 0 10470 800 6 chany_bottom_in[14]
port 57 nsew default input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[15]
port 58 nsew default input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[16]
port 59 nsew default input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[17]
port 60 nsew default input
rlabel metal2 s 12254 0 12310 800 6 chany_bottom_in[18]
port 61 nsew default input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_in[19]
port 62 nsew default input
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[1]
port 63 nsew default input
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_in[2]
port 64 nsew default input
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_in[3]
port 65 nsew default input
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_in[4]
port 66 nsew default input
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_in[5]
port 67 nsew default input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[6]
port 68 nsew default input
rlabel metal2 s 7102 0 7158 800 6 chany_bottom_in[7]
port 69 nsew default input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[8]
port 70 nsew default input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[9]
port 71 nsew default input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_out[0]
port 72 nsew default output
rlabel metal2 s 17866 0 17922 800 6 chany_bottom_out[10]
port 73 nsew default output
rlabel metal2 s 18326 0 18382 800 6 chany_bottom_out[11]
port 74 nsew default output
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[12]
port 75 nsew default output
rlabel metal2 s 19246 0 19302 800 6 chany_bottom_out[13]
port 76 nsew default output
rlabel metal2 s 19706 0 19762 800 6 chany_bottom_out[14]
port 77 nsew default output
rlabel metal2 s 20166 0 20222 800 6 chany_bottom_out[15]
port 78 nsew default output
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_out[16]
port 79 nsew default output
rlabel metal2 s 21086 0 21142 800 6 chany_bottom_out[17]
port 80 nsew default output
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[18]
port 81 nsew default output
rlabel metal2 s 22006 0 22062 800 6 chany_bottom_out[19]
port 82 nsew default output
rlabel metal2 s 13634 0 13690 800 6 chany_bottom_out[1]
port 83 nsew default output
rlabel metal2 s 14094 0 14150 800 6 chany_bottom_out[2]
port 84 nsew default output
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[3]
port 85 nsew default output
rlabel metal2 s 15014 0 15070 800 6 chany_bottom_out[4]
port 86 nsew default output
rlabel metal2 s 15566 0 15622 800 6 chany_bottom_out[5]
port 87 nsew default output
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[6]
port 88 nsew default output
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[7]
port 89 nsew default output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[8]
port 90 nsew default output
rlabel metal2 s 17406 0 17462 800 6 chany_bottom_out[9]
port 91 nsew default output
rlabel metal2 s 3790 22000 3846 22800 6 chany_top_in[0]
port 92 nsew default input
rlabel metal2 s 8390 22000 8446 22800 6 chany_top_in[10]
port 93 nsew default input
rlabel metal2 s 8850 22000 8906 22800 6 chany_top_in[11]
port 94 nsew default input
rlabel metal2 s 9310 22000 9366 22800 6 chany_top_in[12]
port 95 nsew default input
rlabel metal2 s 9770 22000 9826 22800 6 chany_top_in[13]
port 96 nsew default input
rlabel metal2 s 10230 22000 10286 22800 6 chany_top_in[14]
port 97 nsew default input
rlabel metal2 s 10690 22000 10746 22800 6 chany_top_in[15]
port 98 nsew default input
rlabel metal2 s 11150 22000 11206 22800 6 chany_top_in[16]
port 99 nsew default input
rlabel metal2 s 11610 22000 11666 22800 6 chany_top_in[17]
port 100 nsew default input
rlabel metal2 s 11978 22000 12034 22800 6 chany_top_in[18]
port 101 nsew default input
rlabel metal2 s 12438 22000 12494 22800 6 chany_top_in[19]
port 102 nsew default input
rlabel metal2 s 4250 22000 4306 22800 6 chany_top_in[1]
port 103 nsew default input
rlabel metal2 s 4710 22000 4766 22800 6 chany_top_in[2]
port 104 nsew default input
rlabel metal2 s 5170 22000 5226 22800 6 chany_top_in[3]
port 105 nsew default input
rlabel metal2 s 5630 22000 5686 22800 6 chany_top_in[4]
port 106 nsew default input
rlabel metal2 s 6090 22000 6146 22800 6 chany_top_in[5]
port 107 nsew default input
rlabel metal2 s 6550 22000 6606 22800 6 chany_top_in[6]
port 108 nsew default input
rlabel metal2 s 7010 22000 7066 22800 6 chany_top_in[7]
port 109 nsew default input
rlabel metal2 s 7470 22000 7526 22800 6 chany_top_in[8]
port 110 nsew default input
rlabel metal2 s 7930 22000 7986 22800 6 chany_top_in[9]
port 111 nsew default input
rlabel metal2 s 12898 22000 12954 22800 6 chany_top_out[0]
port 112 nsew default output
rlabel metal2 s 17498 22000 17554 22800 6 chany_top_out[10]
port 113 nsew default output
rlabel metal2 s 17958 22000 18014 22800 6 chany_top_out[11]
port 114 nsew default output
rlabel metal2 s 18418 22000 18474 22800 6 chany_top_out[12]
port 115 nsew default output
rlabel metal2 s 18878 22000 18934 22800 6 chany_top_out[13]
port 116 nsew default output
rlabel metal2 s 19338 22000 19394 22800 6 chany_top_out[14]
port 117 nsew default output
rlabel metal2 s 19798 22000 19854 22800 6 chany_top_out[15]
port 118 nsew default output
rlabel metal2 s 20258 22000 20314 22800 6 chany_top_out[16]
port 119 nsew default output
rlabel metal2 s 20718 22000 20774 22800 6 chany_top_out[17]
port 120 nsew default output
rlabel metal2 s 21178 22000 21234 22800 6 chany_top_out[18]
port 121 nsew default output
rlabel metal2 s 21638 22000 21694 22800 6 chany_top_out[19]
port 122 nsew default output
rlabel metal2 s 13358 22000 13414 22800 6 chany_top_out[1]
port 123 nsew default output
rlabel metal2 s 13818 22000 13874 22800 6 chany_top_out[2]
port 124 nsew default output
rlabel metal2 s 14278 22000 14334 22800 6 chany_top_out[3]
port 125 nsew default output
rlabel metal2 s 14738 22000 14794 22800 6 chany_top_out[4]
port 126 nsew default output
rlabel metal2 s 15198 22000 15254 22800 6 chany_top_out[5]
port 127 nsew default output
rlabel metal2 s 15658 22000 15714 22800 6 chany_top_out[6]
port 128 nsew default output
rlabel metal2 s 16118 22000 16174 22800 6 chany_top_out[7]
port 129 nsew default output
rlabel metal2 s 16578 22000 16634 22800 6 chany_top_out[8]
port 130 nsew default output
rlabel metal2 s 17038 22000 17094 22800 6 chany_top_out[9]
port 131 nsew default output
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 132 nsew default input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 133 nsew default input
rlabel metal3 s 0 1096 800 1216 6 left_bottom_grid_pin_36_
port 134 nsew default input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 135 nsew default input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_38_
port 136 nsew default input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 137 nsew default input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_40_
port 138 nsew default input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 139 nsew default input
rlabel metal2 s 22098 22000 22154 22800 6 prog_clk_0_N_in
port 140 nsew default input
rlabel metal2 s 202 22000 258 22800 6 top_left_grid_pin_42_
port 141 nsew default input
rlabel metal2 s 570 22000 626 22800 6 top_left_grid_pin_43_
port 142 nsew default input
rlabel metal2 s 1030 22000 1086 22800 6 top_left_grid_pin_44_
port 143 nsew default input
rlabel metal2 s 1490 22000 1546 22800 6 top_left_grid_pin_45_
port 144 nsew default input
rlabel metal2 s 1950 22000 2006 22800 6 top_left_grid_pin_46_
port 145 nsew default input
rlabel metal2 s 2410 22000 2466 22800 6 top_left_grid_pin_47_
port 146 nsew default input
rlabel metal2 s 2870 22000 2926 22800 6 top_left_grid_pin_48_
port 147 nsew default input
rlabel metal2 s 3330 22000 3386 22800 6 top_left_grid_pin_49_
port 148 nsew default input
rlabel metal2 s 22558 22000 22614 22800 6 top_right_grid_pin_1_
port 149 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 150 nsew power input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 151 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22800 22800
string LEFview TRUE
<< end >>
