* NGSPICE file created from sb_3__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

.subckt sb_3__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ bottom_right_grid_pin_13_
+ bottom_right_grid_pin_15_ bottom_right_grid_pin_1_ bottom_right_grid_pin_3_ bottom_right_grid_pin_5_
+ bottom_right_grid_pin_7_ bottom_right_grid_pin_9_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_12_ left_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ top_right_grid_pin_13_ top_right_grid_pin_15_ top_right_grid_pin_1_ top_right_grid_pin_3_
+ top_right_grid_pin_5_ top_right_grid_pin_7_ top_right_grid_pin_9_ vpwr vgnd
XFILLER_22_144 vpwr vgnd scs8hd_fill_2
XFILLER_22_177 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_85 vpwr vgnd scs8hd_fill_2
XFILLER_26_52 vpwr vgnd scs8hd_fill_2
XFILLER_26_41 vgnd vpwr scs8hd_decap_3
XFILLER_42_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_155 vpwr vgnd scs8hd_fill_2
XFILLER_13_166 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_203 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_1_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_10_147 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_73 vpwr vgnd scs8hd_fill_2
XFILLER_37_95 vpwr vgnd scs8hd_fill_2
XANTENNA__124__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_195 vgnd vpwr scs8hd_decap_12
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _208_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _189_/A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
X_131_ _121_/A _130_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_132 vgnd vpwr scs8hd_decap_4
XANTENNA__110__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_68 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _098_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_85 vgnd vpwr scs8hd_fill_1
XFILLER_34_52 vpwr vgnd scs8hd_fill_2
XFILLER_34_41 vpwr vgnd scs8hd_fill_2
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd vpwr
+ scs8hd_diode_2
X_114_ _113_/Y address[4] _090_/Y _114_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__121__B _119_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_7 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_117 vgnd vpwr scs8hd_decap_3
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_21 vpwr vgnd scs8hd_fill_2
XFILLER_20_65 vpwr vgnd scs8hd_fill_2
XANTENNA__222__A _222_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_96 vgnd vpwr scs8hd_decap_3
XFILLER_29_74 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _193_/Y mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__116__B _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_89 vgnd vpwr scs8hd_decap_3
XFILLER_13_3 vgnd vpwr scs8hd_decap_6
XFILLER_19_150 vpwr vgnd scs8hd_fill_2
XFILLER_34_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_32 vgnd vpwr scs8hd_fill_1
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XFILLER_31_167 vpwr vgnd scs8hd_fill_2
XFILLER_31_101 vpwr vgnd scs8hd_fill_2
XFILLER_16_186 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _126_/X vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_212 vpwr vgnd scs8hd_fill_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _208_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_123 vpwr vgnd scs8hd_fill_2
XFILLER_22_189 vgnd vpwr scs8hd_decap_12
XFILLER_9_105 vpwr vgnd scs8hd_fill_2
XFILLER_42_85 vgnd vpwr scs8hd_decap_8
XFILLER_13_178 vgnd vpwr scs8hd_decap_4
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_182 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _190_/Y mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_104 vgnd vpwr scs8hd_decap_6
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _224_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _102_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
X_130_ _102_/X _130_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_32 vpwr vgnd scs8hd_fill_2
XANTENNA__225__A _225_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_111 vgnd vpwr scs8hd_decap_8
XFILLER_23_87 vgnd vpwr scs8hd_decap_4
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_47 vgnd vpwr scs8hd_decap_4
XFILLER_0_58 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _134_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_67 vpwr vgnd scs8hd_fill_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_65 vgnd vpwr scs8hd_decap_6
X_113_ address[3] _113_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_15_7 vgnd vpwr scs8hd_decap_3
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_37_173 vpwr vgnd scs8hd_fill_2
XFILLER_37_162 vpwr vgnd scs8hd_fill_2
XFILLER_37_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vgnd vpwr scs8hd_decap_8
XFILLER_20_11 vgnd vpwr scs8hd_fill_1
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_20 vpwr vgnd scs8hd_fill_2
XANTENNA__132__B _130_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _192_/A mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_34_110 vpwr vgnd scs8hd_fill_2
XFILLER_19_173 vpwr vgnd scs8hd_fill_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.LATCH_1_.latch data_in _193_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_31_32 vpwr vgnd scs8hd_fill_2
XANTENNA__233__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_198 vgnd vpwr scs8hd_decap_12
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _111_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_224 vpwr vgnd scs8hd_fill_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_102 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_47 vgnd vpwr scs8hd_decap_3
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _196_/Y mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_194 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_127 vpwr vgnd scs8hd_fill_2
XFILLER_12_45 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_31 vpwr vgnd scs8hd_fill_2
XFILLER_37_20 vpwr vgnd scs8hd_fill_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_164 vpwr vgnd scs8hd_fill_2
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_38_6 vgnd vpwr scs8hd_decap_8
XANTENNA__140__B _137_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_55 vgnd vpwr scs8hd_decap_4
XANTENNA__241__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_167 vpwr vgnd scs8hd_fill_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_21 vpwr vgnd scs8hd_fill_2
XFILLER_18_55 vgnd vpwr scs8hd_decap_8
XFILLER_18_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__236__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
X_112_ _103_/A _111_/X _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_108 vgnd vpwr scs8hd_decap_3
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_89 vgnd vpwr scs8hd_decap_3
XFILLER_28_174 vgnd vpwr scs8hd_decap_4
XFILLER_6_69 vpwr vgnd scs8hd_fill_2
XFILLER_19_163 vpwr vgnd scs8hd_fill_2
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_25_177 vgnd vpwr scs8hd_decap_6
XFILLER_25_166 vpwr vgnd scs8hd_fill_2
XFILLER_25_144 vgnd vpwr scs8hd_decap_3
XFILLER_15_12 vgnd vpwr scs8hd_decap_3
XFILLER_15_67 vpwr vgnd scs8hd_fill_2
XFILLER_31_44 vgnd vpwr scs8hd_decap_3
XFILLER_16_122 vgnd vpwr scs8hd_fill_1
XFILLER_31_147 vpwr vgnd scs8hd_fill_2
XFILLER_31_136 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__B _137_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_191 vgnd vpwr scs8hd_decap_12
XFILLER_30_180 vgnd vpwr scs8hd_decap_4
XFILLER_42_76 vgnd vpwr scs8hd_decap_6
XFILLER_42_54 vgnd vpwr scs8hd_decap_8
XFILLER_42_32 vgnd vpwr scs8hd_decap_4
XFILLER_26_77 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XANTENNA__244__A _244_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__138__B _137_/X vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _111_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_68 vgnd vpwr scs8hd_fill_1
XFILLER_18_206 vgnd vpwr scs8hd_decap_8
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_54 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
Xmem_left_track_15.LATCH_0_.latch data_in _204_/A _186_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_187 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB _184_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_188_ _180_/A _163_/A _188_/C _096_/X _188_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__151__B _148_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_212 vpwr vgnd scs8hd_fill_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_4
XFILLER_34_88 vpwr vgnd scs8hd_fill_2
XFILLER_34_77 vgnd vpwr scs8hd_decap_8
X_111_ _111_/A _111_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XFILLER_38_109 vgnd vpwr scs8hd_decap_8
XANTENNA__162__A _111_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_35 vpwr vgnd scs8hd_fill_2
XANTENNA__247__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_20_7 vpwr vgnd scs8hd_fill_2
XFILLER_34_145 vgnd vpwr scs8hd_decap_8
XANTENNA__157__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_40_148 vgnd vpwr scs8hd_decap_4
XFILLER_15_24 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_12 vpwr vgnd scs8hd_fill_2
XFILLER_16_112 vpwr vgnd scs8hd_fill_2
XFILLER_16_134 vgnd vpwr scs8hd_decap_8
XFILLER_16_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_204 vgnd vpwr scs8hd_decap_4
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _191_/Y mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_148 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in _189_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_89 vgnd vpwr scs8hd_decap_3
XFILLER_26_56 vpwr vgnd scs8hd_fill_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_26_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_6
XFILLER_13_159 vgnd vpwr scs8hd_decap_4
XFILLER_21_170 vpwr vgnd scs8hd_fill_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_141 vgnd vpwr scs8hd_fill_1
XANTENNA__154__B _148_/X vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_207 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_77 vgnd vpwr scs8hd_decap_3
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XANTENNA__149__B _148_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _086_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_13 vpwr vgnd scs8hd_fill_2
XFILLER_23_79 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _180_/A _163_/A _188_/C _086_/X _187_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_191 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_9_ mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_35 vgnd vpwr scs8hd_decap_3
XFILLER_34_56 vpwr vgnd scs8hd_fill_2
XFILLER_34_45 vgnd vpwr scs8hd_decap_4
X_110_ address[1] address[2] address[0] _111_/A vgnd vpwr scs8hd_or3_4
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
X_239_ _239_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_93 vpwr vgnd scs8hd_fill_2
XFILLER_20_25 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_78 vpwr vgnd scs8hd_fill_2
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
XFILLER_20_69 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_4
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_143 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_179 vgnd vpwr scs8hd_decap_12
XFILLER_34_168 vgnd vpwr scs8hd_decap_8
XFILLER_34_135 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _162_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_79 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_223 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_216 vgnd vpwr scs8hd_decap_4
XANTENNA__168__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_127 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _190_/A mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_46 vgnd vpwr scs8hd_decap_3
XFILLER_13_138 vgnd vpwr scs8hd_decap_4
XFILLER_42_23 vgnd vpwr scs8hd_decap_8
XFILLER_9_109 vpwr vgnd scs8hd_fill_2
XFILLER_21_182 vgnd vpwr scs8hd_fill_1
XFILLER_3_39 vgnd vpwr scs8hd_decap_8
XANTENNA__170__B _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_252 vpwr vgnd scs8hd_fill_2
XFILLER_27_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _122_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_3
XFILLER_5_145 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _180_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
XFILLER_23_200 vgnd vpwr scs8hd_decap_12
XANTENNA__091__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _194_/Y mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_211 vgnd vpwr scs8hd_decap_3
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
X_186_ _180_/X _163_/A _115_/X _096_/X _186_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_91 vgnd vpwr scs8hd_fill_1
XANTENNA__176__A _172_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.LATCH_0_.latch data_in _200_/A _182_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_238_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
X_169_ _147_/A _163_/X _135_/X _165_/X _169_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_34_3 vpwr vgnd scs8hd_fill_2
XFILLER_37_177 vgnd vpwr scs8hd_decap_6
XFILLER_37_166 vgnd vpwr scs8hd_decap_4
XFILLER_1_72 vpwr vgnd scs8hd_fill_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_29_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_133 vgnd vpwr scs8hd_decap_3
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_114 vgnd vpwr scs8hd_decap_4
XFILLER_19_177 vgnd vpwr scs8hd_decap_6
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_158 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_40_106 vgnd vpwr scs8hd_decap_8
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_25_103 vpwr vgnd scs8hd_fill_2
XFILLER_40_139 vgnd vpwr scs8hd_decap_3
XFILLER_33_191 vgnd vpwr scs8hd_decap_4
XFILLER_33_180 vgnd vpwr scs8hd_decap_3
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_228 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_22_106 vgnd vpwr scs8hd_decap_8
XANTENNA__184__A _180_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_165 vgnd vpwr scs8hd_decap_8
XANTENNA__170__C _135_/X vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_37_35 vpwr vgnd scs8hd_fill_2
XFILLER_37_24 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A address[6] vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_102 vpwr vgnd scs8hd_fill_2
XFILLER_5_113 vpwr vgnd scs8hd_fill_2
XFILLER_5_135 vpwr vgnd scs8hd_fill_2
XFILLER_5_168 vpwr vgnd scs8hd_fill_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XANTENNA__181__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_83 vpwr vgnd scs8hd_fill_2
XFILLER_4_72 vpwr vgnd scs8hd_fill_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_23_212 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
X_185_ _180_/X _163_/A _115_/X _086_/X _185_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_13_70 vpwr vgnd scs8hd_fill_2
XFILLER_36_7 vpwr vgnd scs8hd_fill_2
XANTENNA__176__B _176_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_204 vgnd vpwr scs8hd_decap_8
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_25 vgnd vpwr scs8hd_decap_4
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
XFILLER_40_90 vpwr vgnd scs8hd_fill_2
X_237_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_168_ _147_/A _163_/X _188_/C _167_/X _168_/Y vgnd vpwr scs8hd_nor4_4
X_099_ _103_/A _098_/X _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_156 vgnd vpwr scs8hd_decap_3
XFILLER_37_134 vpwr vgnd scs8hd_fill_2
XFILLER_37_123 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_fill_1
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XANTENNA__097__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
XFILLER_13_9 vgnd vpwr scs8hd_fill_1
XFILLER_19_91 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XFILLER_19_167 vgnd vpwr scs8hd_decap_4
XFILLER_40_129 vgnd vpwr scs8hd_fill_1
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_6 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _188_/C vgnd vpwr scs8hd_diode_2
XANTENNA__184__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_140 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_36 vgnd vpwr scs8hd_fill_1
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_fill_1
XFILLER_16_81 vpwr vgnd scs8hd_fill_2
XANTENNA__170__D _167_/X vgnd vpwr scs8hd_diode_2
XANTENNA__179__B _176_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_28 vgnd vpwr scs8hd_decap_3
XANTENNA__089__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _189_/Y mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XANTENNA__181__C _135_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_62 vgnd vpwr scs8hd_fill_1
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_224 vgnd vpwr scs8hd_decap_12
XANTENNA__091__C _090_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_128 vpwr vgnd scs8hd_fill_2
X_184_ _180_/X _163_/X _092_/X _096_/X _184_/Y vgnd vpwr scs8hd_nor4_4
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__176__C _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_098_ _098_/A _098_/X vgnd vpwr scs8hd_buf_1
X_167_ _096_/X _167_/X vgnd vpwr scs8hd_buf_1
X_236_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__187__B _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_39 vgnd vpwr scs8hd_decap_3
XFILLER_28_113 vgnd vpwr scs8hd_decap_4
XANTENNA__097__B _087_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_50 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_127 vpwr vgnd scs8hd_fill_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_149 vpwr vgnd scs8hd_fill_2
XFILLER_25_127 vpwr vgnd scs8hd_fill_2
XFILLER_15_28 vgnd vpwr scs8hd_decap_4
XFILLER_31_49 vpwr vgnd scs8hd_fill_2
XFILLER_31_16 vgnd vpwr scs8hd_decap_3
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XFILLER_0_204 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_116 vgnd vpwr scs8hd_decap_6
XFILLER_16_149 vgnd vpwr scs8hd_decap_4
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _220_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__184__C _092_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_182 vgnd vpwr scs8hd_fill_1
XANTENNA__168__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_163 vgnd vpwr scs8hd_decap_3
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XFILLER_7_84 vpwr vgnd scs8hd_fill_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XFILLER_26_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_174 vgnd vpwr scs8hd_decap_8
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XFILLER_16_93 vgnd vpwr scs8hd_decap_6
XFILLER_8_145 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_163 vgnd vpwr scs8hd_decap_8
XFILLER_12_174 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__179__C _188_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__181__D _165_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_236 vgnd vpwr scs8hd_decap_8
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_203 vgnd vpwr scs8hd_decap_8
X_183_ _180_/X _163_/X _092_/X _086_/X _183_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_94 vpwr vgnd scs8hd_fill_2
XFILLER_1_162 vpwr vgnd scs8hd_fill_2
XANTENNA__176__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_9_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_235_ _235_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_41_7 vpwr vgnd scs8hd_fill_2
X_097_ address[1] _087_/B _096_/X _098_/A vgnd vpwr scs8hd_or3_4
X_166_ _147_/A _163_/X _188_/C _165_/X _166_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _192_/Y mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_114 vpwr vgnd scs8hd_fill_2
XFILLER_1_31 vpwr vgnd scs8hd_fill_2
XFILLER_1_42 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XANTENNA__187__C _188_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_16 vpwr vgnd scs8hd_fill_2
XFILLER_28_158 vgnd vpwr scs8hd_fill_1
XANTENNA__097__C _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_191 vgnd vpwr scs8hd_decap_12
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_202 vgnd vpwr scs8hd_decap_12
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vgnd vpwr scs8hd_decap_6
XFILLER_19_147 vgnd vpwr scs8hd_fill_1
XFILLER_27_191 vpwr vgnd scs8hd_fill_2
XFILLER_27_180 vgnd vpwr scs8hd_decap_3
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ _118_/A _148_/X _149_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_172 vpwr vgnd scs8hd_fill_2
XFILLER_33_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XFILLER_0_227 vgnd vpwr scs8hd_decap_4
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_21_83 vpwr vgnd scs8hd_fill_2
XANTENNA__184__D _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_120 vgnd vpwr scs8hd_decap_3
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_186 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _209_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_21_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_50 vgnd vpwr scs8hd_fill_1
XFILLER_32_93 vgnd vpwr scs8hd_decap_3
XFILLER_12_186 vgnd vpwr scs8hd_decap_12
XFILLER_35_256 vgnd vpwr scs8hd_decap_12
XFILLER_35_245 vgnd vpwr scs8hd_decap_3
XANTENNA__179__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_16 vgnd vpwr scs8hd_fill_1
XFILLER_5_149 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_182 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_182_ _180_/X address[5] _135_/X _167_/X _182_/Y vgnd vpwr scs8hd_nor4_4
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_7_ mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XANTENNA__100__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_13_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_165_ _086_/X _165_/X vgnd vpwr scs8hd_buf_1
XFILLER_24_61 vpwr vgnd scs8hd_fill_2
X_234_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_4
XFILLER_40_82 vgnd vpwr scs8hd_decap_8
XFILLER_40_71 vpwr vgnd scs8hd_fill_2
X_096_ address[0] _096_/X vgnd vpwr scs8hd_buf_1
XFILLER_34_7 vgnd vpwr scs8hd_decap_3
XANTENNA__187__D _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_76 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_15.LATCH_1_.latch data_in _203_/A _185_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_3_214 vgnd vpwr scs8hd_decap_12
XFILLER_19_50 vpwr vgnd scs8hd_fill_2
XFILLER_19_72 vpwr vgnd scs8hd_fill_2
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
X_148_ _147_/X _148_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_239 vgnd vpwr scs8hd_decap_8
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_114 vgnd vpwr scs8hd_decap_4
XFILLER_12_132 vpwr vgnd scs8hd_fill_2
XFILLER_12_143 vpwr vgnd scs8hd_fill_2
XFILLER_16_62 vgnd vpwr scs8hd_decap_8
XFILLER_32_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_198 vgnd vpwr scs8hd_decap_12
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_268 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_180 vgnd vpwr scs8hd_decap_3
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_117 vpwr vgnd scs8hd_fill_2
XFILLER_5_139 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_83 vpwr vgnd scs8hd_fill_2
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_194 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _180_/X address[5] _135_/X _165_/X _181_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_30 vgnd vpwr scs8hd_decap_6
XFILLER_13_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_142 vgnd vpwr scs8hd_decap_4
XFILLER_38_93 vgnd vpwr scs8hd_decap_4
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_40 vpwr vgnd scs8hd_fill_2
X_164_ _125_/X _188_/C vgnd vpwr scs8hd_buf_1
XFILLER_24_84 vgnd vpwr scs8hd_decap_6
XFILLER_24_73 vpwr vgnd scs8hd_fill_2
X_233_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
X_095_ _118_/A _103_/A _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_7 vgnd vpwr scs8hd_decap_4
XFILLER_37_138 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_226 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_171 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_fill_1
XFILLER_19_95 vpwr vgnd scs8hd_fill_2
XFILLER_19_127 vgnd vpwr scs8hd_decap_3
X_147_ _147_/A _163_/A _092_/X _147_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_182 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_fill_1
XFILLER_24_174 vgnd vpwr scs8hd_decap_12
XFILLER_24_163 vgnd vpwr scs8hd_decap_8
XFILLER_24_152 vgnd vpwr scs8hd_fill_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_152 vpwr vgnd scs8hd_fill_2
XFILLER_30_144 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_163 vpwr vgnd scs8hd_fill_2
XFILLER_15_174 vpwr vgnd scs8hd_fill_2
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _205_/A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_32_51 vpwr vgnd scs8hd_fill_2
XFILLER_8_104 vgnd vpwr scs8hd_decap_8
XFILLER_16_85 vpwr vgnd scs8hd_fill_2
XFILLER_32_84 vpwr vgnd scs8hd_fill_2
XANTENNA__103__B _102_/X vgnd vpwr scs8hd_diode_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_40_250 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_140 vgnd vpwr scs8hd_decap_12
XFILLER_4_66 vgnd vpwr scs8hd_decap_4
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
X_180_ _180_/A _180_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_132 vgnd vpwr scs8hd_decap_4
XFILLER_1_198 vpwr vgnd scs8hd_fill_2
XFILLER_1_187 vpwr vgnd scs8hd_fill_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _103_/A vgnd vpwr scs8hd_diode_2
X_232_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
X_163_ _163_/A _163_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
X_094_ _094_/A _103_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _188_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _121_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_128 vgnd vpwr scs8hd_decap_3
XFILLER_3_238 vgnd vpwr scs8hd_decap_6
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_54 vgnd vpwr scs8hd_decap_8
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XFILLER_27_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_35_84 vpwr vgnd scs8hd_fill_2
XFILLER_35_73 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vpwr vgnd scs8hd_fill_2
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
X_146_ _146_/A _163_/A vgnd vpwr scs8hd_buf_1
XANTENNA__122__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_142 vpwr vgnd scs8hd_fill_2
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
XFILLER_18_194 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _190_/Y mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_8
XFILLER_24_120 vgnd vpwr scs8hd_decap_4
Xmem_left_track_11.LATCH_1_.latch data_in _199_/A _181_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_31 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_7_88 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
X_129_ _098_/X _130_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_41 vpwr vgnd scs8hd_fill_2
XFILLER_12_112 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB _185_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_262 vgnd vpwr scs8hd_decap_12
XFILLER_32_207 vgnd vpwr scs8hd_decap_6
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
Xmem_left_track_7.LATCH_0_.latch data_in _196_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__114__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XFILLER_4_56 vgnd vpwr scs8hd_decap_6
XANTENNA__130__A _102_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XFILLER_13_43 vgnd vpwr scs8hd_fill_1
XFILLER_13_87 vgnd vpwr scs8hd_decap_4
XFILLER_13_98 vgnd vpwr scs8hd_decap_4
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_62 vgnd vpwr scs8hd_decap_8
XANTENNA__109__B _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA__125__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
X_231_ _231_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_10_210 vgnd vpwr scs8hd_decap_4
X_162_ _111_/X _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _089_/X _092_/X _094_/A vgnd vpwr scs8hd_or2_4
XFILLER_37_118 vpwr vgnd scs8hd_fill_2
XFILLER_1_35 vgnd vpwr scs8hd_decap_4
XFILLER_1_46 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_28_107 vgnd vpwr scs8hd_decap_4
XFILLER_10_44 vgnd vpwr scs8hd_decap_6
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_42_154 vgnd vpwr scs8hd_fill_1
XFILLER_35_52 vgnd vpwr scs8hd_decap_6
XFILLER_27_195 vgnd vpwr scs8hd_decap_12
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
X_145_ address[5] _146_/A vgnd vpwr scs8hd_inv_8
XANTENNA__122__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
XFILLER_33_198 vpwr vgnd scs8hd_fill_2
XFILLER_33_187 vpwr vgnd scs8hd_fill_2
XFILLER_33_176 vpwr vgnd scs8hd_fill_2
XFILLER_33_165 vpwr vgnd scs8hd_fill_2
XFILLER_33_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_110 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A _223_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_98 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_30_168 vgnd vpwr scs8hd_decap_3
XFILLER_7_67 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _111_/X vgnd vpwr scs8hd_diode_2
X_128_ _118_/A _130_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_fill_1
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_102 vpwr vgnd scs8hd_fill_2
XFILLER_21_113 vpwr vgnd scs8hd_fill_2
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_29_202 vgnd vpwr scs8hd_decap_12
XFILLER_12_124 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_109 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_274 vgnd vpwr scs8hd_fill_1
XANTENNA__114__C _090_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_241 vgnd vpwr scs8hd_decap_3
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__141__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_182 vgnd vpwr scs8hd_fill_1
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
X_230_ _230_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_24_65 vpwr vgnd scs8hd_fill_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_161_ _108_/X _162_/B _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_75 vgnd vpwr scs8hd_decap_4
X_092_ _091_/X _092_/X vgnd vpwr scs8hd_buf_1
XFILLER_37_108 vgnd vpwr scs8hd_decap_4
XANTENNA__136__A _089_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_163 vgnd vpwr scs8hd_decap_12
XFILLER_19_43 vpwr vgnd scs8hd_fill_2
XFILLER_19_54 vgnd vpwr scs8hd_decap_4
XFILLER_19_76 vpwr vgnd scs8hd_fill_2
XFILLER_42_100 vgnd vpwr scs8hd_decap_12
XFILLER_35_31 vpwr vgnd scs8hd_fill_2
XFILLER_27_130 vgnd vpwr scs8hd_decap_3
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _221_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_144_ address[6] _147_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_144 vgnd vpwr scs8hd_decap_8
XFILLER_24_133 vpwr vgnd scs8hd_fill_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_125 vgnd vpwr scs8hd_decap_4
XFILLER_30_103 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__133__B _130_/B vgnd vpwr scs8hd_diode_2
X_127_ _126_/X _130_/B vgnd vpwr scs8hd_buf_1
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_29_214 vgnd vpwr scs8hd_decap_12
XFILLER_12_147 vgnd vpwr scs8hd_decap_4
XFILLER_32_76 vpwr vgnd scs8hd_fill_2
XANTENNA__234__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XFILLER_20_180 vgnd vpwr scs8hd_decap_12
XANTENNA__144__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_32 vpwr vgnd scs8hd_fill_2
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_165 vgnd vpwr scs8hd_decap_6
XANTENNA__139__A _098_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _203_/A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XFILLER_1_146 vgnd vpwr scs8hd_fill_1
XANTENNA__125__C _090_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XANTENNA__141__B _137_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.LATCH_0_.latch data_in _192_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_091_ address[3] address[4] _090_/Y _091_/X vgnd vpwr scs8hd_or3_4
XFILLER_40_32 vgnd vpwr scs8hd_decap_4
X_160_ _121_/A _162_/B _160_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XANTENNA__242__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _135_/X vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_175 vgnd vpwr scs8hd_fill_1
XFILLER_36_120 vgnd vpwr scs8hd_decap_4
XFILLER_19_22 vgnd vpwr scs8hd_decap_4
XFILLER_19_99 vgnd vpwr scs8hd_decap_4
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_42_134 vgnd vpwr scs8hd_decap_12
XFILLER_42_112 vgnd vpwr scs8hd_fill_1
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XFILLER_27_175 vgnd vpwr scs8hd_decap_3
XANTENNA__237__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
X_143_ _111_/X _137_/X _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XFILLER_33_123 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_131 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_189 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
XFILLER_15_167 vgnd vpwr scs8hd_decap_4
XFILLER_15_178 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_126_ _089_/X _125_/X _126_/X vgnd vpwr scs8hd_or2_4
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_226 vgnd vpwr scs8hd_decap_12
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_22 vpwr vgnd scs8hd_fill_2
XFILLER_16_89 vgnd vpwr scs8hd_decap_3
XFILLER_32_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_11_170 vgnd vpwr scs8hd_fill_1
XFILLER_11_181 vpwr vgnd scs8hd_fill_2
XANTENNA__160__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
X_109_ _103_/A _108_/X _109_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_11 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA__245__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_40_221 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_133 vpwr vgnd scs8hd_fill_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_221 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _137_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_38_87 vgnd vpwr scs8hd_decap_3
XFILLER_38_32 vgnd vpwr scs8hd_decap_4
XFILLER_13_243 vgnd vpwr scs8hd_fill_1
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_39_162 vpwr vgnd scs8hd_fill_2
XFILLER_39_151 vgnd vpwr scs8hd_decap_8
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
X_090_ enable _090_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_27 vgnd vpwr scs8hd_fill_1
XANTENNA__152__B _148_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_69 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _206_/A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_27_154 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_42_146 vgnd vpwr scs8hd_decap_8
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_88 vpwr vgnd scs8hd_fill_2
XFILLER_35_77 vpwr vgnd scs8hd_fill_2
XFILLER_35_66 vpwr vgnd scs8hd_fill_2
XFILLER_27_187 vpwr vgnd scs8hd_fill_2
X_142_ _108_/X _137_/X _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _223_/A vgnd vpwr scs8hd_inv_1
XFILLER_33_146 vpwr vgnd scs8hd_fill_2
XANTENNA__147__B _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_165 vgnd vpwr scs8hd_decap_8
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vgnd vpwr scs8hd_decap_8
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_13 vpwr vgnd scs8hd_fill_2
XFILLER_21_35 vgnd vpwr scs8hd_fill_1
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_21_79 vpwr vgnd scs8hd_fill_2
XANTENNA__248__A _248_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_135 vpwr vgnd scs8hd_fill_2
X_125_ address[3] _125_/B _090_/Y _125_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_7 vgnd vpwr scs8hd_decap_3
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_205 vgnd vpwr scs8hd_decap_8
XANTENNA__158__A _098_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XFILLER_29_238 vgnd vpwr scs8hd_decap_6
XFILLER_16_46 vpwr vgnd scs8hd_fill_2
XFILLER_32_45 vgnd vpwr scs8hd_decap_4
XFILLER_12_105 vgnd vpwr scs8hd_decap_4
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _106_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
X_108_ _107_/X _108_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_120 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_fill_1
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _244_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_233 vgnd vpwr scs8hd_decap_8
XANTENNA__155__B _146_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _147_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_192 vpwr vgnd scs8hd_fill_2
XANTENNA__166__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_35 vgnd vpwr scs8hd_decap_3
XFILLER_24_13 vpwr vgnd scs8hd_fill_2
XFILLER_14_90 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_6
XFILLER_35_12 vpwr vgnd scs8hd_fill_2
XFILLER_27_100 vpwr vgnd scs8hd_fill_2
X_141_ _121_/A _137_/X _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_114 vgnd vpwr scs8hd_decap_4
XANTENNA__147__C _092_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_25 vgnd vpwr scs8hd_decap_4
XFILLER_15_103 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
X_124_ address[4] _125_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _162_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_191 vgnd vpwr scs8hd_decap_12
XANTENNA__174__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_117 vgnd vpwr scs8hd_decap_3
XANTENNA__084__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_12_128 vpwr vgnd scs8hd_fill_2
XFILLER_20_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
X_107_ address[1] address[2] _086_/A _107_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_176 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_6
XFILLER_26_209 vgnd vpwr scs8hd_decap_4
XANTENNA__169__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_231 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA__155__C _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_15 vpwr vgnd scs8hd_fill_2
XFILLER_22_201 vgnd vpwr scs8hd_decap_12
XFILLER_13_26 vpwr vgnd scs8hd_fill_2
XFILLER_38_23 vgnd vpwr scs8hd_decap_8
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_182 vgnd vpwr scs8hd_decap_4
XANTENNA__166__B _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _180_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _201_/A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_24_69 vpwr vgnd scs8hd_fill_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.INVTX1_2_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_46 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_145 vpwr vgnd scs8hd_fill_2
XFILLER_36_134 vpwr vgnd scs8hd_fill_2
XFILLER_36_112 vgnd vpwr scs8hd_fill_1
XANTENNA__177__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_58 vgnd vpwr scs8hd_fill_1
XFILLER_35_35 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_27_167 vpwr vgnd scs8hd_fill_2
X_140_ _102_/X _137_/X _140_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_3_ mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_101 vpwr vgnd scs8hd_fill_2
XFILLER_18_112 vgnd vpwr scs8hd_decap_8
XFILLER_18_145 vgnd vpwr scs8hd_decap_4
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_137 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _205_/Y mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_107 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_123_ _111_/X _119_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_11_92 vpwr vgnd scs8hd_fill_2
XFILLER_16_7 vgnd vpwr scs8hd_decap_3
XANTENNA__174__B _176_/B vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _120_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_140 vpwr vgnd scs8hd_fill_2
XFILLER_11_173 vgnd vpwr scs8hd_decap_8
XFILLER_7_155 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
X_106_ _103_/A _121_/A _106_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _180_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_71 vpwr vgnd scs8hd_fill_2
XFILLER_27_14 vgnd vpwr scs8hd_decap_3
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_91 vpwr vgnd scs8hd_fill_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_191 vgnd vpwr scs8hd_decap_4
XFILLER_3_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_79 vgnd vpwr scs8hd_decap_8
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XANTENNA__166__C _188_/C vgnd vpwr scs8hd_diode_2
XANTENNA__182__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_40_36 vgnd vpwr scs8hd_fill_1
XFILLER_6_209 vgnd vpwr scs8hd_decap_4
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_40_58 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_231 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_179 vgnd vpwr scs8hd_decap_12
XFILLER_36_124 vgnd vpwr scs8hd_fill_1
Xmem_left_track_7.LATCH_1_.latch data_in _195_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__177__B _176_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_135 vpwr vgnd scs8hd_fill_2
XFILLER_27_113 vgnd vpwr scs8hd_decap_3
XFILLER_42_116 vgnd vpwr scs8hd_decap_8
XFILLER_35_58 vgnd vpwr scs8hd_fill_1
XANTENNA__087__B _087_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_135 vgnd vpwr scs8hd_fill_1
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__188__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_2_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_24_116 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_122_ _108_/X _119_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _204_/A mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__174__C _092_/X vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_26 vgnd vpwr scs8hd_decap_3
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_163 vpwr vgnd scs8hd_fill_2
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
X_105_ _104_/X _121_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_101 vpwr vgnd scs8hd_fill_2
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XANTENNA__169__C _135_/X vgnd vpwr scs8hd_diode_2
XANTENNA__185__B _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_211 vgnd vpwr scs8hd_decap_3
XANTENNA__095__B _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vpwr vgnd scs8hd_fill_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_38_47 vgnd vpwr scs8hd_decap_12
XFILLER_13_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_0_173 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__166__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__182__C _135_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vpwr vgnd scs8hd_fill_2
XFILLER_5_51 vgnd vpwr scs8hd_decap_4
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_39_166 vgnd vpwr scs8hd_decap_12
XFILLER_39_111 vgnd vpwr scs8hd_decap_3
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_243 vgnd vpwr scs8hd_fill_1
XFILLER_39_90 vpwr vgnd scs8hd_fill_2
XFILLER_39_7 vgnd vpwr scs8hd_decap_4
XANTENNA__177__C _115_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__087__C _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_48 vpwr vgnd scs8hd_fill_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _207_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_91 vgnd vpwr scs8hd_decap_8
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__188__B _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_52 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_17 vpwr vgnd scs8hd_fill_2
XFILLER_15_139 vpwr vgnd scs8hd_fill_2
X_121_ _121_/A _119_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_8
XFILLER_12_109 vgnd vpwr scs8hd_fill_1
XFILLER_20_131 vpwr vgnd scs8hd_fill_2
XFILLER_20_142 vgnd vpwr scs8hd_decap_8
Xmem_left_track_17.LATCH_0_.latch data_in _206_/A _188_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _100_/Y address[2] _096_/X _104_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XANTENNA__169__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XANTENNA__185__C _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_40_226 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_6
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_116 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_3
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_13_215 vgnd vpwr scs8hd_decap_12
XFILLER_0_196 vgnd vpwr scs8hd_decap_4
XANTENNA__182__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_39_178 vgnd vpwr scs8hd_decap_4
XFILLER_39_134 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_17 vgnd vpwr scs8hd_decap_4
XFILLER_14_61 vgnd vpwr scs8hd_decap_8
XFILLER_30_93 vgnd vpwr scs8hd_fill_1
XFILLER_30_71 vpwr vgnd scs8hd_fill_2
XFILLER_30_60 vgnd vpwr scs8hd_decap_4
XFILLER_36_104 vpwr vgnd scs8hd_fill_2
XANTENNA__177__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_16 vgnd vpwr scs8hd_decap_4
XFILLER_19_39 vpwr vgnd scs8hd_fill_2
XFILLER_35_181 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_129 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _199_/A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_82 vpwr vgnd scs8hd_fill_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__188__C _188_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_97 vgnd vpwr scs8hd_decap_3
XFILLER_32_195 vgnd vpwr scs8hd_decap_12
XFILLER_32_184 vgnd vpwr scs8hd_decap_8
XFILLER_32_173 vgnd vpwr scs8hd_decap_8
Xmem_left_track_3.LATCH_1_.latch data_in _191_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _102_/X _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_173 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_decap_4
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_81 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
X_103_ _103_/A _102_/X _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_114 vgnd vpwr scs8hd_decap_4
XFILLER_7_136 vgnd vpwr scs8hd_decap_6
XFILLER_22_61 vpwr vgnd scs8hd_fill_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _203_/Y mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XANTENNA__185__D _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_180 vgnd vpwr scs8hd_decap_8
XFILLER_27_28 vpwr vgnd scs8hd_fill_2
XFILLER_40_238 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vpwr vgnd scs8hd_fill_2
XFILLER_3_161 vpwr vgnd scs8hd_fill_2
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_19 vgnd vpwr scs8hd_decap_4
XFILLER_13_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_0_142 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_28_71 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_40 vgnd vpwr scs8hd_fill_1
XFILLER_14_73 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_149 vgnd vpwr scs8hd_decap_4
XFILLER_36_138 vpwr vgnd scs8hd_fill_2
XFILLER_36_116 vpwr vgnd scs8hd_fill_2
XFILLER_29_190 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _100_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_19_18 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_127 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XFILLER_41_130 vpwr vgnd scs8hd_fill_2
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_3_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_8
XANTENNA__188__D _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_160 vpwr vgnd scs8hd_fill_2
XFILLER_17_171 vpwr vgnd scs8hd_fill_2
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XFILLER_23_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _207_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_41 vgnd vpwr scs8hd_fill_1
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_248_ _248_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_179_ _172_/X _176_/B _188_/C _167_/X _179_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_16_19 vpwr vgnd scs8hd_fill_2
XFILLER_32_18 vpwr vgnd scs8hd_fill_2
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
X_102_ _102_/A _102_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_159 vpwr vgnd scs8hd_fill_2
XFILLER_11_166 vgnd vpwr scs8hd_decap_4
XFILLER_22_40 vpwr vgnd scs8hd_fill_2
XFILLER_22_73 vpwr vgnd scs8hd_fill_2
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_34_203 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _202_/A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_129 vpwr vgnd scs8hd_fill_2
XFILLER_17_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _100_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_13.LATCH_0_.latch data_in _202_/A _184_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_239 vgnd vpwr scs8hd_decap_4
XFILLER_28_83 vpwr vgnd scs8hd_fill_2
XFILLER_28_61 vgnd vpwr scs8hd_decap_4
XFILLER_0_187 vgnd vpwr scs8hd_fill_1
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_98 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _154_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_18 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _206_/Y mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _225_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_84 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XANTENNA__101__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_1_ mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_7_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_4
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
X_247_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__107__A address[1] vgnd vpwr scs8hd_diode_2
X_178_ _172_/X _176_/B _188_/C _165_/X _178_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_37_234 vpwr vgnd scs8hd_fill_2
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_167 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _100_/Y address[2] _086_/X _102_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_105 vgnd vpwr scs8hd_decap_4
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_108 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_30 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XANTENNA__104__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__120__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _197_/A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_40 vpwr vgnd scs8hd_fill_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _114_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_55 vgnd vpwr scs8hd_fill_1
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_181 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _162_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_20 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XANTENNA__101__C _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_94 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_173 vpwr vgnd scs8hd_fill_2
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_3
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_6
XFILLER_2_45 vgnd vpwr scs8hd_decap_4
XANTENNA__112__B _111_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vpwr vgnd scs8hd_fill_2
XFILLER_32_143 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_10 vpwr vgnd scs8hd_fill_2
XFILLER_11_21 vpwr vgnd scs8hd_fill_2
XFILLER_36_62 vpwr vgnd scs8hd_fill_2
XFILLER_14_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
X_246_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B address[2] vgnd vpwr scs8hd_diode_2
X_177_ _172_/X _176_/B _115_/X _167_/X _177_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_42_6 vgnd vpwr scs8hd_decap_12
XANTENNA__123__A _111_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vgnd vpwr scs8hd_decap_3
XFILLER_20_113 vgnd vpwr scs8hd_fill_1
XFILLER_20_135 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
X_100_ address[1] _100_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_20 vpwr vgnd scs8hd_fill_2
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_150 vgnd vpwr scs8hd_fill_1
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
X_229_ _229_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_53 vgnd vpwr scs8hd_decap_6
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_33_85 vpwr vgnd scs8hd_fill_2
XANTENNA__104__C _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_142 vgnd vpwr scs8hd_decap_4
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _201_/Y mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _119_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_39_138 vpwr vgnd scs8hd_fill_2
XFILLER_39_116 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_193 vgnd vpwr scs8hd_decap_12
XFILLER_14_32 vgnd vpwr scs8hd_decap_8
XFILLER_30_64 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_39_62 vpwr vgnd scs8hd_fill_2
XFILLER_36_108 vgnd vpwr scs8hd_decap_4
XFILLER_29_160 vgnd vpwr scs8hd_decap_4
XANTENNA__126__A _089_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_185 vgnd vpwr scs8hd_decap_12
XFILLER_26_174 vgnd vpwr scs8hd_decap_8
XFILLER_26_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_130 vgnd vpwr scs8hd_decap_4
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_155 vgnd vpwr scs8hd_decap_12
XFILLER_41_74 vpwr vgnd scs8hd_fill_2
XFILLER_41_30 vpwr vgnd scs8hd_fill_2
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_86 vpwr vgnd scs8hd_fill_2
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XFILLER_32_122 vpwr vgnd scs8hd_fill_2
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_144 vpwr vgnd scs8hd_fill_2
XFILLER_23_177 vgnd vpwr scs8hd_decap_6
XFILLER_23_188 vgnd vpwr scs8hd_decap_12
XFILLER_11_44 vgnd vpwr scs8hd_decap_4
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
XFILLER_36_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_245_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__107__C _086_/A vgnd vpwr scs8hd_diode_2
X_176_ _172_/X _176_/B _115_/X _165_/X _176_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__123__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__224__A _224_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_fill_1
XFILLER_22_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_8
XFILLER_8_67 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _113_/Y vgnd vpwr scs8hd_diode_2
X_228_ _228_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
X_159_ _102_/X _162_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_140 vgnd vpwr scs8hd_decap_4
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_209 vgnd vpwr scs8hd_decap_12
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_198 vpwr vgnd scs8hd_fill_2
XFILLER_3_187 vpwr vgnd scs8hd_fill_2
XFILLER_3_176 vpwr vgnd scs8hd_fill_2
XFILLER_3_165 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _098_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _200_/A mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_102 vgnd vpwr scs8hd_decap_3
XFILLER_28_97 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB _186_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_79 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_44 vpwr vgnd scs8hd_fill_2
XANTENNA__232__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_150 vgnd vpwr scs8hd_decap_4
XANTENNA__126__B _125_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _108_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_134 vgnd vpwr scs8hd_fill_1
XPHY_76 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_65 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_197 vgnd vpwr scs8hd_decap_12
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_167 vgnd vpwr scs8hd_decap_12
XFILLER_41_53 vpwr vgnd scs8hd_fill_2
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _204_/Y mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_1_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_142 vgnd vpwr scs8hd_decap_4
XFILLER_17_164 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_23_134 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_244_ _244_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
X_175_ _172_/X _176_/B _092_/X _167_/X _175_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB _183_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_171 vpwr vgnd scs8hd_fill_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_28_204 vgnd vpwr scs8hd_decap_8
XFILLER_11_115 vgnd vpwr scs8hd_decap_4
XFILLER_11_159 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_227_ _227_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__134__B _125_/B vgnd vpwr scs8hd_diode_2
X_089_ address[6] address[5] _089_/X vgnd vpwr scs8hd_or2_4
X_158_ _098_/X _162_/B _158_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
XANTENNA__150__A _098_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_207 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_32 vpwr vgnd scs8hd_fill_2
XFILLER_33_10 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_111 vgnd vpwr scs8hd_decap_4
XFILLER_12_9 vgnd vpwr scs8hd_decap_8
XANTENNA__129__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_169 vpwr vgnd scs8hd_fill_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_28_87 vgnd vpwr scs8hd_decap_3
XFILLER_12_210 vgnd vpwr scs8hd_decap_4
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_58 vgnd vpwr scs8hd_decap_3
Xmem_left_track_17.LATCH_1_.latch data_in _205_/A _187_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _195_/A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_42 vpwr vgnd scs8hd_fill_2
XFILLER_30_88 vpwr vgnd scs8hd_fill_2
XFILLER_39_53 vgnd vpwr scs8hd_decap_6
XFILLER_29_184 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _137_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _219_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_209 vgnd vpwr scs8hd_decap_4
XFILLER_26_110 vgnd vpwr scs8hd_decap_6
XFILLER_41_179 vgnd vpwr scs8hd_decap_4
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_25_99 vpwr vgnd scs8hd_fill_2
XFILLER_25_66 vgnd vpwr scs8hd_decap_3
XFILLER_25_33 vpwr vgnd scs8hd_fill_2
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XANTENNA__243__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_253 vgnd vpwr scs8hd_decap_12
XFILLER_1_242 vpwr vgnd scs8hd_fill_2
XFILLER_17_110 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_3
XANTENNA__238__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_102 vgnd vpwr scs8hd_decap_3
X_243_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_14_124 vpwr vgnd scs8hd_fill_2
XFILLER_14_157 vgnd vpwr scs8hd_decap_8
XFILLER_14_168 vgnd vpwr scs8hd_decap_8
XFILLER_14_179 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
X_174_ _172_/X _176_/B _092_/X _165_/X _174_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_238 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A _147_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ _192_/A mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_11_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_15_ mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_226_ _226_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__134__C _090_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _118_/A _162_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B _148_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_197 vgnd vpwr scs8hd_decap_12
X_088_ _087_/X _118_/A vgnd vpwr scs8hd_buf_1
XFILLER_25_219 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_34 vgnd vpwr scs8hd_decap_4
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_134 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_211 vgnd vpwr scs8hd_decap_3
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_11 vgnd vpwr scs8hd_fill_1
XANTENNA__246__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_130 vgnd vpwr scs8hd_decap_4
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XFILLER_5_207 vgnd vpwr scs8hd_decap_12
XFILLER_39_21 vgnd vpwr scs8hd_decap_6
XFILLER_30_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _199_/Y mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_130 vpwr vgnd scs8hd_fill_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_5_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_177 vpwr vgnd scs8hd_fill_2
XFILLER_35_166 vpwr vgnd scs8hd_fill_2
XFILLER_25_12 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
XFILLER_41_103 vpwr vgnd scs8hd_fill_2
XFILLER_41_22 vgnd vpwr scs8hd_fill_1
XFILLER_41_11 vpwr vgnd scs8hd_fill_2
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_49 vgnd vpwr scs8hd_fill_1
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_265 vgnd vpwr scs8hd_decap_12
XFILLER_32_158 vgnd vpwr scs8hd_decap_6
XANTENNA__153__B _148_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_103 vpwr vgnd scs8hd_fill_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_23_169 vpwr vgnd scs8hd_fill_2
XFILLER_11_25 vgnd vpwr scs8hd_decap_12
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
XFILLER_36_66 vpwr vgnd scs8hd_fill_2
XFILLER_36_11 vgnd vpwr scs8hd_decap_4
X_242_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_173_ address[5] _176_/B vgnd vpwr scs8hd_buf_1
XFILLER_37_228 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _198_/A mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__164__A _125_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_140 vgnd vpwr scs8hd_decap_3
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XFILLER_13_191 vgnd vpwr scs8hd_decap_12
XFILLER_3_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_24 vgnd vpwr scs8hd_decap_4
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_225_ _225_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
X_087_ address[1] _087_/B _086_/X _087_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_110 vpwr vgnd scs8hd_fill_2
X_156_ _155_/X _162_/B vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_7 vgnd vpwr scs8hd_decap_8
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _102_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_13 vpwr vgnd scs8hd_fill_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_79 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
X_139_ _098_/X _137_/X _139_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__B _162_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XFILLER_28_67 vpwr vgnd scs8hd_fill_2
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _180_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_69 vpwr vgnd scs8hd_fill_2
XFILLER_30_35 vpwr vgnd scs8hd_fill_2
XFILLER_5_219 vgnd vpwr scs8hd_decap_12
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_145 vpwr vgnd scs8hd_fill_2
XFILLER_35_123 vpwr vgnd scs8hd_fill_2
XANTENNA__167__A _096_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_13.LATCH_1_.latch data_in _201_/A _183_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_167 vgnd vpwr scs8hd_decap_4
XFILLER_26_145 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_126 vpwr vgnd scs8hd_fill_2
XFILLER_41_34 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_78 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_126 vgnd vpwr scs8hd_decap_4
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XFILLER_17_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _099_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_126 vpwr vgnd scs8hd_fill_2
XFILLER_23_148 vpwr vgnd scs8hd_fill_2
XFILLER_11_37 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_89 vgnd vpwr scs8hd_fill_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_241_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
X_172_ _180_/A _172_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XFILLER_20_107 vgnd vpwr scs8hd_decap_6
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _202_/Y mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_36 vpwr vgnd scs8hd_fill_2
XFILLER_22_69 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A enable vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch data_in _198_/A _179_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_224_ _224_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_086_ _086_/A _086_/X vgnd vpwr scs8hd_buf_1
X_155_ address[6] _146_/A _115_/X _155_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_140 vgnd vpwr scs8hd_decap_4
XFILLER_10_151 vpwr vgnd scs8hd_fill_2
XANTENNA__159__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A _172_/X vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XANTENNA__085__A address[0] vgnd vpwr scs8hd_diode_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_207_ _207_/HI _207_/LO vgnd vpwr scs8hd_conb_1
X_138_ _118_/A _137_/X _138_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_180 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_206 vgnd vpwr scs8hd_decap_8
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_143 vpwr vgnd scs8hd_fill_2
XFILLER_14_48 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_5_ mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__183__A _180_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _248_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_41_57 vpwr vgnd scs8hd_fill_2
XANTENNA__093__A _089_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_146 vgnd vpwr scs8hd_fill_1
XFILLER_32_149 vgnd vpwr scs8hd_fill_1
XFILLER_32_105 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _193_/A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_80 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XFILLER_31_171 vpwr vgnd scs8hd_fill_2
XFILLER_36_24 vgnd vpwr scs8hd_decap_6
XANTENNA__088__A _087_/X vgnd vpwr scs8hd_diode_2
X_240_ _240_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vgnd vpwr scs8hd_decap_4
X_171_ _147_/A _180_/A vgnd vpwr scs8hd_inv_8
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _161_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_175 vgnd vpwr scs8hd_decap_8
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_119 vgnd vpwr scs8hd_fill_1
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
X_223_ _223_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
X_085_ address[0] _086_/A vgnd vpwr scs8hd_inv_8
XFILLER_6_123 vpwr vgnd scs8hd_fill_2
XFILLER_6_167 vgnd vpwr scs8hd_decap_4
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
XFILLER_10_174 vgnd vpwr scs8hd_decap_12
X_154_ _111_/X _148_/X _154_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _197_/Y mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XANTENNA__175__B _176_/B vgnd vpwr scs8hd_diode_2
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_25 vgnd vpwr scs8hd_decap_4
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ _190_/A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_148 vpwr vgnd scs8hd_fill_2
XFILLER_3_115 vgnd vpwr scs8hd_fill_1
XFILLER_30_203 vgnd vpwr scs8hd_decap_8
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
X_137_ _136_/X _137_/X vgnd vpwr scs8hd_buf_1
XFILLER_23_91 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vgnd vpwr scs8hd_fill_1
XANTENNA__186__A _180_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _222_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_36 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_79 vgnd vpwr scs8hd_decap_8
XFILLER_39_46 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XFILLER_35_103 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA__183__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_139 vpwr vgnd scs8hd_fill_2
XFILLER_34_191 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_41_47 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B _092_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_202 vgnd vpwr scs8hd_decap_8
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_139 vpwr vgnd scs8hd_fill_2
XFILLER_25_191 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _118_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__178__B _176_/B vgnd vpwr scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_14_128 vpwr vgnd scs8hd_fill_2
X_170_ _147_/A _163_/X _135_/X _167_/X _170_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_left_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_9_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_109 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_231 vgnd vpwr scs8hd_decap_12
X_222_ _222_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_102 vgnd vpwr scs8hd_decap_8
XFILLER_10_186 vgnd vpwr scs8hd_decap_12
X_153_ _108_/X _148_/X _153_/Y vgnd vpwr scs8hd_nor2_4
X_084_ address[2] _087_/B vgnd vpwr scs8hd_inv_8
XFILLER_6_146 vgnd vpwr scs8hd_decap_4
XFILLER_12_71 vpwr vgnd scs8hd_fill_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_15_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__175__C _092_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _196_/A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_201 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
Xmem_left_track_5.LATCH_0_.latch data_in _194_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_136_ _089_/X _135_/X _136_/X vgnd vpwr scs8hd_or2_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__186__B _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
X_119_ _098_/X _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vpwr vgnd scs8hd_fill_2
XFILLER_14_28 vgnd vpwr scs8hd_decap_3
XFILLER_29_156 vpwr vgnd scs8hd_fill_2
XFILLER_29_134 vgnd vpwr scs8hd_decap_3
XFILLER_20_82 vgnd vpwr scs8hd_decap_4
XFILLER_29_91 vgnd vpwr scs8hd_decap_3
XANTENNA__183__C _092_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vgnd vpwr scs8hd_decap_3
XFILLER_26_126 vpwr vgnd scs8hd_fill_2
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XFILLER_41_107 vgnd vpwr scs8hd_decap_4
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_26 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__178__C _188_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_151 vgnd vpwr scs8hd_decap_3
XFILLER_23_107 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_36_48 vgnd vpwr scs8hd_decap_8
XFILLER_14_107 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_140 vpwr vgnd scs8hd_fill_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_81 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_13_ mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_28 vgnd vpwr scs8hd_fill_1
XANTENNA__099__B _098_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_243 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
X_152_ _121_/A _148_/X _152_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_198 vgnd vpwr scs8hd_decap_12
XFILLER_37_91 vpwr vgnd scs8hd_fill_2
XFILLER_33_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA__175__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_191 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _200_/Y mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
X_135_ _134_/X _135_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__186__C _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XFILLER_9_84 vpwr vgnd scs8hd_fill_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_8
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
X_118_ _118_/A _119_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_157 vgnd vpwr scs8hd_decap_12
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XFILLER_30_39 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_179 vgnd vpwr scs8hd_decap_4
XFILLER_29_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_61 vpwr vgnd scs8hd_fill_2
XFILLER_35_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__183__D _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_149 vgnd vpwr scs8hd_decap_4
XFILLER_26_116 vgnd vpwr scs8hd_fill_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_17_138 vpwr vgnd scs8hd_fill_2
XFILLER_40_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__178__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_14_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _191_/A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
X_151_ _102_/X _148_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_144 vgnd vpwr scs8hd_fill_1
XFILLER_12_40 vpwr vgnd scs8hd_fill_2
XFILLER_12_62 vgnd vpwr scs8hd_decap_6
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_214 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
X_134_ _113_/Y _125_/B _090_/Y _134_/X vgnd vpwr scs8hd_or3_4
XFILLER_23_83 vpwr vgnd scs8hd_fill_2
XFILLER_2_184 vgnd vpwr scs8hd_decap_4
XFILLER_2_151 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__186__D _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_8
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _195_/Y mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd vpwr
+ scs8hd_diode_2
X_117_ _116_/X _119_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XFILLER_38_169 vgnd vpwr scs8hd_decap_12
XFILLER_38_147 vgnd vpwr scs8hd_decap_6
XFILLER_15_3 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.LATCH_0_.latch data_in _190_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_128 vpwr vgnd scs8hd_fill_2
XFILLER_26_106 vpwr vgnd scs8hd_fill_2
XFILLER_25_29 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_1_249 vpwr vgnd scs8hd_fill_2
XFILLER_32_109 vpwr vgnd scs8hd_fill_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XFILLER_15_84 vpwr vgnd scs8hd_fill_2
XFILLER_31_83 vgnd vpwr scs8hd_decap_3
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _192_/Y mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_197 vgnd vpwr scs8hd_decap_12
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _098_/X _148_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_123 vpwr vgnd scs8hd_fill_2
XFILLER_6_127 vpwr vgnd scs8hd_fill_2
XFILLER_10_167 vgnd vpwr scs8hd_decap_4
XFILLER_33_226 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_29 vgnd vpwr scs8hd_fill_1
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _187_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
X_133_ _111_/X _130_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_51 vpwr vgnd scs8hd_fill_2
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_9_53 vgnd vpwr scs8hd_decap_8
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _194_/A mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_40 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _089_/X _115_/X _116_/X vgnd vpwr scs8hd_or2_4
XANTENNA__105__A _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_126 vpwr vgnd scs8hd_fill_2
XFILLER_30_19 vpwr vgnd scs8hd_fill_2
XFILLER_39_17 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_107 vpwr vgnd scs8hd_fill_2
XFILLER_28_192 vgnd vpwr scs8hd_decap_12
XFILLER_28_181 vgnd vpwr scs8hd_decap_8
XFILLER_28_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_65 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_195 vgnd vpwr scs8hd_decap_12
XFILLER_25_173 vpwr vgnd scs8hd_fill_2
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_25_140 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _198_/Y mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_31_143 vpwr vgnd scs8hd_fill_2
XFILLER_31_132 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XFILLER_36_18 vgnd vpwr scs8hd_decap_4
XFILLER_22_165 vgnd vpwr scs8hd_decap_12
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_3
XFILLER_42_72 vpwr vgnd scs8hd_fill_2
XFILLER_42_50 vgnd vpwr scs8hd_fill_1
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_9_158 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vgnd vpwr scs8hd_decap_4
XFILLER_13_187 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_12_20 vgnd vpwr scs8hd_decap_8
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_50 vgnd vpwr scs8hd_decap_4
XFILLER_33_238 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _107_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
X_132_ _108_/X _130_/B _132_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_197 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__110__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_115_ _114_/X _115_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in _197_/A _178_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_29 vpwr vgnd scs8hd_fill_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vgnd vpwr scs8hd_decap_3
XFILLER_29_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_86 vgnd vpwr scs8hd_fill_1
XANTENNA__116__A _089_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_19 vgnd vpwr scs8hd_fill_1
XFILLER_1_218 vgnd vpwr scs8hd_decap_12
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_40_144 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_97 vgnd vpwr scs8hd_decap_4
XFILLER_16_163 vgnd vpwr scs8hd_decap_8
XFILLER_16_174 vgnd vpwr scs8hd_decap_12
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_200 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _209_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

