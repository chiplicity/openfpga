VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2984.540 BY 2974.160 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.510 2927.720 67.790 2930.120 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 89.720 51.880 90.320 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 105.360 2935.480 105.960 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 59.120 51.880 59.720 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 121.000 51.880 121.600 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.850 2927.720 104.130 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 214.160 51.880 214.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 229.120 2935.480 229.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.030 44.120 188.310 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 244.760 51.880 245.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 270.600 2935.480 271.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.230 44.120 243.510 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 250.130 2927.720 250.410 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 276.040 51.880 276.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 307.320 51.880 307.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 337.920 51.880 338.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 146.840 2935.480 147.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.890 44.120 299.170 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 286.470 2927.720 286.750 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 369.200 51.880 369.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 311.400 2935.480 312.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.810 2927.720 323.090 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 399.800 51.880 400.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.550 44.120 354.830 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 431.080 51.880 431.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 462.360 51.880 462.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 492.960 51.880 493.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 187.640 2935.480 188.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 524.240 51.880 524.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 352.880 2935.480 353.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 555.520 51.880 556.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.610 2927.720 359.890 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.950 2927.720 396.230 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 394.360 2935.480 394.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 435.160 2935.480 435.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 432.750 2927.720 433.030 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 586.120 51.880 586.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 469.090 2927.720 469.370 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.190 2927.720 140.470 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.890 2927.720 506.170 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.750 44.120 410.030 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 617.400 51.880 618.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.230 2927.720 542.510 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 648.680 51.880 649.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 578.570 2927.720 578.850 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 615.370 2927.720 615.650 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 651.710 2927.720 651.990 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 679.280 51.880 679.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 688.510 2927.720 688.790 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.170 44.120 77.450 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 710.560 51.880 711.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 476.640 2935.480 477.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.850 2927.720 725.130 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 741.160 51.880 741.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 517.440 2935.480 518.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 772.440 51.880 773.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 803.720 51.880 804.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 834.320 51.880 834.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 761.190 2927.720 761.470 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 865.600 51.880 866.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 151.600 51.880 152.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.410 44.120 465.690 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 521.070 44.120 521.350 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 797.990 2927.720 798.270 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 558.920 2935.480 559.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 896.880 51.880 897.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.270 44.120 576.550 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 600.400 2935.480 601.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 834.330 2927.720 834.610 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.930 44.120 632.210 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 927.480 51.880 928.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.370 44.120 132.650 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 958.760 51.880 959.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 990.040 51.880 990.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 687.590 44.120 687.870 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1020.640 51.880 1021.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.790 44.120 743.070 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 871.130 2927.720 871.410 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 798.450 44.120 798.730 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1051.920 51.880 1052.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1082.520 51.880 1083.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 641.200 2935.480 641.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 182.880 51.880 183.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.470 2927.720 907.750 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1113.800 51.880 1114.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 682.680 2935.480 683.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1145.080 51.880 1145.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 854.110 44.120 854.390 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 724.160 2935.480 724.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 764.960 2935.480 765.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.270 2927.720 944.550 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.610 2927.720 980.890 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1016.950 2927.720 1017.230 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.990 2927.720 177.270 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 806.440 2935.480 807.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 847.240 2935.480 847.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1175.680 51.880 1176.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 888.720 2935.480 889.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1053.750 2927.720 1054.030 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1090.090 2927.720 1090.370 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.330 2927.720 213.610 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.890 2927.720 1127.170 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 964.970 44.120 965.250 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1272.710 2927.720 1272.990 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1238.240 51.880 1238.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1268.840 51.880 1269.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1300.120 51.880 1300.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.630 44.120 1020.910 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1309.510 2927.720 1309.790 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1094.760 2935.480 1095.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1331.400 51.880 1332.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1136.240 2935.480 1136.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 930.200 2935.480 930.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1345.850 2927.720 1346.130 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1177.040 2935.480 1177.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.650 2927.720 1382.930 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1362.000 51.880 1362.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.830 44.120 1076.110 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.490 44.120 1131.770 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1218.520 2935.480 1219.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1393.280 51.880 1393.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.150 44.120 1187.430 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1423.880 51.880 1424.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1163.230 2927.720 1163.510 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1242.350 44.120 1242.630 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1455.160 51.880 1455.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1260.000 2935.480 1260.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1298.010 44.120 1298.290 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1300.800 2935.480 1301.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1353.670 44.120 1353.950 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.990 2927.720 1419.270 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.330 2927.720 1455.610 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1492.130 2927.720 1492.410 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1408.870 44.120 1409.150 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 971.000 2935.480 971.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1342.280 2935.480 1342.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1383.760 2935.480 1384.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1486.440 51.880 1487.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1528.470 2927.720 1528.750 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1517.040 51.880 1517.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1424.560 2935.480 1425.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1548.320 51.880 1548.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1579.600 51.880 1580.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1464.530 44.120 1464.810 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1565.270 2927.720 1565.550 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1199.570 2927.720 1199.850 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1466.040 2935.480 1466.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1520.190 44.120 1520.470 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1601.610 2927.720 1601.890 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1507.520 2935.480 1508.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1637.950 2927.720 1638.230 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1548.320 2935.480 1548.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1610.200 51.880 1610.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1589.800 2935.480 1590.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1575.390 44.120 1575.670 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1641.480 51.880 1642.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1236.370 2927.720 1236.650 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1631.050 44.120 1631.330 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1630.600 2935.480 1631.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1674.750 2927.720 1675.030 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1672.080 51.880 1672.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1672.080 2935.480 1672.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1711.090 2927.720 1711.370 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1703.360 51.880 1703.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1713.560 2935.480 1714.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1734.640 51.880 1735.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1747.890 2927.720 1748.170 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1206.960 51.880 1207.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1784.230 2927.720 1784.510 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1754.360 2935.480 1754.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1821.030 2927.720 1821.310 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.370 2927.720 1857.650 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1795.840 2935.480 1796.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1765.240 51.880 1765.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1837.320 2935.480 1837.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.710 2927.720 1893.990 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1686.250 44.120 1686.530 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1741.910 44.120 1742.190 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1012.480 2935.480 1013.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1878.120 2935.480 1878.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1930.510 2927.720 1930.790 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1966.850 2927.720 1967.130 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1797.570 44.120 1797.850 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2003.650 2927.720 2003.930 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1796.520 51.880 1797.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1827.800 51.880 1828.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1858.400 51.880 1859.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1919.600 2935.480 1920.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1960.400 2935.480 1961.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 909.310 44.120 909.590 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1852.770 44.120 1853.050 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1889.680 51.880 1890.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2001.880 2935.480 2002.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1908.430 44.120 1908.710 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1920.960 51.880 1921.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2039.990 2927.720 2040.270 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 1053.960 2935.480 1054.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2043.360 2935.480 2043.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2044.720 51.880 2045.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2019.290 44.120 2019.570 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2074.950 44.120 2075.230 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2186.270 2927.720 2186.550 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2076.000 51.880 2076.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2167.120 2935.480 2167.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2106.600 51.880 2107.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2137.880 51.880 2138.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2207.920 2935.480 2208.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2169.160 51.880 2169.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1951.560 51.880 1952.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2199.760 51.880 2200.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2249.400 2935.480 2250.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2290.200 2935.480 2290.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2231.040 51.880 2231.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2130.610 44.120 2130.890 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2185.810 44.120 2186.090 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2222.610 2927.720 2222.890 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2262.320 51.880 2262.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2331.680 2935.480 2332.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2292.920 51.880 2293.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1964.090 44.120 1964.370 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2324.200 51.880 2324.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2259.410 2927.720 2259.690 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2354.800 51.880 2355.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2295.750 2927.720 2296.030 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2332.090 2927.720 2332.370 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2386.080 51.880 2386.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2417.360 51.880 2417.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2373.160 2935.480 2373.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2241.470 44.120 2241.750 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2413.960 2935.480 2414.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2076.330 2927.720 2076.610 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2455.440 2935.480 2456.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2297.130 44.120 2297.410 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2447.960 51.880 2448.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2479.240 51.880 2479.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2352.330 44.120 2352.610 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2368.890 2927.720 2369.170 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2496.920 2935.480 2497.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2407.990 44.120 2408.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.230 2927.720 2405.510 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2537.720 2935.480 2538.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2084.160 2935.480 2084.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2442.030 2927.720 2442.310 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2478.370 2927.720 2478.650 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2514.710 2927.720 2514.990 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2551.510 2927.720 2551.790 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2510.520 51.880 2511.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2587.850 2927.720 2588.130 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2579.200 2935.480 2579.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2541.120 51.880 2541.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2463.650 44.120 2463.930 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2624.650 2927.720 2624.930 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2125.640 2935.480 2126.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2572.400 51.880 2573.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2620.000 2935.480 2620.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2661.480 2935.480 2662.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2603.680 51.880 2604.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2660.990 2927.720 2661.270 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2518.850 44.120 2519.130 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2697.790 2927.720 2698.070 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2574.510 44.120 2574.790 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2630.170 44.120 2630.450 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2702.960 2935.480 2703.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2113.130 2927.720 2113.410 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2743.760 2935.480 2744.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2685.370 44.120 2685.650 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2741.030 44.120 2741.310 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2785.240 2935.480 2785.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2826.720 2935.480 2827.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2734.130 2927.720 2734.410 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2634.280 51.880 2634.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2770.470 2927.720 2770.750 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2807.270 2927.720 2807.550 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2843.610 2927.720 2843.890 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2149.470 2927.720 2149.750 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2665.560 51.880 2666.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2696.160 51.880 2696.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2796.690 44.120 2796.970 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2727.440 51.880 2728.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2758.720 51.880 2759.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2880.410 2927.720 2880.690 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2867.520 2935.480 2868.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2933.080 2909.000 2935.480 2909.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.890 44.120 2852.170 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2916.750 2927.720 2917.030 2930.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1982.840 51.880 1983.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2907.550 44.120 2907.830 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2789.320 51.880 2789.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2820.600 51.880 2821.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2851.880 51.880 2852.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2882.480 51.880 2883.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2913.760 51.880 2914.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2013.440 51.880 2014.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2933.080 64.560 2935.480 65.160 ;
    END
  END prog_clk
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 2959.540 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 2984.540 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 99.670 58.825 2879.580 2912.615 ;
      LAYER met1 ;
        RECT 63.350 46.880 2919.810 2914.360 ;
      LAYER met2 ;
        RECT 63.370 2927.440 67.230 2927.730 ;
        RECT 68.070 2927.440 103.570 2927.730 ;
        RECT 104.410 2927.440 139.910 2927.730 ;
        RECT 140.750 2927.440 176.710 2927.730 ;
        RECT 177.550 2927.440 213.050 2927.730 ;
        RECT 213.890 2927.440 249.850 2927.730 ;
        RECT 250.690 2927.440 286.190 2927.730 ;
        RECT 287.030 2927.440 322.530 2927.730 ;
        RECT 323.370 2927.440 359.330 2927.730 ;
        RECT 360.170 2927.440 395.670 2927.730 ;
        RECT 396.510 2927.440 432.470 2927.730 ;
        RECT 433.310 2927.440 468.810 2927.730 ;
        RECT 469.650 2927.440 505.610 2927.730 ;
        RECT 506.450 2927.440 541.950 2927.730 ;
        RECT 542.790 2927.440 578.290 2927.730 ;
        RECT 579.130 2927.440 615.090 2927.730 ;
        RECT 615.930 2927.440 651.430 2927.730 ;
        RECT 652.270 2927.440 688.230 2927.730 ;
        RECT 689.070 2927.440 724.570 2927.730 ;
        RECT 725.410 2927.440 760.910 2927.730 ;
        RECT 761.750 2927.440 797.710 2927.730 ;
        RECT 798.550 2927.440 834.050 2927.730 ;
        RECT 834.890 2927.440 870.850 2927.730 ;
        RECT 871.690 2927.440 907.190 2927.730 ;
        RECT 908.030 2927.440 943.990 2927.730 ;
        RECT 944.830 2927.440 980.330 2927.730 ;
        RECT 981.170 2927.440 1016.670 2927.730 ;
        RECT 1017.510 2927.440 1053.470 2927.730 ;
        RECT 1054.310 2927.440 1089.810 2927.730 ;
        RECT 1090.650 2927.440 1126.610 2927.730 ;
        RECT 1127.450 2927.440 1162.950 2927.730 ;
        RECT 1163.790 2927.440 1199.290 2927.730 ;
        RECT 1200.130 2927.440 1236.090 2927.730 ;
        RECT 1236.930 2927.440 1272.430 2927.730 ;
        RECT 1273.270 2927.440 1309.230 2927.730 ;
        RECT 1310.070 2927.440 1345.570 2927.730 ;
        RECT 1346.410 2927.440 1382.370 2927.730 ;
        RECT 1383.210 2927.440 1418.710 2927.730 ;
        RECT 1419.550 2927.440 1455.050 2927.730 ;
        RECT 1455.890 2927.440 1491.850 2927.730 ;
        RECT 1492.690 2927.440 1528.190 2927.730 ;
        RECT 1529.030 2927.440 1564.990 2927.730 ;
        RECT 1565.830 2927.440 1601.330 2927.730 ;
        RECT 1602.170 2927.440 1637.670 2927.730 ;
        RECT 1638.510 2927.440 1674.470 2927.730 ;
        RECT 1675.310 2927.440 1710.810 2927.730 ;
        RECT 1711.650 2927.440 1747.610 2927.730 ;
        RECT 1748.450 2927.440 1783.950 2927.730 ;
        RECT 1784.790 2927.440 1820.750 2927.730 ;
        RECT 1821.590 2927.440 1857.090 2927.730 ;
        RECT 1857.930 2927.440 1893.430 2927.730 ;
        RECT 1894.270 2927.440 1930.230 2927.730 ;
        RECT 1931.070 2927.440 1966.570 2927.730 ;
        RECT 1967.410 2927.440 2003.370 2927.730 ;
        RECT 2004.210 2927.440 2039.710 2927.730 ;
        RECT 2040.550 2927.440 2076.050 2927.730 ;
        RECT 2076.890 2927.440 2112.850 2927.730 ;
        RECT 2113.690 2927.440 2149.190 2927.730 ;
        RECT 2150.030 2927.440 2185.990 2927.730 ;
        RECT 2186.830 2927.440 2222.330 2927.730 ;
        RECT 2223.170 2927.440 2259.130 2927.730 ;
        RECT 2259.970 2927.440 2295.470 2927.730 ;
        RECT 2296.310 2927.440 2331.810 2927.730 ;
        RECT 2332.650 2927.440 2368.610 2927.730 ;
        RECT 2369.450 2927.440 2404.950 2927.730 ;
        RECT 2405.790 2927.440 2441.750 2927.730 ;
        RECT 2442.590 2927.440 2478.090 2927.730 ;
        RECT 2478.930 2927.440 2514.430 2927.730 ;
        RECT 2515.270 2927.440 2551.230 2927.730 ;
        RECT 2552.070 2927.440 2587.570 2927.730 ;
        RECT 2588.410 2927.440 2624.370 2927.730 ;
        RECT 2625.210 2927.440 2660.710 2927.730 ;
        RECT 2661.550 2927.440 2697.510 2927.730 ;
        RECT 2698.350 2927.440 2733.850 2927.730 ;
        RECT 2734.690 2927.440 2770.190 2927.730 ;
        RECT 2771.030 2927.440 2806.990 2927.730 ;
        RECT 2807.830 2927.440 2843.330 2927.730 ;
        RECT 2844.170 2927.440 2880.130 2927.730 ;
        RECT 2880.970 2927.440 2916.470 2927.730 ;
        RECT 2917.310 2927.440 2919.790 2927.730 ;
        RECT 63.370 46.800 2919.790 2927.440 ;
        RECT 63.370 46.520 76.890 46.800 ;
        RECT 77.730 46.520 132.090 46.800 ;
        RECT 132.930 46.520 187.750 46.800 ;
        RECT 188.590 46.520 242.950 46.800 ;
        RECT 243.790 46.520 298.610 46.800 ;
        RECT 299.450 46.520 354.270 46.800 ;
        RECT 355.110 46.520 409.470 46.800 ;
        RECT 410.310 46.520 465.130 46.800 ;
        RECT 465.970 46.520 520.790 46.800 ;
        RECT 521.630 46.520 575.990 46.800 ;
        RECT 576.830 46.520 631.650 46.800 ;
        RECT 632.490 46.520 687.310 46.800 ;
        RECT 688.150 46.520 742.510 46.800 ;
        RECT 743.350 46.520 798.170 46.800 ;
        RECT 799.010 46.520 853.830 46.800 ;
        RECT 854.670 46.520 909.030 46.800 ;
        RECT 909.870 46.520 964.690 46.800 ;
        RECT 965.530 46.520 1020.350 46.800 ;
        RECT 1021.190 46.520 1075.550 46.800 ;
        RECT 1076.390 46.520 1131.210 46.800 ;
        RECT 1132.050 46.520 1186.870 46.800 ;
        RECT 1187.710 46.520 1242.070 46.800 ;
        RECT 1242.910 46.520 1297.730 46.800 ;
        RECT 1298.570 46.520 1353.390 46.800 ;
        RECT 1354.230 46.520 1408.590 46.800 ;
        RECT 1409.430 46.520 1464.250 46.800 ;
        RECT 1465.090 46.520 1519.910 46.800 ;
        RECT 1520.750 46.520 1575.110 46.800 ;
        RECT 1575.950 46.520 1630.770 46.800 ;
        RECT 1631.610 46.520 1685.970 46.800 ;
        RECT 1686.810 46.520 1741.630 46.800 ;
        RECT 1742.470 46.520 1797.290 46.800 ;
        RECT 1798.130 46.520 1852.490 46.800 ;
        RECT 1853.330 46.520 1908.150 46.800 ;
        RECT 1908.990 46.520 1963.810 46.800 ;
        RECT 1964.650 46.520 2019.010 46.800 ;
        RECT 2019.850 46.520 2074.670 46.800 ;
        RECT 2075.510 46.520 2130.330 46.800 ;
        RECT 2131.170 46.520 2185.530 46.800 ;
        RECT 2186.370 46.520 2241.190 46.800 ;
        RECT 2242.030 46.520 2296.850 46.800 ;
        RECT 2297.690 46.520 2352.050 46.800 ;
        RECT 2352.890 46.520 2407.710 46.800 ;
        RECT 2408.550 46.520 2463.370 46.800 ;
        RECT 2464.210 46.520 2518.570 46.800 ;
        RECT 2519.410 46.520 2574.230 46.800 ;
        RECT 2575.070 46.520 2629.890 46.800 ;
        RECT 2630.730 46.520 2685.090 46.800 ;
        RECT 2685.930 46.520 2740.750 46.800 ;
        RECT 2741.590 46.520 2796.410 46.800 ;
        RECT 2797.250 46.520 2851.610 46.800 ;
        RECT 2852.450 46.520 2907.270 46.800 ;
        RECT 2908.110 46.520 2919.790 46.800 ;
      LAYER met3 ;
        RECT 52.280 2913.360 2933.080 2914.225 ;
        RECT 51.880 2910.000 2933.080 2913.360 ;
        RECT 51.880 2908.600 2932.680 2910.000 ;
        RECT 51.880 2883.480 2933.080 2908.600 ;
        RECT 52.280 2882.080 2933.080 2883.480 ;
        RECT 51.880 2868.520 2933.080 2882.080 ;
        RECT 51.880 2867.120 2932.680 2868.520 ;
        RECT 51.880 2852.880 2933.080 2867.120 ;
        RECT 52.280 2851.480 2933.080 2852.880 ;
        RECT 51.880 2827.720 2933.080 2851.480 ;
        RECT 51.880 2826.320 2932.680 2827.720 ;
        RECT 51.880 2821.600 2933.080 2826.320 ;
        RECT 52.280 2820.200 2933.080 2821.600 ;
        RECT 51.880 2790.320 2933.080 2820.200 ;
        RECT 52.280 2788.920 2933.080 2790.320 ;
        RECT 51.880 2786.240 2933.080 2788.920 ;
        RECT 51.880 2784.840 2932.680 2786.240 ;
        RECT 51.880 2759.720 2933.080 2784.840 ;
        RECT 52.280 2758.320 2933.080 2759.720 ;
        RECT 51.880 2744.760 2933.080 2758.320 ;
        RECT 51.880 2743.360 2932.680 2744.760 ;
        RECT 51.880 2728.440 2933.080 2743.360 ;
        RECT 52.280 2727.040 2933.080 2728.440 ;
        RECT 51.880 2703.960 2933.080 2727.040 ;
        RECT 51.880 2702.560 2932.680 2703.960 ;
        RECT 51.880 2697.160 2933.080 2702.560 ;
        RECT 52.280 2695.760 2933.080 2697.160 ;
        RECT 51.880 2666.560 2933.080 2695.760 ;
        RECT 52.280 2665.160 2933.080 2666.560 ;
        RECT 51.880 2662.480 2933.080 2665.160 ;
        RECT 51.880 2661.080 2932.680 2662.480 ;
        RECT 51.880 2635.280 2933.080 2661.080 ;
        RECT 52.280 2633.880 2933.080 2635.280 ;
        RECT 51.880 2621.000 2933.080 2633.880 ;
        RECT 51.880 2619.600 2932.680 2621.000 ;
        RECT 51.880 2604.680 2933.080 2619.600 ;
        RECT 52.280 2603.280 2933.080 2604.680 ;
        RECT 51.880 2580.200 2933.080 2603.280 ;
        RECT 51.880 2578.800 2932.680 2580.200 ;
        RECT 51.880 2573.400 2933.080 2578.800 ;
        RECT 52.280 2572.000 2933.080 2573.400 ;
        RECT 51.880 2542.120 2933.080 2572.000 ;
        RECT 52.280 2540.720 2933.080 2542.120 ;
        RECT 51.880 2538.720 2933.080 2540.720 ;
        RECT 51.880 2537.320 2932.680 2538.720 ;
        RECT 51.880 2511.520 2933.080 2537.320 ;
        RECT 52.280 2510.120 2933.080 2511.520 ;
        RECT 51.880 2497.920 2933.080 2510.120 ;
        RECT 51.880 2496.520 2932.680 2497.920 ;
        RECT 51.880 2480.240 2933.080 2496.520 ;
        RECT 52.280 2478.840 2933.080 2480.240 ;
        RECT 51.880 2456.440 2933.080 2478.840 ;
        RECT 51.880 2455.040 2932.680 2456.440 ;
        RECT 51.880 2448.960 2933.080 2455.040 ;
        RECT 52.280 2447.560 2933.080 2448.960 ;
        RECT 51.880 2418.360 2933.080 2447.560 ;
        RECT 52.280 2416.960 2933.080 2418.360 ;
        RECT 51.880 2414.960 2933.080 2416.960 ;
        RECT 51.880 2413.560 2932.680 2414.960 ;
        RECT 51.880 2387.080 2933.080 2413.560 ;
        RECT 52.280 2385.680 2933.080 2387.080 ;
        RECT 51.880 2374.160 2933.080 2385.680 ;
        RECT 51.880 2372.760 2932.680 2374.160 ;
        RECT 51.880 2355.800 2933.080 2372.760 ;
        RECT 52.280 2354.400 2933.080 2355.800 ;
        RECT 51.880 2332.680 2933.080 2354.400 ;
        RECT 51.880 2331.280 2932.680 2332.680 ;
        RECT 51.880 2325.200 2933.080 2331.280 ;
        RECT 52.280 2323.800 2933.080 2325.200 ;
        RECT 51.880 2293.920 2933.080 2323.800 ;
        RECT 52.280 2292.520 2933.080 2293.920 ;
        RECT 51.880 2291.200 2933.080 2292.520 ;
        RECT 51.880 2289.800 2932.680 2291.200 ;
        RECT 51.880 2263.320 2933.080 2289.800 ;
        RECT 52.280 2261.920 2933.080 2263.320 ;
        RECT 51.880 2250.400 2933.080 2261.920 ;
        RECT 51.880 2249.000 2932.680 2250.400 ;
        RECT 51.880 2232.040 2933.080 2249.000 ;
        RECT 52.280 2230.640 2933.080 2232.040 ;
        RECT 51.880 2208.920 2933.080 2230.640 ;
        RECT 51.880 2207.520 2932.680 2208.920 ;
        RECT 51.880 2200.760 2933.080 2207.520 ;
        RECT 52.280 2199.360 2933.080 2200.760 ;
        RECT 51.880 2170.160 2933.080 2199.360 ;
        RECT 52.280 2168.760 2933.080 2170.160 ;
        RECT 51.880 2168.120 2933.080 2168.760 ;
        RECT 51.880 2166.720 2932.680 2168.120 ;
        RECT 51.880 2138.880 2933.080 2166.720 ;
        RECT 52.280 2137.480 2933.080 2138.880 ;
        RECT 51.880 2126.640 2933.080 2137.480 ;
        RECT 51.880 2125.240 2932.680 2126.640 ;
        RECT 51.880 2107.600 2933.080 2125.240 ;
        RECT 52.280 2106.200 2933.080 2107.600 ;
        RECT 51.880 2085.160 2933.080 2106.200 ;
        RECT 51.880 2083.760 2932.680 2085.160 ;
        RECT 51.880 2077.000 2933.080 2083.760 ;
        RECT 52.280 2075.600 2933.080 2077.000 ;
        RECT 51.880 2045.720 2933.080 2075.600 ;
        RECT 52.280 2044.360 2933.080 2045.720 ;
        RECT 52.280 2044.320 2932.680 2044.360 ;
        RECT 51.880 2042.960 2932.680 2044.320 ;
        RECT 51.880 2014.440 2933.080 2042.960 ;
        RECT 52.280 2013.040 2933.080 2014.440 ;
        RECT 51.880 2002.880 2933.080 2013.040 ;
        RECT 51.880 2001.480 2932.680 2002.880 ;
        RECT 51.880 1983.840 2933.080 2001.480 ;
        RECT 52.280 1982.440 2933.080 1983.840 ;
        RECT 51.880 1961.400 2933.080 1982.440 ;
        RECT 51.880 1960.000 2932.680 1961.400 ;
        RECT 51.880 1952.560 2933.080 1960.000 ;
        RECT 52.280 1951.160 2933.080 1952.560 ;
        RECT 51.880 1921.960 2933.080 1951.160 ;
        RECT 52.280 1920.600 2933.080 1921.960 ;
        RECT 52.280 1920.560 2932.680 1920.600 ;
        RECT 51.880 1919.200 2932.680 1920.560 ;
        RECT 51.880 1890.680 2933.080 1919.200 ;
        RECT 52.280 1889.280 2933.080 1890.680 ;
        RECT 51.880 1879.120 2933.080 1889.280 ;
        RECT 51.880 1877.720 2932.680 1879.120 ;
        RECT 51.880 1859.400 2933.080 1877.720 ;
        RECT 52.280 1858.000 2933.080 1859.400 ;
        RECT 51.880 1838.320 2933.080 1858.000 ;
        RECT 51.880 1836.920 2932.680 1838.320 ;
        RECT 51.880 1828.800 2933.080 1836.920 ;
        RECT 52.280 1827.400 2933.080 1828.800 ;
        RECT 51.880 1797.520 2933.080 1827.400 ;
        RECT 52.280 1796.840 2933.080 1797.520 ;
        RECT 52.280 1796.120 2932.680 1796.840 ;
        RECT 51.880 1795.440 2932.680 1796.120 ;
        RECT 51.880 1766.240 2933.080 1795.440 ;
        RECT 52.280 1764.840 2933.080 1766.240 ;
        RECT 51.880 1755.360 2933.080 1764.840 ;
        RECT 51.880 1753.960 2932.680 1755.360 ;
        RECT 51.880 1735.640 2933.080 1753.960 ;
        RECT 52.280 1734.240 2933.080 1735.640 ;
        RECT 51.880 1714.560 2933.080 1734.240 ;
        RECT 51.880 1713.160 2932.680 1714.560 ;
        RECT 51.880 1704.360 2933.080 1713.160 ;
        RECT 52.280 1702.960 2933.080 1704.360 ;
        RECT 51.880 1673.080 2933.080 1702.960 ;
        RECT 52.280 1671.680 2932.680 1673.080 ;
        RECT 51.880 1642.480 2933.080 1671.680 ;
        RECT 52.280 1641.080 2933.080 1642.480 ;
        RECT 51.880 1631.600 2933.080 1641.080 ;
        RECT 51.880 1630.200 2932.680 1631.600 ;
        RECT 51.880 1611.200 2933.080 1630.200 ;
        RECT 52.280 1609.800 2933.080 1611.200 ;
        RECT 51.880 1590.800 2933.080 1609.800 ;
        RECT 51.880 1589.400 2932.680 1590.800 ;
        RECT 51.880 1580.600 2933.080 1589.400 ;
        RECT 52.280 1579.200 2933.080 1580.600 ;
        RECT 51.880 1549.320 2933.080 1579.200 ;
        RECT 52.280 1547.920 2932.680 1549.320 ;
        RECT 51.880 1518.040 2933.080 1547.920 ;
        RECT 52.280 1516.640 2933.080 1518.040 ;
        RECT 51.880 1508.520 2933.080 1516.640 ;
        RECT 51.880 1507.120 2932.680 1508.520 ;
        RECT 51.880 1487.440 2933.080 1507.120 ;
        RECT 52.280 1486.040 2933.080 1487.440 ;
        RECT 51.880 1467.040 2933.080 1486.040 ;
        RECT 51.880 1465.640 2932.680 1467.040 ;
        RECT 51.880 1456.160 2933.080 1465.640 ;
        RECT 52.280 1454.760 2933.080 1456.160 ;
        RECT 51.880 1425.560 2933.080 1454.760 ;
        RECT 51.880 1424.880 2932.680 1425.560 ;
        RECT 52.280 1424.160 2932.680 1424.880 ;
        RECT 52.280 1423.480 2933.080 1424.160 ;
        RECT 51.880 1394.280 2933.080 1423.480 ;
        RECT 52.280 1392.880 2933.080 1394.280 ;
        RECT 51.880 1384.760 2933.080 1392.880 ;
        RECT 51.880 1383.360 2932.680 1384.760 ;
        RECT 51.880 1363.000 2933.080 1383.360 ;
        RECT 52.280 1361.600 2933.080 1363.000 ;
        RECT 51.880 1343.280 2933.080 1361.600 ;
        RECT 51.880 1341.880 2932.680 1343.280 ;
        RECT 51.880 1332.400 2933.080 1341.880 ;
        RECT 52.280 1331.000 2933.080 1332.400 ;
        RECT 51.880 1301.800 2933.080 1331.000 ;
        RECT 51.880 1301.120 2932.680 1301.800 ;
        RECT 52.280 1300.400 2932.680 1301.120 ;
        RECT 52.280 1299.720 2933.080 1300.400 ;
        RECT 51.880 1269.840 2933.080 1299.720 ;
        RECT 52.280 1268.440 2933.080 1269.840 ;
        RECT 51.880 1261.000 2933.080 1268.440 ;
        RECT 51.880 1259.600 2932.680 1261.000 ;
        RECT 51.880 1239.240 2933.080 1259.600 ;
        RECT 52.280 1237.840 2933.080 1239.240 ;
        RECT 51.880 1219.520 2933.080 1237.840 ;
        RECT 51.880 1218.120 2932.680 1219.520 ;
        RECT 51.880 1207.960 2933.080 1218.120 ;
        RECT 52.280 1206.560 2933.080 1207.960 ;
        RECT 51.880 1178.040 2933.080 1206.560 ;
        RECT 51.880 1176.680 2932.680 1178.040 ;
        RECT 52.280 1176.640 2932.680 1176.680 ;
        RECT 52.280 1175.280 2933.080 1176.640 ;
        RECT 51.880 1146.080 2933.080 1175.280 ;
        RECT 52.280 1144.680 2933.080 1146.080 ;
        RECT 51.880 1137.240 2933.080 1144.680 ;
        RECT 51.880 1135.840 2932.680 1137.240 ;
        RECT 51.880 1114.800 2933.080 1135.840 ;
        RECT 52.280 1113.400 2933.080 1114.800 ;
        RECT 51.880 1095.760 2933.080 1113.400 ;
        RECT 51.880 1094.360 2932.680 1095.760 ;
        RECT 51.880 1083.520 2933.080 1094.360 ;
        RECT 52.280 1082.120 2933.080 1083.520 ;
        RECT 51.880 1054.960 2933.080 1082.120 ;
        RECT 51.880 1053.560 2932.680 1054.960 ;
        RECT 51.880 1052.920 2933.080 1053.560 ;
        RECT 52.280 1051.520 2933.080 1052.920 ;
        RECT 51.880 1021.640 2933.080 1051.520 ;
        RECT 52.280 1020.240 2933.080 1021.640 ;
        RECT 51.880 1013.480 2933.080 1020.240 ;
        RECT 51.880 1012.080 2932.680 1013.480 ;
        RECT 51.880 991.040 2933.080 1012.080 ;
        RECT 52.280 989.640 2933.080 991.040 ;
        RECT 51.880 972.000 2933.080 989.640 ;
        RECT 51.880 970.600 2932.680 972.000 ;
        RECT 51.880 959.760 2933.080 970.600 ;
        RECT 52.280 958.360 2933.080 959.760 ;
        RECT 51.880 931.200 2933.080 958.360 ;
        RECT 51.880 929.800 2932.680 931.200 ;
        RECT 51.880 928.480 2933.080 929.800 ;
        RECT 52.280 927.080 2933.080 928.480 ;
        RECT 51.880 897.880 2933.080 927.080 ;
        RECT 52.280 896.480 2933.080 897.880 ;
        RECT 51.880 889.720 2933.080 896.480 ;
        RECT 51.880 888.320 2932.680 889.720 ;
        RECT 51.880 866.600 2933.080 888.320 ;
        RECT 52.280 865.200 2933.080 866.600 ;
        RECT 51.880 848.240 2933.080 865.200 ;
        RECT 51.880 846.840 2932.680 848.240 ;
        RECT 51.880 835.320 2933.080 846.840 ;
        RECT 52.280 833.920 2933.080 835.320 ;
        RECT 51.880 807.440 2933.080 833.920 ;
        RECT 51.880 806.040 2932.680 807.440 ;
        RECT 51.880 804.720 2933.080 806.040 ;
        RECT 52.280 803.320 2933.080 804.720 ;
        RECT 51.880 773.440 2933.080 803.320 ;
        RECT 52.280 772.040 2933.080 773.440 ;
        RECT 51.880 765.960 2933.080 772.040 ;
        RECT 51.880 764.560 2932.680 765.960 ;
        RECT 51.880 742.160 2933.080 764.560 ;
        RECT 52.280 740.760 2933.080 742.160 ;
        RECT 51.880 725.160 2933.080 740.760 ;
        RECT 51.880 723.760 2932.680 725.160 ;
        RECT 51.880 711.560 2933.080 723.760 ;
        RECT 52.280 710.160 2933.080 711.560 ;
        RECT 51.880 683.680 2933.080 710.160 ;
        RECT 51.880 682.280 2932.680 683.680 ;
        RECT 51.880 680.280 2933.080 682.280 ;
        RECT 52.280 678.880 2933.080 680.280 ;
        RECT 51.880 649.680 2933.080 678.880 ;
        RECT 52.280 648.280 2933.080 649.680 ;
        RECT 51.880 642.200 2933.080 648.280 ;
        RECT 51.880 640.800 2932.680 642.200 ;
        RECT 51.880 618.400 2933.080 640.800 ;
        RECT 52.280 617.000 2933.080 618.400 ;
        RECT 51.880 601.400 2933.080 617.000 ;
        RECT 51.880 600.000 2932.680 601.400 ;
        RECT 51.880 587.120 2933.080 600.000 ;
        RECT 52.280 585.720 2933.080 587.120 ;
        RECT 51.880 559.920 2933.080 585.720 ;
        RECT 51.880 558.520 2932.680 559.920 ;
        RECT 51.880 556.520 2933.080 558.520 ;
        RECT 52.280 555.120 2933.080 556.520 ;
        RECT 51.880 525.240 2933.080 555.120 ;
        RECT 52.280 523.840 2933.080 525.240 ;
        RECT 51.880 518.440 2933.080 523.840 ;
        RECT 51.880 517.040 2932.680 518.440 ;
        RECT 51.880 493.960 2933.080 517.040 ;
        RECT 52.280 492.560 2933.080 493.960 ;
        RECT 51.880 477.640 2933.080 492.560 ;
        RECT 51.880 476.240 2932.680 477.640 ;
        RECT 51.880 463.360 2933.080 476.240 ;
        RECT 52.280 461.960 2933.080 463.360 ;
        RECT 51.880 436.160 2933.080 461.960 ;
        RECT 51.880 434.760 2932.680 436.160 ;
        RECT 51.880 432.080 2933.080 434.760 ;
        RECT 52.280 430.680 2933.080 432.080 ;
        RECT 51.880 400.800 2933.080 430.680 ;
        RECT 52.280 399.400 2933.080 400.800 ;
        RECT 51.880 395.360 2933.080 399.400 ;
        RECT 51.880 393.960 2932.680 395.360 ;
        RECT 51.880 370.200 2933.080 393.960 ;
        RECT 52.280 368.800 2933.080 370.200 ;
        RECT 51.880 353.880 2933.080 368.800 ;
        RECT 51.880 352.480 2932.680 353.880 ;
        RECT 51.880 338.920 2933.080 352.480 ;
        RECT 52.280 337.520 2933.080 338.920 ;
        RECT 51.880 312.400 2933.080 337.520 ;
        RECT 51.880 311.000 2932.680 312.400 ;
        RECT 51.880 308.320 2933.080 311.000 ;
        RECT 52.280 306.920 2933.080 308.320 ;
        RECT 51.880 277.040 2933.080 306.920 ;
        RECT 52.280 275.640 2933.080 277.040 ;
        RECT 51.880 271.600 2933.080 275.640 ;
        RECT 51.880 270.200 2932.680 271.600 ;
        RECT 51.880 245.760 2933.080 270.200 ;
        RECT 52.280 244.360 2933.080 245.760 ;
        RECT 51.880 230.120 2933.080 244.360 ;
        RECT 51.880 228.720 2932.680 230.120 ;
        RECT 51.880 215.160 2933.080 228.720 ;
        RECT 52.280 213.760 2933.080 215.160 ;
        RECT 51.880 188.640 2933.080 213.760 ;
        RECT 51.880 187.240 2932.680 188.640 ;
        RECT 51.880 183.880 2933.080 187.240 ;
        RECT 52.280 182.480 2933.080 183.880 ;
        RECT 51.880 152.600 2933.080 182.480 ;
        RECT 52.280 151.200 2933.080 152.600 ;
        RECT 51.880 147.840 2933.080 151.200 ;
        RECT 51.880 146.440 2932.680 147.840 ;
        RECT 51.880 122.000 2933.080 146.440 ;
        RECT 52.280 120.600 2933.080 122.000 ;
        RECT 51.880 106.360 2933.080 120.600 ;
        RECT 51.880 104.960 2932.680 106.360 ;
        RECT 51.880 90.720 2933.080 104.960 ;
        RECT 52.280 89.320 2933.080 90.720 ;
        RECT 51.880 65.560 2933.080 89.320 ;
        RECT 51.880 64.160 2932.680 65.560 ;
        RECT 51.880 60.120 2933.080 64.160 ;
        RECT 52.280 59.255 2933.080 60.120 ;
      LAYER met4 ;
        RECT 0.000 0.000 2984.540 2974.160 ;
      LAYER met5 ;
        RECT 0.000 139.200 2984.540 2974.160 ;
  END
END fpga_top
END LIBRARY

