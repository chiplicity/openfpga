VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 2.400 116.920 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 1.400 140.000 2.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.960 140.000 30.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 33.360 140.000 33.960 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 36.080 140.000 36.680 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.800 140.000 39.400 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 42.200 140.000 42.800 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.920 140.000 45.520 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 47.640 140.000 48.240 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 50.360 140.000 50.960 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 53.760 140.000 54.360 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 56.480 140.000 57.080 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.120 140.000 4.720 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 9.560 140.000 10.160 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 12.960 140.000 13.560 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.680 140.000 16.280 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 21.800 140.000 22.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 24.520 140.000 25.120 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 27.240 140.000 27.840 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 59.200 140.000 59.800 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 88.440 140.000 89.040 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 91.840 140.000 92.440 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 94.560 140.000 95.160 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 97.280 140.000 97.880 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 100.000 140.000 100.600 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 103.400 140.000 104.000 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 106.120 140.000 106.720 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.840 140.000 109.440 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.960 140.000 115.560 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 62.600 140.000 63.200 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 65.320 140.000 65.920 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 68.040 140.000 68.640 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 71.440 140.000 72.040 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.160 140.000 74.760 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 76.880 140.000 77.480 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 79.600 140.000 80.200 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 83.000 140.000 83.600 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 85.720 140.000 86.320 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 137.600 4.970 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 137.600 39.010 140.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 137.600 42.230 140.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 137.600 45.910 140.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 137.600 49.130 140.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 137.600 52.810 140.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 137.600 56.030 140.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 137.600 59.710 140.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 137.600 62.930 140.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 137.600 66.150 140.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 137.600 8.190 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 137.600 11.870 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 137.600 15.090 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 137.600 18.770 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 137.600 21.990 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 137.600 25.210 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 137.600 28.890 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 137.600 32.110 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 137.600 35.790 140.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 137.600 73.050 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 137.600 107.090 140.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 137.600 110.770 140.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 137.600 113.990 140.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 137.600 117.670 140.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 137.600 120.890 140.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 137.600 124.110 140.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 137.600 127.790 140.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 137.600 131.010 140.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.410 137.600 134.690 140.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 137.600 137.910 140.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 137.600 76.730 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 137.600 79.950 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 137.600 83.170 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 137.600 86.850 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 137.600 90.070 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 137.600 93.750 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 137.600 96.970 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 137.600 100.650 140.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 137.600 103.870 140.000 ;
    END
  END chany_top_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 2.400 23.760 ;
    END
  END prog_clk
  PIN right_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 117.680 140.000 118.280 ;
    END
  END right_top_grid_pin_42_
  PIN right_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 120.400 140.000 121.000 ;
    END
  END right_top_grid_pin_43_
  PIN right_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 123.800 140.000 124.400 ;
    END
  END right_top_grid_pin_44_
  PIN right_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END right_top_grid_pin_45_
  PIN right_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END right_top_grid_pin_46_
  PIN right_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 132.640 140.000 133.240 ;
    END
  END right_top_grid_pin_47_
  PIN right_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 135.360 140.000 135.960 ;
    END
  END right_top_grid_pin_48_
  PIN right_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 138.080 140.000 138.680 ;
    END
  END right_top_grid_pin_49_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 137.600 1.750 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 5.520 2.760 134.320 128.080 ;
      LAYER met2 ;
        RECT 2.030 137.320 4.410 138.565 ;
        RECT 5.250 137.320 7.630 138.565 ;
        RECT 8.470 137.320 11.310 138.565 ;
        RECT 12.150 137.320 14.530 138.565 ;
        RECT 15.370 137.320 18.210 138.565 ;
        RECT 19.050 137.320 21.430 138.565 ;
        RECT 22.270 137.320 24.650 138.565 ;
        RECT 25.490 137.320 28.330 138.565 ;
        RECT 29.170 137.320 31.550 138.565 ;
        RECT 32.390 137.320 35.230 138.565 ;
        RECT 36.070 137.320 38.450 138.565 ;
        RECT 39.290 137.320 41.670 138.565 ;
        RECT 42.510 137.320 45.350 138.565 ;
        RECT 46.190 137.320 48.570 138.565 ;
        RECT 49.410 137.320 52.250 138.565 ;
        RECT 53.090 137.320 55.470 138.565 ;
        RECT 56.310 137.320 59.150 138.565 ;
        RECT 59.990 137.320 62.370 138.565 ;
        RECT 63.210 137.320 65.590 138.565 ;
        RECT 66.430 137.320 69.270 138.565 ;
        RECT 70.110 137.320 72.490 138.565 ;
        RECT 73.330 137.320 76.170 138.565 ;
        RECT 77.010 137.320 79.390 138.565 ;
        RECT 80.230 137.320 82.610 138.565 ;
        RECT 83.450 137.320 86.290 138.565 ;
        RECT 87.130 137.320 89.510 138.565 ;
        RECT 90.350 137.320 93.190 138.565 ;
        RECT 94.030 137.320 96.410 138.565 ;
        RECT 97.250 137.320 100.090 138.565 ;
        RECT 100.930 137.320 103.310 138.565 ;
        RECT 104.150 137.320 106.530 138.565 ;
        RECT 107.370 137.320 110.210 138.565 ;
        RECT 111.050 137.320 113.430 138.565 ;
        RECT 114.270 137.320 117.110 138.565 ;
        RECT 117.950 137.320 120.330 138.565 ;
        RECT 121.170 137.320 123.550 138.565 ;
        RECT 124.390 137.320 127.230 138.565 ;
        RECT 128.070 137.320 130.450 138.565 ;
        RECT 131.290 137.320 134.130 138.565 ;
        RECT 134.970 137.320 137.350 138.565 ;
        RECT 1.470 2.680 137.910 137.320 ;
        RECT 2.030 1.515 4.410 2.680 ;
        RECT 5.250 1.515 7.630 2.680 ;
        RECT 8.470 1.515 11.310 2.680 ;
        RECT 12.150 1.515 14.530 2.680 ;
        RECT 15.370 1.515 18.210 2.680 ;
        RECT 19.050 1.515 21.430 2.680 ;
        RECT 22.270 1.515 24.650 2.680 ;
        RECT 25.490 1.515 28.330 2.680 ;
        RECT 29.170 1.515 31.550 2.680 ;
        RECT 32.390 1.515 35.230 2.680 ;
        RECT 36.070 1.515 38.450 2.680 ;
        RECT 39.290 1.515 41.670 2.680 ;
        RECT 42.510 1.515 45.350 2.680 ;
        RECT 46.190 1.515 48.570 2.680 ;
        RECT 49.410 1.515 52.250 2.680 ;
        RECT 53.090 1.515 55.470 2.680 ;
        RECT 56.310 1.515 59.150 2.680 ;
        RECT 59.990 1.515 62.370 2.680 ;
        RECT 63.210 1.515 65.590 2.680 ;
        RECT 66.430 1.515 69.270 2.680 ;
        RECT 70.110 1.515 72.490 2.680 ;
        RECT 73.330 1.515 76.170 2.680 ;
        RECT 77.010 1.515 79.390 2.680 ;
        RECT 80.230 1.515 82.610 2.680 ;
        RECT 83.450 1.515 86.290 2.680 ;
        RECT 87.130 1.515 89.510 2.680 ;
        RECT 90.350 1.515 93.190 2.680 ;
        RECT 94.030 1.515 96.410 2.680 ;
        RECT 97.250 1.515 100.090 2.680 ;
        RECT 100.930 1.515 103.310 2.680 ;
        RECT 104.150 1.515 106.530 2.680 ;
        RECT 107.370 1.515 110.210 2.680 ;
        RECT 111.050 1.515 113.430 2.680 ;
        RECT 114.270 1.515 117.110 2.680 ;
        RECT 117.950 1.515 120.330 2.680 ;
        RECT 121.170 1.515 123.550 2.680 ;
        RECT 124.390 1.515 127.230 2.680 ;
        RECT 128.070 1.515 130.450 2.680 ;
        RECT 131.290 1.515 134.130 2.680 ;
        RECT 134.970 1.515 137.350 2.680 ;
      LAYER met3 ;
        RECT 1.445 137.680 137.200 138.545 ;
        RECT 1.445 136.360 137.935 137.680 ;
        RECT 1.445 134.960 137.200 136.360 ;
        RECT 1.445 133.640 137.935 134.960 ;
        RECT 1.445 132.240 137.200 133.640 ;
        RECT 1.445 130.240 137.935 132.240 ;
        RECT 1.445 128.840 137.200 130.240 ;
        RECT 1.445 127.520 137.935 128.840 ;
        RECT 1.445 126.120 137.200 127.520 ;
        RECT 1.445 124.800 137.935 126.120 ;
        RECT 1.445 123.400 137.200 124.800 ;
        RECT 1.445 121.400 137.935 123.400 ;
        RECT 1.445 120.000 137.200 121.400 ;
        RECT 1.445 118.680 137.935 120.000 ;
        RECT 1.445 117.320 137.200 118.680 ;
        RECT 2.800 117.280 137.200 117.320 ;
        RECT 2.800 115.960 137.935 117.280 ;
        RECT 2.800 115.920 137.200 115.960 ;
        RECT 1.445 114.560 137.200 115.920 ;
        RECT 1.445 113.240 137.935 114.560 ;
        RECT 1.445 111.840 137.200 113.240 ;
        RECT 1.445 109.840 137.935 111.840 ;
        RECT 1.445 108.440 137.200 109.840 ;
        RECT 1.445 107.120 137.935 108.440 ;
        RECT 1.445 105.720 137.200 107.120 ;
        RECT 1.445 104.400 137.935 105.720 ;
        RECT 1.445 103.000 137.200 104.400 ;
        RECT 1.445 101.000 137.935 103.000 ;
        RECT 1.445 99.600 137.200 101.000 ;
        RECT 1.445 98.280 137.935 99.600 ;
        RECT 1.445 96.880 137.200 98.280 ;
        RECT 1.445 95.560 137.935 96.880 ;
        RECT 1.445 94.160 137.200 95.560 ;
        RECT 1.445 92.840 137.935 94.160 ;
        RECT 1.445 91.440 137.200 92.840 ;
        RECT 1.445 89.440 137.935 91.440 ;
        RECT 1.445 88.040 137.200 89.440 ;
        RECT 1.445 86.720 137.935 88.040 ;
        RECT 1.445 85.320 137.200 86.720 ;
        RECT 1.445 84.000 137.935 85.320 ;
        RECT 1.445 82.600 137.200 84.000 ;
        RECT 1.445 80.600 137.935 82.600 ;
        RECT 1.445 79.200 137.200 80.600 ;
        RECT 1.445 77.880 137.935 79.200 ;
        RECT 1.445 76.480 137.200 77.880 ;
        RECT 1.445 75.160 137.935 76.480 ;
        RECT 1.445 73.760 137.200 75.160 ;
        RECT 1.445 72.440 137.935 73.760 ;
        RECT 1.445 71.040 137.200 72.440 ;
        RECT 1.445 70.400 137.935 71.040 ;
        RECT 2.800 69.040 137.935 70.400 ;
        RECT 2.800 69.000 137.200 69.040 ;
        RECT 1.445 67.640 137.200 69.000 ;
        RECT 1.445 66.320 137.935 67.640 ;
        RECT 1.445 64.920 137.200 66.320 ;
        RECT 1.445 63.600 137.935 64.920 ;
        RECT 1.445 62.200 137.200 63.600 ;
        RECT 1.445 60.200 137.935 62.200 ;
        RECT 1.445 58.800 137.200 60.200 ;
        RECT 1.445 57.480 137.935 58.800 ;
        RECT 1.445 56.080 137.200 57.480 ;
        RECT 1.445 54.760 137.935 56.080 ;
        RECT 1.445 53.360 137.200 54.760 ;
        RECT 1.445 51.360 137.935 53.360 ;
        RECT 1.445 49.960 137.200 51.360 ;
        RECT 1.445 48.640 137.935 49.960 ;
        RECT 1.445 47.240 137.200 48.640 ;
        RECT 1.445 45.920 137.935 47.240 ;
        RECT 1.445 44.520 137.200 45.920 ;
        RECT 1.445 43.200 137.935 44.520 ;
        RECT 1.445 41.800 137.200 43.200 ;
        RECT 1.445 39.800 137.935 41.800 ;
        RECT 1.445 38.400 137.200 39.800 ;
        RECT 1.445 37.080 137.935 38.400 ;
        RECT 1.445 35.680 137.200 37.080 ;
        RECT 1.445 34.360 137.935 35.680 ;
        RECT 1.445 32.960 137.200 34.360 ;
        RECT 1.445 30.960 137.935 32.960 ;
        RECT 1.445 29.560 137.200 30.960 ;
        RECT 1.445 28.240 137.935 29.560 ;
        RECT 1.445 26.840 137.200 28.240 ;
        RECT 1.445 25.520 137.935 26.840 ;
        RECT 1.445 24.160 137.200 25.520 ;
        RECT 2.800 24.120 137.200 24.160 ;
        RECT 2.800 22.800 137.935 24.120 ;
        RECT 2.800 22.760 137.200 22.800 ;
        RECT 1.445 21.400 137.200 22.760 ;
        RECT 1.445 19.400 137.935 21.400 ;
        RECT 1.445 18.000 137.200 19.400 ;
        RECT 1.445 16.680 137.935 18.000 ;
        RECT 1.445 15.280 137.200 16.680 ;
        RECT 1.445 13.960 137.935 15.280 ;
        RECT 1.445 12.560 137.200 13.960 ;
        RECT 1.445 10.560 137.935 12.560 ;
        RECT 1.445 9.160 137.200 10.560 ;
        RECT 1.445 7.840 137.935 9.160 ;
        RECT 1.445 6.440 137.200 7.840 ;
        RECT 1.445 5.120 137.935 6.440 ;
        RECT 1.445 3.720 137.200 5.120 ;
        RECT 1.445 2.400 137.935 3.720 ;
        RECT 1.445 1.535 137.200 2.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_0__1_
END LIBRARY

