magic
tech sky130A
magscale 1 2
timestamp 1604669128
<< locali >>
rect 7297 22559 7331 22729
rect 2237 16983 2271 17289
rect 6469 14943 6503 15045
rect 11897 8823 11931 9129
<< viali >>
rect 7941 25381 7975 25415
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 3065 25313 3099 25347
rect 4629 25313 4663 25347
rect 4721 25245 4755 25279
rect 4813 25245 4847 25279
rect 5825 25245 5859 25279
rect 6929 25245 6963 25279
rect 2053 25177 2087 25211
rect 1593 25109 1627 25143
rect 2421 25109 2455 25143
rect 2697 25109 2731 25143
rect 4261 25109 4295 25143
rect 7849 25109 7883 25143
rect 12909 25109 12943 25143
rect 1869 24905 1903 24939
rect 5089 24905 5123 24939
rect 2329 24837 2363 24871
rect 3065 24769 3099 24803
rect 4629 24769 4663 24803
rect 5365 24769 5399 24803
rect 6193 24769 6227 24803
rect 8309 24769 8343 24803
rect 12265 24769 12299 24803
rect 12909 24769 12943 24803
rect 13093 24769 13127 24803
rect 1409 24701 1443 24735
rect 2789 24701 2823 24735
rect 3525 24701 3559 24735
rect 4353 24701 4387 24735
rect 5549 24701 5583 24735
rect 9597 24701 9631 24735
rect 9689 24701 9723 24735
rect 3893 24633 3927 24667
rect 7665 24633 7699 24667
rect 8217 24633 8251 24667
rect 9229 24633 9263 24667
rect 9934 24633 9968 24667
rect 12817 24633 12851 24667
rect 1593 24565 1627 24599
rect 2421 24565 2455 24599
rect 2881 24565 2915 24599
rect 3985 24565 4019 24599
rect 4445 24565 4479 24599
rect 5733 24565 5767 24599
rect 7297 24565 7331 24599
rect 7757 24565 7791 24599
rect 8125 24565 8159 24599
rect 11069 24565 11103 24599
rect 11805 24565 11839 24599
rect 12449 24565 12483 24599
rect 1685 24361 1719 24395
rect 2513 24361 2547 24395
rect 7021 24361 7055 24395
rect 10149 24361 10183 24395
rect 15669 24361 15703 24395
rect 17325 24361 17359 24395
rect 21833 24361 21867 24395
rect 22937 24361 22971 24395
rect 24041 24361 24075 24395
rect 3157 24293 3191 24327
rect 3893 24293 3927 24327
rect 7941 24293 7975 24327
rect 4988 24225 5022 24259
rect 7849 24225 7883 24259
rect 10057 24225 10091 24259
rect 11345 24225 11379 24259
rect 11612 24225 11646 24259
rect 15485 24225 15519 24259
rect 17141 24225 17175 24259
rect 21649 24225 21683 24259
rect 22753 24225 22787 24259
rect 23857 24225 23891 24259
rect 2053 24157 2087 24191
rect 2605 24157 2639 24191
rect 2789 24157 2823 24191
rect 4721 24157 4755 24191
rect 8033 24157 8067 24191
rect 9505 24157 9539 24191
rect 10333 24157 10367 24191
rect 7389 24089 7423 24123
rect 2145 24021 2179 24055
rect 4353 24021 4387 24055
rect 6101 24021 6135 24055
rect 7481 24021 7515 24055
rect 9689 24021 9723 24055
rect 12725 24021 12759 24055
rect 1685 23817 1719 23851
rect 4353 23817 4387 23851
rect 4905 23817 4939 23851
rect 8125 23817 8159 23851
rect 9229 23817 9263 23851
rect 9689 23817 9723 23851
rect 11161 23817 11195 23851
rect 11713 23817 11747 23851
rect 16405 23817 16439 23851
rect 18613 23817 18647 23851
rect 19717 23817 19751 23851
rect 21925 23817 21959 23851
rect 24961 23817 24995 23851
rect 20821 23749 20855 23783
rect 23857 23749 23891 23783
rect 4813 23681 4847 23715
rect 5365 23681 5399 23715
rect 5457 23681 5491 23715
rect 7665 23681 7699 23715
rect 8677 23681 8711 23715
rect 2145 23613 2179 23647
rect 5273 23613 5307 23647
rect 7481 23613 7515 23647
rect 7573 23613 7607 23647
rect 9781 23613 9815 23647
rect 13737 23613 13771 23647
rect 16221 23613 16255 23647
rect 18429 23613 18463 23647
rect 18981 23613 19015 23647
rect 19533 23613 19567 23647
rect 20085 23613 20119 23647
rect 20637 23613 20671 23647
rect 21741 23613 21775 23647
rect 22293 23613 22327 23647
rect 23673 23613 23707 23647
rect 24593 23613 24627 23647
rect 24777 23613 24811 23647
rect 25329 23613 25363 23647
rect 2412 23545 2446 23579
rect 10026 23545 10060 23579
rect 12081 23545 12115 23579
rect 13982 23545 14016 23579
rect 21281 23545 21315 23579
rect 24225 23545 24259 23579
rect 2053 23477 2087 23511
rect 3525 23477 3559 23511
rect 5917 23477 5951 23511
rect 6561 23477 6595 23511
rect 7113 23477 7147 23511
rect 8769 23477 8803 23511
rect 12725 23477 12759 23511
rect 13553 23477 13587 23511
rect 15117 23477 15151 23511
rect 15669 23477 15703 23511
rect 16865 23477 16899 23511
rect 17233 23477 17267 23511
rect 21557 23477 21591 23511
rect 22753 23477 22787 23511
rect 2329 23273 2363 23307
rect 2973 23273 3007 23307
rect 3893 23273 3927 23307
rect 4537 23273 4571 23307
rect 6653 23273 6687 23307
rect 7021 23273 7055 23307
rect 8493 23273 8527 23307
rect 9505 23273 9539 23307
rect 13185 23273 13219 23307
rect 15485 23273 15519 23307
rect 16773 23273 16807 23307
rect 18061 23273 18095 23307
rect 21097 23273 21131 23307
rect 22385 23273 22419 23307
rect 23489 23273 23523 23307
rect 2421 23205 2455 23239
rect 10149 23205 10183 23239
rect 12072 23205 12106 23239
rect 4629 23137 4663 23171
rect 4885 23137 4919 23171
rect 7113 23137 7147 23171
rect 7380 23137 7414 23171
rect 10057 23137 10091 23171
rect 11805 23137 11839 23171
rect 15301 23137 15335 23171
rect 16589 23137 16623 23171
rect 17877 23137 17911 23171
rect 18889 23137 18923 23171
rect 20913 23137 20947 23171
rect 22201 23137 22235 23171
rect 23305 23137 23339 23171
rect 2513 23069 2547 23103
rect 10241 23069 10275 23103
rect 19073 23001 19107 23035
rect 1777 22933 1811 22967
rect 1961 22933 1995 22967
rect 6009 22933 6043 22967
rect 9689 22933 9723 22967
rect 10793 22933 10827 22967
rect 13829 22933 13863 22967
rect 4629 22729 4663 22763
rect 7113 22729 7147 22763
rect 7297 22729 7331 22763
rect 7481 22729 7515 22763
rect 9689 22729 9723 22763
rect 11437 22729 11471 22763
rect 11805 22729 11839 22763
rect 12173 22729 12207 22763
rect 14933 22729 14967 22763
rect 16313 22729 16347 22763
rect 16957 22729 16991 22763
rect 5825 22593 5859 22627
rect 6653 22593 6687 22627
rect 10425 22661 10459 22695
rect 10885 22593 10919 22627
rect 10977 22593 11011 22627
rect 2237 22525 2271 22559
rect 4261 22525 4295 22559
rect 5549 22525 5583 22559
rect 7297 22525 7331 22559
rect 7665 22525 7699 22559
rect 13553 22525 13587 22559
rect 16129 22525 16163 22559
rect 16589 22525 16623 22559
rect 2482 22457 2516 22491
rect 5089 22457 5123 22491
rect 5641 22457 5675 22491
rect 7910 22457 7944 22491
rect 12449 22457 12483 22491
rect 13369 22457 13403 22491
rect 13820 22457 13854 22491
rect 18245 22457 18279 22491
rect 1593 22389 1627 22423
rect 2053 22389 2087 22423
rect 3617 22389 3651 22423
rect 5181 22389 5215 22423
rect 6285 22389 6319 22423
rect 9045 22389 9079 22423
rect 10333 22389 10367 22423
rect 10793 22389 10827 22423
rect 13093 22389 13127 22423
rect 15577 22389 15611 22423
rect 18889 22389 18923 22423
rect 20913 22389 20947 22423
rect 22201 22389 22235 22423
rect 23305 22389 23339 22423
rect 1685 22185 1719 22219
rect 2145 22185 2179 22219
rect 4721 22185 4755 22219
rect 5457 22185 5491 22219
rect 6469 22185 6503 22219
rect 6929 22185 6963 22219
rect 7573 22185 7607 22219
rect 7941 22185 7975 22219
rect 8677 22185 8711 22219
rect 9689 22185 9723 22219
rect 10701 22185 10735 22219
rect 12909 22185 12943 22219
rect 5365 22117 5399 22151
rect 2881 22049 2915 22083
rect 6009 22049 6043 22083
rect 8125 22049 8159 22083
rect 9505 22049 9539 22083
rect 10517 22049 10551 22083
rect 11069 22049 11103 22083
rect 2237 21981 2271 22015
rect 2421 21981 2455 22015
rect 3617 21981 3651 22015
rect 4353 21981 4387 22015
rect 5549 21981 5583 22015
rect 7021 21981 7055 22015
rect 7205 21981 7239 22015
rect 11161 21981 11195 22015
rect 11345 21981 11379 22015
rect 13001 21981 13035 22015
rect 13185 21981 13219 22015
rect 1777 21845 1811 21879
rect 3341 21845 3375 21879
rect 4997 21845 5031 21879
rect 6561 21845 6595 21879
rect 8309 21845 8343 21879
rect 12541 21845 12575 21879
rect 13553 21845 13587 21879
rect 1593 21641 1627 21675
rect 2053 21641 2087 21675
rect 2421 21641 2455 21675
rect 4353 21641 4387 21675
rect 6561 21641 6595 21675
rect 6837 21641 6871 21675
rect 7849 21641 7883 21675
rect 11069 21641 11103 21675
rect 12265 21641 12299 21675
rect 12725 21641 12759 21675
rect 14565 21641 14599 21675
rect 10793 21573 10827 21607
rect 11897 21573 11931 21607
rect 3157 21505 3191 21539
rect 3709 21505 3743 21539
rect 3801 21505 3835 21539
rect 5733 21505 5767 21539
rect 7297 21505 7331 21539
rect 7481 21505 7515 21539
rect 1409 21437 1443 21471
rect 5089 21437 5123 21471
rect 5641 21437 5675 21471
rect 6285 21437 6319 21471
rect 7205 21437 7239 21471
rect 8585 21437 8619 21471
rect 8841 21437 8875 21471
rect 13185 21437 13219 21471
rect 3617 21369 3651 21403
rect 4721 21369 4755 21403
rect 13452 21369 13486 21403
rect 2789 21301 2823 21335
rect 3249 21301 3283 21335
rect 5181 21301 5215 21335
rect 5549 21301 5583 21335
rect 8401 21301 8435 21335
rect 9965 21301 9999 21335
rect 11345 21301 11379 21335
rect 13001 21301 13035 21335
rect 1593 21097 1627 21131
rect 3433 21097 3467 21131
rect 6469 21097 6503 21131
rect 10333 21097 10367 21131
rect 10793 21097 10827 21131
rect 11529 21097 11563 21131
rect 14105 21097 14139 21131
rect 1961 21029 1995 21063
rect 6828 21029 6862 21063
rect 12992 21029 13026 21063
rect 1409 20961 1443 20995
rect 2513 20961 2547 20995
rect 3157 20961 3191 20995
rect 4344 20961 4378 20995
rect 9689 20961 9723 20995
rect 4077 20893 4111 20927
rect 6561 20893 6595 20927
rect 11621 20893 11655 20927
rect 11805 20893 11839 20927
rect 12725 20893 12759 20927
rect 2697 20825 2731 20859
rect 8861 20825 8895 20859
rect 2329 20757 2363 20791
rect 3801 20757 3835 20791
rect 5457 20757 5491 20791
rect 6009 20757 6043 20791
rect 7941 20757 7975 20791
rect 8585 20757 8619 20791
rect 9873 20757 9907 20791
rect 11161 20757 11195 20791
rect 12541 20757 12575 20791
rect 1593 20553 1627 20587
rect 3341 20553 3375 20587
rect 3985 20553 4019 20587
rect 5549 20553 5583 20587
rect 6193 20553 6227 20587
rect 7297 20553 7331 20587
rect 9873 20553 9907 20587
rect 11345 20553 11379 20587
rect 11897 20553 11931 20587
rect 12449 20553 12483 20587
rect 13829 20553 13863 20587
rect 1961 20417 1995 20451
rect 4997 20417 5031 20451
rect 10241 20417 10275 20451
rect 10793 20417 10827 20451
rect 10885 20417 10919 20451
rect 12265 20417 12299 20451
rect 12909 20417 12943 20451
rect 13093 20417 13127 20451
rect 14565 20417 14599 20451
rect 15025 20417 15059 20451
rect 2228 20349 2262 20383
rect 4813 20349 4847 20383
rect 6837 20349 6871 20383
rect 7849 20349 7883 20383
rect 8116 20349 8150 20383
rect 12817 20349 12851 20383
rect 14473 20349 14507 20383
rect 4353 20281 4387 20315
rect 4905 20281 4939 20315
rect 7665 20281 7699 20315
rect 10701 20281 10735 20315
rect 13461 20281 13495 20315
rect 14381 20281 14415 20315
rect 4445 20213 4479 20247
rect 6653 20213 6687 20247
rect 7021 20213 7055 20247
rect 9229 20213 9263 20247
rect 10333 20213 10367 20247
rect 14013 20213 14047 20247
rect 2881 20009 2915 20043
rect 3433 20009 3467 20043
rect 4537 20009 4571 20043
rect 5365 20009 5399 20043
rect 5457 20009 5491 20043
rect 8033 20009 8067 20043
rect 10425 20009 10459 20043
rect 11805 20009 11839 20043
rect 12265 20009 12299 20043
rect 13737 20009 13771 20043
rect 14289 20009 14323 20043
rect 6898 19941 6932 19975
rect 1501 19873 1535 19907
rect 1768 19873 1802 19907
rect 6653 19873 6687 19907
rect 9689 19873 9723 19907
rect 11161 19873 11195 19907
rect 12357 19873 12391 19907
rect 12624 19873 12658 19907
rect 5549 19805 5583 19839
rect 11253 19805 11287 19839
rect 11437 19805 11471 19839
rect 15301 19805 15335 19839
rect 3801 19669 3835 19703
rect 4905 19669 4939 19703
rect 4997 19669 5031 19703
rect 6009 19669 6043 19703
rect 9413 19669 9447 19703
rect 9873 19669 9907 19703
rect 10793 19669 10827 19703
rect 2605 19465 2639 19499
rect 2973 19465 3007 19499
rect 3157 19465 3191 19499
rect 4721 19465 4755 19499
rect 11437 19465 11471 19499
rect 11897 19465 11931 19499
rect 13829 19465 13863 19499
rect 2237 19329 2271 19363
rect 3617 19329 3651 19363
rect 3709 19329 3743 19363
rect 5365 19329 5399 19363
rect 8125 19329 8159 19363
rect 2053 19261 2087 19295
rect 3525 19261 3559 19295
rect 5181 19261 5215 19295
rect 5273 19261 5307 19295
rect 5825 19261 5859 19295
rect 6193 19261 6227 19295
rect 7389 19261 7423 19295
rect 7941 19261 7975 19295
rect 8953 19261 8987 19295
rect 9045 19261 9079 19295
rect 12265 19261 12299 19295
rect 12449 19261 12483 19295
rect 14933 19261 14967 19295
rect 15393 19261 15427 19295
rect 8585 19193 8619 19227
rect 9290 19193 9324 19227
rect 12716 19193 12750 19227
rect 1593 19125 1627 19159
rect 1961 19125 1995 19159
rect 4353 19125 4387 19159
rect 4813 19125 4847 19159
rect 6653 19125 6687 19159
rect 7481 19125 7515 19159
rect 7849 19125 7883 19159
rect 10425 19125 10459 19159
rect 11069 19125 11103 19159
rect 15117 19125 15151 19159
rect 15945 19125 15979 19159
rect 1685 18921 1719 18955
rect 3157 18921 3191 18955
rect 3525 18921 3559 18955
rect 4721 18921 4755 18955
rect 7665 18921 7699 18955
rect 9137 18921 9171 18955
rect 10425 18921 10459 18955
rect 13001 18921 13035 18955
rect 13461 18921 13495 18955
rect 5426 18853 5460 18887
rect 9413 18853 9447 18887
rect 2145 18785 2179 18819
rect 4077 18785 4111 18819
rect 5181 18785 5215 18819
rect 7205 18785 7239 18819
rect 8033 18785 8067 18819
rect 8125 18785 8159 18819
rect 10784 18785 10818 18819
rect 13369 18785 13403 18819
rect 2237 18717 2271 18751
rect 2329 18717 2363 18751
rect 7573 18717 7607 18751
rect 8309 18717 8343 18751
rect 10517 18717 10551 18751
rect 13553 18717 13587 18751
rect 15301 18717 15335 18751
rect 16313 18717 16347 18751
rect 12909 18649 12943 18683
rect 1777 18581 1811 18615
rect 2881 18581 2915 18615
rect 4261 18581 4295 18615
rect 5089 18581 5123 18615
rect 6561 18581 6595 18615
rect 9965 18581 9999 18615
rect 11897 18581 11931 18615
rect 12541 18581 12575 18615
rect 14013 18581 14047 18615
rect 2053 18377 2087 18411
rect 3617 18377 3651 18411
rect 4261 18377 4295 18411
rect 8217 18377 8251 18411
rect 9321 18377 9355 18411
rect 11437 18377 11471 18411
rect 12265 18377 12299 18411
rect 13369 18377 13403 18411
rect 23857 18377 23891 18411
rect 8861 18309 8895 18343
rect 13093 18309 13127 18343
rect 14933 18309 14967 18343
rect 2237 18241 2271 18275
rect 5365 18241 5399 18275
rect 6101 18241 6135 18275
rect 9137 18241 9171 18275
rect 9781 18241 9815 18275
rect 9965 18241 9999 18275
rect 12449 18241 12483 18275
rect 2504 18173 2538 18207
rect 4629 18173 4663 18207
rect 5089 18173 5123 18207
rect 5825 18173 5859 18207
rect 6653 18173 6687 18207
rect 6837 18173 6871 18207
rect 9689 18173 9723 18207
rect 10885 18173 10919 18207
rect 11805 18173 11839 18207
rect 13553 18173 13587 18207
rect 16313 18173 16347 18207
rect 23673 18173 23707 18207
rect 24133 18173 24167 18207
rect 5181 18105 5215 18139
rect 7082 18105 7116 18139
rect 13820 18105 13854 18139
rect 1685 18037 1719 18071
rect 4721 18037 4755 18071
rect 10609 18037 10643 18071
rect 11069 18037 11103 18071
rect 16497 18037 16531 18071
rect 16957 18037 16991 18071
rect 2237 17833 2271 17867
rect 2329 17833 2363 17867
rect 3341 17833 3375 17867
rect 3801 17833 3835 17867
rect 4261 17833 4295 17867
rect 6101 17833 6135 17867
rect 7665 17833 7699 17867
rect 9413 17833 9447 17867
rect 11989 17833 12023 17867
rect 13461 17833 13495 17867
rect 17049 17833 17083 17867
rect 7573 17765 7607 17799
rect 8769 17765 8803 17799
rect 10854 17765 10888 17799
rect 1869 17697 1903 17731
rect 2697 17697 2731 17731
rect 4721 17697 4755 17731
rect 4988 17697 5022 17731
rect 8033 17697 8067 17731
rect 10609 17697 10643 17731
rect 15669 17697 15703 17731
rect 16865 17697 16899 17731
rect 17877 17697 17911 17731
rect 2789 17629 2823 17663
rect 2973 17629 3007 17663
rect 8125 17629 8159 17663
rect 8309 17629 8343 17663
rect 13553 17629 13587 17663
rect 13737 17629 13771 17663
rect 14105 17629 14139 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 13093 17561 13127 17595
rect 15301 17561 15335 17595
rect 6929 17493 6963 17527
rect 9873 17493 9907 17527
rect 12909 17493 12943 17527
rect 18061 17493 18095 17527
rect 1593 17289 1627 17323
rect 2053 17289 2087 17323
rect 2237 17289 2271 17323
rect 2329 17289 2363 17323
rect 3525 17289 3559 17323
rect 4261 17289 4295 17323
rect 5365 17289 5399 17323
rect 7573 17289 7607 17323
rect 10517 17289 10551 17323
rect 11437 17289 11471 17323
rect 12265 17289 12299 17323
rect 14197 17289 14231 17323
rect 14841 17289 14875 17323
rect 17233 17289 17267 17323
rect 18521 17289 18555 17323
rect 1409 17085 1443 17119
rect 2697 17221 2731 17255
rect 3157 17221 3191 17255
rect 8585 17221 8619 17255
rect 8953 17221 8987 17255
rect 4169 17153 4203 17187
rect 4813 17153 4847 17187
rect 7113 17153 7147 17187
rect 8125 17153 8159 17187
rect 9137 17153 9171 17187
rect 18061 17153 18095 17187
rect 2513 17085 2547 17119
rect 4629 17085 4663 17119
rect 7941 17085 7975 17119
rect 8033 17085 8067 17119
rect 9404 17085 9438 17119
rect 12817 17085 12851 17119
rect 15301 17085 15335 17119
rect 15568 17085 15602 17119
rect 6009 17017 6043 17051
rect 13084 17017 13118 17051
rect 2237 16949 2271 16983
rect 4721 16949 4755 16983
rect 5641 16949 5675 16983
rect 6561 16949 6595 16983
rect 7389 16949 7423 16983
rect 11161 16949 11195 16983
rect 12725 16949 12759 16983
rect 15209 16949 15243 16983
rect 16681 16949 16715 16983
rect 1409 16745 1443 16779
rect 2329 16745 2363 16779
rect 2881 16745 2915 16779
rect 3893 16745 3927 16779
rect 5181 16745 5215 16779
rect 8033 16745 8067 16779
rect 9229 16745 9263 16779
rect 9873 16745 9907 16779
rect 11437 16745 11471 16779
rect 11989 16745 12023 16779
rect 13829 16745 13863 16779
rect 14289 16745 14323 16779
rect 15485 16745 15519 16779
rect 15853 16745 15887 16779
rect 16129 16745 16163 16779
rect 19349 16745 19383 16779
rect 4353 16677 4387 16711
rect 8493 16677 8527 16711
rect 13461 16677 13495 16711
rect 15117 16677 15151 16711
rect 16926 16677 16960 16711
rect 2789 16609 2823 16643
rect 5089 16609 5123 16643
rect 6377 16609 6411 16643
rect 6837 16609 6871 16643
rect 7757 16609 7791 16643
rect 8401 16609 8435 16643
rect 9689 16609 9723 16643
rect 10609 16609 10643 16643
rect 10793 16609 10827 16643
rect 12357 16609 12391 16643
rect 14105 16609 14139 16643
rect 15301 16609 15335 16643
rect 19165 16609 19199 16643
rect 3065 16541 3099 16575
rect 5365 16541 5399 16575
rect 6929 16541 6963 16575
rect 7021 16541 7055 16575
rect 8677 16541 8711 16575
rect 12449 16541 12483 16575
rect 12633 16541 12667 16575
rect 16681 16541 16715 16575
rect 4721 16473 4755 16507
rect 1961 16405 1995 16439
rect 2421 16405 2455 16439
rect 3525 16405 3559 16439
rect 5733 16405 5767 16439
rect 6469 16405 6503 16439
rect 10241 16405 10275 16439
rect 10977 16405 11011 16439
rect 13185 16405 13219 16439
rect 18061 16405 18095 16439
rect 4721 16201 4755 16235
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 8033 16201 8067 16235
rect 9045 16201 9079 16235
rect 11621 16201 11655 16235
rect 13093 16201 13127 16235
rect 16037 16201 16071 16235
rect 19901 16201 19935 16235
rect 20637 16201 20671 16235
rect 4445 16133 4479 16167
rect 6929 16133 6963 16167
rect 2237 16065 2271 16099
rect 3893 16065 3927 16099
rect 5733 16065 5767 16099
rect 7389 16065 7423 16099
rect 7573 16065 7607 16099
rect 8493 16065 8527 16099
rect 9413 16065 9447 16099
rect 10057 16065 10091 16099
rect 13553 16065 13587 16099
rect 13737 16065 13771 16099
rect 2053 15997 2087 16031
rect 3617 15997 3651 16031
rect 5641 15997 5675 16031
rect 11069 15997 11103 16031
rect 14657 15997 14691 16031
rect 14924 15997 14958 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 19073 15997 19107 16031
rect 19533 15997 19567 16031
rect 20453 15997 20487 16031
rect 21005 15997 21039 16031
rect 2145 15929 2179 15963
rect 3157 15929 3191 15963
rect 9873 15929 9907 15963
rect 13461 15929 13495 15963
rect 14197 15929 14231 15963
rect 1685 15861 1719 15895
rect 2789 15861 2823 15895
rect 3249 15861 3283 15895
rect 3709 15861 3743 15895
rect 5181 15861 5215 15895
rect 5549 15861 5583 15895
rect 7297 15861 7331 15895
rect 9505 15861 9539 15895
rect 9965 15861 9999 15895
rect 10609 15861 10643 15895
rect 10977 15861 11011 15895
rect 11253 15861 11287 15895
rect 12081 15861 12115 15895
rect 12909 15861 12943 15895
rect 14565 15861 14599 15895
rect 16681 15861 16715 15895
rect 17049 15861 17083 15895
rect 18245 15861 18279 15895
rect 19257 15861 19291 15895
rect 2881 15657 2915 15691
rect 3525 15657 3559 15691
rect 4629 15657 4663 15691
rect 7205 15657 7239 15691
rect 8309 15657 8343 15691
rect 8953 15657 8987 15691
rect 12357 15657 12391 15691
rect 14197 15657 14231 15691
rect 14749 15657 14783 15691
rect 15485 15657 15519 15691
rect 16129 15657 16163 15691
rect 17785 15657 17819 15691
rect 7021 15589 7055 15623
rect 8585 15589 8619 15623
rect 10578 15589 10612 15623
rect 13185 15589 13219 15623
rect 1768 15521 1802 15555
rect 4721 15521 4755 15555
rect 4988 15521 5022 15555
rect 7573 15521 7607 15555
rect 15301 15521 15335 15555
rect 15761 15521 15795 15555
rect 16672 15521 16706 15555
rect 1501 15453 1535 15487
rect 7665 15453 7699 15487
rect 7849 15453 7883 15487
rect 10333 15453 10367 15487
rect 13277 15453 13311 15487
rect 13369 15453 13403 15487
rect 16405 15453 16439 15487
rect 12817 15385 12851 15419
rect 3893 15317 3927 15351
rect 6101 15317 6135 15351
rect 9413 15317 9447 15351
rect 9965 15317 9999 15351
rect 11713 15317 11747 15351
rect 1593 15113 1627 15147
rect 2421 15113 2455 15147
rect 4813 15113 4847 15147
rect 8217 15113 8251 15147
rect 8769 15113 8803 15147
rect 11161 15113 11195 15147
rect 12265 15113 12299 15147
rect 17417 15113 17451 15147
rect 19625 15113 19659 15147
rect 4261 15045 4295 15079
rect 6469 15045 6503 15079
rect 6653 15045 6687 15079
rect 6285 14977 6319 15011
rect 16957 14977 16991 15011
rect 1409 14909 1443 14943
rect 2881 14909 2915 14943
rect 3148 14909 3182 14943
rect 5365 14909 5399 14943
rect 6469 14909 6503 14943
rect 6837 14909 6871 14943
rect 7104 14909 7138 14943
rect 9781 14909 9815 14943
rect 13829 14909 13863 14943
rect 13921 14909 13955 14943
rect 19441 14909 19475 14943
rect 19901 14909 19935 14943
rect 2053 14841 2087 14875
rect 2789 14841 2823 14875
rect 9229 14841 9263 14875
rect 10048 14841 10082 14875
rect 12817 14841 12851 14875
rect 14166 14841 14200 14875
rect 15945 14841 15979 14875
rect 16773 14841 16807 14875
rect 5273 14773 5307 14807
rect 5549 14773 5583 14807
rect 9689 14773 9723 14807
rect 12909 14773 12943 14807
rect 13369 14773 13403 14807
rect 15301 14773 15335 14807
rect 16221 14773 16255 14807
rect 16405 14773 16439 14807
rect 16865 14773 16899 14807
rect 17785 14773 17819 14807
rect 1869 14569 1903 14603
rect 2421 14569 2455 14603
rect 4445 14569 4479 14603
rect 4537 14569 4571 14603
rect 7481 14569 7515 14603
rect 10057 14569 10091 14603
rect 10793 14569 10827 14603
rect 14013 14569 14047 14603
rect 15301 14569 15335 14603
rect 15669 14569 15703 14603
rect 16865 14569 16899 14603
rect 2789 14501 2823 14535
rect 3893 14501 3927 14535
rect 6368 14501 6402 14535
rect 12072 14501 12106 14535
rect 16313 14501 16347 14535
rect 2881 14433 2915 14467
rect 6108 14433 6142 14467
rect 8401 14433 8435 14467
rect 10149 14433 10183 14467
rect 11805 14433 11839 14467
rect 16773 14433 16807 14467
rect 1409 14365 1443 14399
rect 3065 14365 3099 14399
rect 4629 14365 4663 14399
rect 8585 14365 8619 14399
rect 10241 14365 10275 14399
rect 15761 14365 15795 14399
rect 15853 14365 15887 14399
rect 4077 14297 4111 14331
rect 9229 14297 9263 14331
rect 2329 14229 2363 14263
rect 3433 14229 3467 14263
rect 5089 14229 5123 14263
rect 5457 14229 5491 14263
rect 6009 14229 6043 14263
rect 8033 14229 8067 14263
rect 9689 14229 9723 14263
rect 13185 14229 13219 14263
rect 15025 14229 15059 14263
rect 1593 14025 1627 14059
rect 4353 14025 4387 14059
rect 5365 14025 5399 14059
rect 6193 14025 6227 14059
rect 6561 14025 6595 14059
rect 7389 14025 7423 14059
rect 8953 14025 8987 14059
rect 11437 14025 11471 14059
rect 12173 14025 12207 14059
rect 15209 14025 15243 14059
rect 15761 14025 15795 14059
rect 16313 14025 16347 14059
rect 17417 14025 17451 14059
rect 4169 13957 4203 13991
rect 7021 13957 7055 13991
rect 11161 13957 11195 13991
rect 2697 13889 2731 13923
rect 3249 13889 3283 13923
rect 3433 13889 3467 13923
rect 4997 13889 5031 13923
rect 8033 13889 8067 13923
rect 8217 13889 8251 13923
rect 9137 13889 9171 13923
rect 12449 13889 12483 13923
rect 16773 13889 16807 13923
rect 16957 13889 16991 13923
rect 1409 13821 1443 13855
rect 4813 13821 4847 13855
rect 7941 13821 7975 13855
rect 8585 13821 8619 13855
rect 13737 13821 13771 13855
rect 13829 13821 13863 13855
rect 2329 13753 2363 13787
rect 3157 13753 3191 13787
rect 9404 13753 9438 13787
rect 13369 13753 13403 13787
rect 14096 13753 14130 13787
rect 2789 13685 2823 13719
rect 4721 13685 4755 13719
rect 5733 13685 5767 13719
rect 7573 13685 7607 13719
rect 10517 13685 10551 13719
rect 11897 13685 11931 13719
rect 16129 13685 16163 13719
rect 16681 13685 16715 13719
rect 3157 13481 3191 13515
rect 3893 13481 3927 13515
rect 4445 13481 4479 13515
rect 5089 13481 5123 13515
rect 5917 13481 5951 13515
rect 6285 13481 6319 13515
rect 7665 13481 7699 13515
rect 8125 13481 8159 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 14013 13481 14047 13515
rect 15025 13481 15059 13515
rect 16957 13481 16991 13515
rect 19441 13481 19475 13515
rect 21097 13481 21131 13515
rect 2513 13413 2547 13447
rect 4537 13413 4571 13447
rect 5825 13345 5859 13379
rect 7481 13345 7515 13379
rect 10057 13345 10091 13379
rect 12245 13345 12279 13379
rect 15844 13345 15878 13379
rect 18317 13345 18351 13379
rect 20913 13345 20947 13379
rect 2605 13277 2639 13311
rect 2697 13277 2731 13311
rect 4629 13277 4663 13311
rect 6377 13277 6411 13311
rect 6561 13277 6595 13311
rect 8585 13277 8619 13311
rect 10241 13277 10275 13311
rect 11989 13277 12023 13311
rect 15577 13277 15611 13311
rect 18061 13277 18095 13311
rect 1593 13141 1627 13175
rect 1961 13141 1995 13175
rect 2145 13141 2179 13175
rect 4077 13141 4111 13175
rect 7021 13141 7055 13175
rect 7297 13141 7331 13175
rect 9505 13141 9539 13175
rect 13369 13141 13403 13175
rect 3985 12937 4019 12971
rect 4997 12937 5031 12971
rect 6561 12937 6595 12971
rect 8769 12937 8803 12971
rect 9229 12937 9263 12971
rect 10609 12937 10643 12971
rect 11529 12937 11563 12971
rect 11897 12937 11931 12971
rect 12173 12937 12207 12971
rect 12449 12937 12483 12971
rect 14013 12937 14047 12971
rect 16405 12937 16439 12971
rect 21281 12937 21315 12971
rect 22477 12937 22511 12971
rect 4629 12869 4663 12903
rect 2605 12801 2639 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 7389 12801 7423 12835
rect 9781 12801 9815 12835
rect 10241 12801 10275 12835
rect 12909 12801 12943 12835
rect 13093 12801 13127 12835
rect 13553 12801 13587 12835
rect 14657 12801 14691 12835
rect 17049 12801 17083 12835
rect 1409 12733 1443 12767
rect 2145 12733 2179 12767
rect 2861 12733 2895 12767
rect 5549 12733 5583 12767
rect 8401 12733 8435 12767
rect 9689 12733 9723 12767
rect 12817 12733 12851 12767
rect 14473 12733 14507 12767
rect 18889 12733 18923 12767
rect 20913 12733 20947 12767
rect 21097 12733 21131 12767
rect 21557 12733 21591 12767
rect 22293 12733 22327 12767
rect 22753 12733 22787 12767
rect 7297 12665 7331 12699
rect 9137 12665 9171 12699
rect 9597 12665 9631 12699
rect 10793 12665 10827 12699
rect 13921 12665 13955 12699
rect 14381 12665 14415 12699
rect 15301 12665 15335 12699
rect 16313 12665 16347 12699
rect 16773 12665 16807 12699
rect 18061 12665 18095 12699
rect 1593 12597 1627 12631
rect 2513 12597 2547 12631
rect 5181 12597 5215 12631
rect 6193 12597 6227 12631
rect 6837 12597 6871 12631
rect 7205 12597 7239 12631
rect 7849 12597 7883 12631
rect 15669 12597 15703 12631
rect 16865 12597 16899 12631
rect 17417 12597 17451 12631
rect 18521 12597 18555 12631
rect 3249 12393 3283 12427
rect 3893 12393 3927 12427
rect 4261 12393 4295 12427
rect 4629 12393 4663 12427
rect 6837 12393 6871 12427
rect 9321 12393 9355 12427
rect 9689 12393 9723 12427
rect 11253 12393 11287 12427
rect 11621 12393 11655 12427
rect 12541 12393 12575 12427
rect 12909 12393 12943 12427
rect 13369 12393 13403 12427
rect 15853 12393 15887 12427
rect 16405 12393 16439 12427
rect 21925 12393 21959 12427
rect 2881 12325 2915 12359
rect 5702 12325 5736 12359
rect 10149 12325 10183 12359
rect 16948 12325 16982 12359
rect 2145 12257 2179 12291
rect 2237 12257 2271 12291
rect 4077 12257 4111 12291
rect 5273 12257 5307 12291
rect 5457 12257 5491 12291
rect 8309 12257 8343 12291
rect 10057 12257 10091 12291
rect 11713 12257 11747 12291
rect 14013 12257 14047 12291
rect 15669 12257 15703 12291
rect 21741 12257 21775 12291
rect 2421 12189 2455 12223
rect 8401 12189 8435 12223
rect 8585 12189 8619 12223
rect 10333 12189 10367 12223
rect 11805 12189 11839 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 16681 12189 16715 12223
rect 1685 12121 1719 12155
rect 7757 12121 7791 12155
rect 18061 12121 18095 12155
rect 1777 12053 1811 12087
rect 7481 12053 7515 12087
rect 7941 12053 7975 12087
rect 13645 12053 13679 12087
rect 15485 12053 15519 12087
rect 4077 11849 4111 11883
rect 5181 11849 5215 11883
rect 6285 11849 6319 11883
rect 8309 11849 8343 11883
rect 10793 11849 10827 11883
rect 11253 11849 11287 11883
rect 12725 11849 12759 11883
rect 16037 11849 16071 11883
rect 17141 11849 17175 11883
rect 18061 11849 18095 11883
rect 7849 11781 7883 11815
rect 4721 11713 4755 11747
rect 5733 11713 5767 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 8493 11713 8527 11747
rect 15577 11713 15611 11747
rect 16497 11713 16531 11747
rect 16681 11713 16715 11747
rect 18613 11713 18647 11747
rect 1961 11645 1995 11679
rect 2053 11645 2087 11679
rect 2320 11645 2354 11679
rect 8749 11645 8783 11679
rect 13277 11645 13311 11679
rect 18521 11645 18555 11679
rect 19073 11645 19107 11679
rect 4997 11577 5031 11611
rect 5641 11577 5675 11611
rect 6561 11577 6595 11611
rect 7205 11577 7239 11611
rect 10425 11577 10459 11611
rect 12173 11577 12207 11611
rect 13544 11577 13578 11611
rect 17785 11577 17819 11611
rect 18429 11577 18463 11611
rect 3433 11509 3467 11543
rect 5549 11509 5583 11543
rect 6837 11509 6871 11543
rect 9873 11509 9907 11543
rect 11345 11509 11379 11543
rect 11805 11509 11839 11543
rect 13093 11509 13127 11543
rect 14657 11509 14691 11543
rect 15853 11509 15887 11543
rect 16405 11509 16439 11543
rect 17417 11509 17451 11543
rect 21741 11509 21775 11543
rect 1593 11305 1627 11339
rect 1961 11305 1995 11339
rect 2421 11305 2455 11339
rect 2881 11305 2915 11339
rect 3525 11305 3559 11339
rect 3801 11305 3835 11339
rect 5549 11305 5583 11339
rect 6009 11305 6043 11339
rect 8217 11305 8251 11339
rect 8585 11305 8619 11339
rect 8861 11305 8895 11339
rect 9873 11305 9907 11339
rect 13369 11305 13403 11339
rect 16681 11305 16715 11339
rect 17969 11305 18003 11339
rect 6460 11237 6494 11271
rect 9229 11237 9263 11271
rect 11152 11237 11186 11271
rect 13737 11237 13771 11271
rect 18337 11237 18371 11271
rect 1409 11169 1443 11203
rect 2789 11169 2823 11203
rect 4445 11169 4479 11203
rect 4537 11169 4571 11203
rect 6193 11169 6227 11203
rect 14473 11169 14507 11203
rect 15568 11169 15602 11203
rect 17785 11169 17819 11203
rect 3065 11101 3099 11135
rect 4629 11101 4663 11135
rect 10885 11101 10919 11135
rect 13829 11101 13863 11135
rect 13921 11101 13955 11135
rect 15301 11101 15335 11135
rect 2329 11033 2363 11067
rect 4077 11033 4111 11067
rect 5273 11033 5307 11067
rect 10425 11033 10459 11067
rect 12909 11033 12943 11067
rect 13277 11033 13311 11067
rect 7573 10965 7607 10999
rect 12265 10965 12299 10999
rect 17233 10965 17267 10999
rect 3525 10761 3559 10795
rect 6193 10761 6227 10795
rect 6653 10761 6687 10795
rect 8677 10761 8711 10795
rect 11161 10761 11195 10795
rect 13829 10761 13863 10795
rect 15209 10761 15243 10795
rect 16221 10761 16255 10795
rect 16957 10761 16991 10795
rect 18521 10761 18555 10795
rect 7113 10693 7147 10727
rect 11713 10693 11747 10727
rect 12173 10693 12207 10727
rect 15117 10693 15151 10727
rect 7297 10625 7331 10659
rect 12449 10625 12483 10659
rect 15761 10625 15795 10659
rect 1593 10557 1627 10591
rect 3985 10557 4019 10591
rect 4077 10557 4111 10591
rect 9689 10557 9723 10591
rect 9781 10557 9815 10591
rect 10037 10557 10071 10591
rect 16589 10557 16623 10591
rect 16773 10557 16807 10591
rect 17233 10557 17267 10591
rect 18337 10557 18371 10591
rect 18889 10557 18923 10591
rect 1860 10489 1894 10523
rect 4344 10489 4378 10523
rect 7564 10489 7598 10523
rect 9321 10489 9355 10523
rect 12694 10489 12728 10523
rect 14749 10489 14783 10523
rect 15577 10489 15611 10523
rect 2973 10421 3007 10455
rect 5457 10421 5491 10455
rect 15669 10421 15703 10455
rect 17785 10421 17819 10455
rect 1869 10217 1903 10251
rect 2421 10217 2455 10251
rect 3893 10217 3927 10251
rect 4629 10217 4663 10251
rect 4905 10217 4939 10251
rect 8677 10217 8711 10251
rect 9505 10217 9539 10251
rect 9689 10217 9723 10251
rect 10977 10217 11011 10251
rect 13277 10217 13311 10251
rect 13461 10217 13495 10251
rect 13921 10217 13955 10251
rect 17141 10217 17175 10251
rect 18429 10217 18463 10251
rect 2329 10149 2363 10183
rect 3525 10149 3559 10183
rect 5426 10149 5460 10183
rect 16006 10149 16040 10183
rect 2789 10081 2823 10115
rect 4077 10081 4111 10115
rect 5181 10081 5215 10115
rect 7573 10081 7607 10115
rect 8033 10081 8067 10115
rect 10057 10081 10091 10115
rect 11621 10081 11655 10115
rect 11713 10081 11747 10115
rect 13829 10081 13863 10115
rect 18245 10081 18279 10115
rect 1409 10013 1443 10047
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 7205 10013 7239 10047
rect 8125 10013 8159 10047
rect 8217 10013 8251 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 11805 10013 11839 10047
rect 12817 10013 12851 10047
rect 14105 10013 14139 10047
rect 15761 10013 15795 10047
rect 7665 9945 7699 9979
rect 11253 9945 11287 9979
rect 14473 9945 14507 9979
rect 6561 9877 6595 9911
rect 9137 9877 9171 9911
rect 12541 9877 12575 9911
rect 15577 9877 15611 9911
rect 2789 9673 2823 9707
rect 3525 9673 3559 9707
rect 5365 9673 5399 9707
rect 11253 9673 11287 9707
rect 13921 9673 13955 9707
rect 14289 9673 14323 9707
rect 16313 9673 16347 9707
rect 18245 9673 18279 9707
rect 1409 9605 1443 9639
rect 2421 9605 2455 9639
rect 3157 9605 3191 9639
rect 6285 9605 6319 9639
rect 7573 9605 7607 9639
rect 8033 9605 8067 9639
rect 9045 9605 9079 9639
rect 18521 9605 18555 9639
rect 2053 9537 2087 9571
rect 6837 9537 6871 9571
rect 8493 9537 8527 9571
rect 8677 9537 8711 9571
rect 10057 9537 10091 9571
rect 10241 9537 10275 9571
rect 13001 9537 13035 9571
rect 14381 9537 14415 9571
rect 16865 9537 16899 9571
rect 1777 9469 1811 9503
rect 2973 9469 3007 9503
rect 3893 9469 3927 9503
rect 3985 9469 4019 9503
rect 4241 9469 4275 9503
rect 18061 9469 18095 9503
rect 18889 9469 18923 9503
rect 11345 9401 11379 9435
rect 12173 9401 12207 9435
rect 12817 9401 12851 9435
rect 14626 9401 14660 9435
rect 1869 9333 1903 9367
rect 6009 9333 6043 9367
rect 7849 9333 7883 9367
rect 8401 9333 8435 9367
rect 9413 9333 9447 9367
rect 9597 9333 9631 9367
rect 9965 9333 9999 9367
rect 10609 9333 10643 9367
rect 11805 9333 11839 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 13461 9333 13495 9367
rect 15761 9333 15795 9367
rect 1593 9129 1627 9163
rect 1961 9129 1995 9163
rect 2329 9129 2363 9163
rect 2973 9129 3007 9163
rect 3893 9129 3927 9163
rect 4261 9129 4295 9163
rect 4629 9129 4663 9163
rect 5549 9129 5583 9163
rect 8033 9129 8067 9163
rect 11713 9129 11747 9163
rect 11897 9129 11931 9163
rect 13553 9129 13587 9163
rect 14105 9129 14139 9163
rect 14473 9129 14507 9163
rect 15761 9129 15795 9163
rect 16773 9129 16807 9163
rect 3341 9061 3375 9095
rect 6898 9061 6932 9095
rect 8677 9061 8711 9095
rect 9934 9061 9968 9095
rect 1409 8993 1443 9027
rect 2513 8993 2547 9027
rect 5457 8993 5491 9027
rect 6653 8993 6687 9027
rect 9689 8993 9723 9027
rect 5733 8925 5767 8959
rect 8953 8925 8987 8959
rect 2697 8857 2731 8891
rect 5089 8857 5123 8891
rect 15301 9061 15335 9095
rect 12429 8993 12463 9027
rect 16589 8993 16623 9027
rect 12173 8925 12207 8959
rect 9505 8789 9539 8823
rect 11069 8789 11103 8823
rect 11897 8789 11931 8823
rect 11989 8789 12023 8823
rect 1593 8585 1627 8619
rect 1961 8585 1995 8619
rect 5457 8585 5491 8619
rect 5917 8585 5951 8619
rect 6561 8585 6595 8619
rect 10241 8585 10275 8619
rect 10793 8585 10827 8619
rect 11897 8585 11931 8619
rect 12725 8585 12759 8619
rect 14289 8585 14323 8619
rect 16589 8585 16623 8619
rect 5181 8517 5215 8551
rect 9321 8517 9355 8551
rect 6929 8449 6963 8483
rect 10609 8449 10643 8483
rect 11253 8449 11287 8483
rect 11437 8449 11471 8483
rect 12909 8449 12943 8483
rect 1409 8381 1443 8415
rect 2605 8381 2639 8415
rect 7941 8381 7975 8415
rect 8197 8381 8231 8415
rect 11161 8381 11195 8415
rect 13165 8381 13199 8415
rect 9873 8313 9907 8347
rect 12173 8313 12207 8347
rect 7481 8245 7515 8279
rect 7757 8245 7791 8279
rect 1593 8041 1627 8075
rect 2237 8041 2271 8075
rect 8033 8041 8067 8075
rect 9873 8041 9907 8075
rect 11713 8041 11747 8075
rect 12265 8041 12299 8075
rect 13001 8041 13035 8075
rect 1869 7973 1903 8007
rect 1409 7905 1443 7939
rect 10333 7905 10367 7939
rect 10600 7905 10634 7939
rect 1685 7497 1719 7531
rect 10333 7497 10367 7531
rect 10701 7497 10735 7531
rect 9689 7361 9723 7395
rect 10609 5321 10643 5355
rect 9229 5117 9263 5151
rect 9137 5049 9171 5083
rect 9496 5049 9530 5083
rect 9229 4437 9263 4471
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 2130 25372 2136 25424
rect 2188 25412 2194 25424
rect 2774 25412 2780 25424
rect 2188 25384 2780 25412
rect 2188 25372 2194 25384
rect 2774 25372 2780 25384
rect 2832 25372 2838 25424
rect 3418 25372 3424 25424
rect 3476 25412 3482 25424
rect 7929 25415 7987 25421
rect 7929 25412 7941 25415
rect 3476 25384 7941 25412
rect 3476 25372 3482 25384
rect 7929 25381 7941 25384
rect 7975 25381 7987 25415
rect 7929 25375 7987 25381
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 1762 25344 1768 25356
rect 1443 25316 1768 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 1762 25304 1768 25316
rect 1820 25304 1826 25356
rect 2314 25304 2320 25356
rect 2372 25344 2378 25356
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 2372 25316 2513 25344
rect 2372 25304 2378 25316
rect 2501 25313 2513 25316
rect 2547 25313 2559 25347
rect 3050 25344 3056 25356
rect 3011 25316 3056 25344
rect 2501 25307 2559 25313
rect 3050 25304 3056 25316
rect 3108 25304 3114 25356
rect 4617 25347 4675 25353
rect 4617 25313 4629 25347
rect 4663 25344 4675 25347
rect 4663 25316 5120 25344
rect 4663 25313 4675 25316
rect 4617 25307 4675 25313
rect 5092 25288 5120 25316
rect 4706 25276 4712 25288
rect 4667 25248 4712 25276
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 4801 25279 4859 25285
rect 4801 25245 4813 25279
rect 4847 25245 4859 25279
rect 4801 25239 4859 25245
rect 1394 25168 1400 25220
rect 1452 25208 1458 25220
rect 2041 25211 2099 25217
rect 2041 25208 2053 25211
rect 1452 25180 2053 25208
rect 1452 25168 1458 25180
rect 2041 25177 2053 25180
rect 2087 25208 2099 25211
rect 2590 25208 2596 25220
rect 2087 25180 2596 25208
rect 2087 25177 2099 25180
rect 2041 25171 2099 25177
rect 2590 25168 2596 25180
rect 2648 25168 2654 25220
rect 4614 25168 4620 25220
rect 4672 25208 4678 25220
rect 4816 25208 4844 25239
rect 5074 25236 5080 25288
rect 5132 25276 5138 25288
rect 5813 25279 5871 25285
rect 5813 25276 5825 25279
rect 5132 25248 5825 25276
rect 5132 25236 5138 25248
rect 5813 25245 5825 25248
rect 5859 25245 5871 25279
rect 6914 25276 6920 25288
rect 6875 25248 6920 25276
rect 5813 25239 5871 25245
rect 6914 25236 6920 25248
rect 6972 25236 6978 25288
rect 4672 25180 4844 25208
rect 4672 25168 4678 25180
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 2406 25140 2412 25152
rect 2367 25112 2412 25140
rect 2406 25100 2412 25112
rect 2464 25100 2470 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2774 25140 2780 25152
rect 2731 25112 2780 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2774 25100 2780 25112
rect 2832 25100 2838 25152
rect 4249 25143 4307 25149
rect 4249 25109 4261 25143
rect 4295 25140 4307 25143
rect 6086 25140 6092 25152
rect 4295 25112 6092 25140
rect 4295 25109 4307 25112
rect 4249 25103 4307 25109
rect 6086 25100 6092 25112
rect 6144 25100 6150 25152
rect 7834 25140 7840 25152
rect 7795 25112 7840 25140
rect 7834 25100 7840 25112
rect 7892 25100 7898 25152
rect 12897 25143 12955 25149
rect 12897 25109 12909 25143
rect 12943 25140 12955 25143
rect 13078 25140 13084 25152
rect 12943 25112 13084 25140
rect 12943 25109 12955 25112
rect 12897 25103 12955 25109
rect 13078 25100 13084 25112
rect 13136 25100 13142 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1762 24896 1768 24948
rect 1820 24936 1826 24948
rect 1857 24939 1915 24945
rect 1857 24936 1869 24939
rect 1820 24908 1869 24936
rect 1820 24896 1826 24908
rect 1857 24905 1869 24908
rect 1903 24936 1915 24939
rect 5074 24936 5080 24948
rect 1903 24908 2452 24936
rect 1903 24905 1915 24908
rect 1857 24899 1915 24905
rect 2314 24868 2320 24880
rect 2275 24840 2320 24868
rect 2314 24828 2320 24840
rect 2372 24828 2378 24880
rect 2424 24868 2452 24908
rect 2976 24908 4752 24936
rect 5035 24908 5080 24936
rect 2976 24868 3004 24908
rect 4724 24868 4752 24908
rect 5074 24896 5080 24908
rect 5132 24896 5138 24948
rect 5350 24896 5356 24948
rect 5408 24896 5414 24948
rect 5368 24868 5396 24896
rect 2424 24840 3004 24868
rect 3068 24840 4660 24868
rect 4724 24840 5396 24868
rect 2406 24760 2412 24812
rect 2464 24800 2470 24812
rect 3068 24809 3096 24840
rect 4632 24809 4660 24840
rect 3053 24803 3111 24809
rect 3053 24800 3065 24803
rect 2464 24772 3065 24800
rect 2464 24760 2470 24772
rect 3053 24769 3065 24772
rect 3099 24769 3111 24803
rect 3053 24763 3111 24769
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24800 4675 24803
rect 5353 24803 5411 24809
rect 5353 24800 5365 24803
rect 4663 24772 5365 24800
rect 4663 24769 4675 24772
rect 4617 24763 4675 24769
rect 5353 24769 5365 24772
rect 5399 24769 5411 24803
rect 6178 24800 6184 24812
rect 5353 24763 5411 24769
rect 5552 24772 6184 24800
rect 1394 24732 1400 24744
rect 1355 24704 1400 24732
rect 1394 24692 1400 24704
rect 1452 24692 1458 24744
rect 2498 24692 2504 24744
rect 2556 24692 2562 24744
rect 2777 24735 2835 24741
rect 2777 24701 2789 24735
rect 2823 24732 2835 24735
rect 2866 24732 2872 24744
rect 2823 24704 2872 24732
rect 2823 24701 2835 24704
rect 2777 24695 2835 24701
rect 2866 24692 2872 24704
rect 2924 24692 2930 24744
rect 3510 24732 3516 24744
rect 3423 24704 3516 24732
rect 3510 24692 3516 24704
rect 3568 24732 3574 24744
rect 4341 24735 4399 24741
rect 4341 24732 4353 24735
rect 3568 24704 4353 24732
rect 3568 24692 3574 24704
rect 4341 24701 4353 24704
rect 4387 24732 4399 24735
rect 4982 24732 4988 24744
rect 4387 24704 4988 24732
rect 4387 24701 4399 24704
rect 4341 24695 4399 24701
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 5552 24741 5580 24772
rect 6178 24760 6184 24772
rect 6236 24760 6242 24812
rect 7374 24760 7380 24812
rect 7432 24800 7438 24812
rect 8297 24803 8355 24809
rect 8297 24800 8309 24803
rect 7432 24772 8309 24800
rect 7432 24760 7438 24772
rect 8297 24769 8309 24772
rect 8343 24769 8355 24803
rect 12250 24800 12256 24812
rect 12211 24772 12256 24800
rect 8297 24763 8355 24769
rect 12250 24760 12256 24772
rect 12308 24800 12314 24812
rect 12897 24803 12955 24809
rect 12897 24800 12909 24803
rect 12308 24772 12909 24800
rect 12308 24760 12314 24772
rect 12897 24769 12909 24772
rect 12943 24769 12955 24803
rect 13078 24800 13084 24812
rect 13039 24772 13084 24800
rect 12897 24763 12955 24769
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 5537 24735 5595 24741
rect 5537 24701 5549 24735
rect 5583 24701 5595 24735
rect 5537 24695 5595 24701
rect 9585 24735 9643 24741
rect 9585 24701 9597 24735
rect 9631 24732 9643 24735
rect 9677 24735 9735 24741
rect 9677 24732 9689 24735
rect 9631 24704 9689 24732
rect 9631 24701 9643 24704
rect 9585 24695 9643 24701
rect 9677 24701 9689 24704
rect 9723 24732 9735 24735
rect 9766 24732 9772 24744
rect 9723 24704 9772 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 9766 24692 9772 24704
rect 9824 24692 9830 24744
rect 1762 24624 1768 24676
rect 1820 24664 1826 24676
rect 2516 24664 2544 24692
rect 1820 24636 2544 24664
rect 3881 24667 3939 24673
rect 1820 24624 1826 24636
rect 3881 24633 3893 24667
rect 3927 24664 3939 24667
rect 7653 24667 7711 24673
rect 3927 24636 4476 24664
rect 3927 24633 3939 24636
rect 3881 24627 3939 24633
rect 4448 24608 4476 24636
rect 7653 24633 7665 24667
rect 7699 24664 7711 24667
rect 8202 24664 8208 24676
rect 7699 24636 8208 24664
rect 7699 24633 7711 24636
rect 7653 24627 7711 24633
rect 8202 24624 8208 24636
rect 8260 24624 8266 24676
rect 9217 24667 9275 24673
rect 9217 24633 9229 24667
rect 9263 24664 9275 24667
rect 9922 24667 9980 24673
rect 9922 24664 9934 24667
rect 9263 24636 9934 24664
rect 9263 24633 9275 24636
rect 9217 24627 9275 24633
rect 9922 24633 9934 24636
rect 9968 24664 9980 24667
rect 10042 24664 10048 24676
rect 9968 24636 10048 24664
rect 9968 24633 9980 24636
rect 9922 24627 9980 24633
rect 10042 24624 10048 24636
rect 10100 24624 10106 24676
rect 12805 24667 12863 24673
rect 12805 24664 12817 24667
rect 11808 24636 12817 24664
rect 11808 24608 11836 24636
rect 12805 24633 12817 24636
rect 12851 24633 12863 24667
rect 12805 24627 12863 24633
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 2314 24596 2320 24608
rect 1627 24568 2320 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 2314 24556 2320 24568
rect 2372 24556 2378 24608
rect 2409 24599 2467 24605
rect 2409 24565 2421 24599
rect 2455 24596 2467 24599
rect 2498 24596 2504 24608
rect 2455 24568 2504 24596
rect 2455 24565 2467 24568
rect 2409 24559 2467 24565
rect 2498 24556 2504 24568
rect 2556 24556 2562 24608
rect 2869 24599 2927 24605
rect 2869 24565 2881 24599
rect 2915 24596 2927 24599
rect 3050 24596 3056 24608
rect 2915 24568 3056 24596
rect 2915 24565 2927 24568
rect 2869 24559 2927 24565
rect 3050 24556 3056 24568
rect 3108 24556 3114 24608
rect 3970 24596 3976 24608
rect 3931 24568 3976 24596
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 4430 24596 4436 24608
rect 4391 24568 4436 24596
rect 4430 24556 4436 24568
rect 4488 24556 4494 24608
rect 5534 24556 5540 24608
rect 5592 24596 5598 24608
rect 5721 24599 5779 24605
rect 5721 24596 5733 24599
rect 5592 24568 5733 24596
rect 5592 24556 5598 24568
rect 5721 24565 5733 24568
rect 5767 24565 5779 24599
rect 5721 24559 5779 24565
rect 7285 24599 7343 24605
rect 7285 24565 7297 24599
rect 7331 24596 7343 24599
rect 7374 24596 7380 24608
rect 7331 24568 7380 24596
rect 7331 24565 7343 24568
rect 7285 24559 7343 24565
rect 7374 24556 7380 24568
rect 7432 24556 7438 24608
rect 7742 24596 7748 24608
rect 7703 24568 7748 24596
rect 7742 24556 7748 24568
rect 7800 24556 7806 24608
rect 7834 24556 7840 24608
rect 7892 24596 7898 24608
rect 8113 24599 8171 24605
rect 8113 24596 8125 24599
rect 7892 24568 8125 24596
rect 7892 24556 7898 24568
rect 8113 24565 8125 24568
rect 8159 24565 8171 24599
rect 8113 24559 8171 24565
rect 11057 24599 11115 24605
rect 11057 24565 11069 24599
rect 11103 24596 11115 24599
rect 11146 24596 11152 24608
rect 11103 24568 11152 24596
rect 11103 24565 11115 24568
rect 11057 24559 11115 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 11790 24596 11796 24608
rect 11751 24568 11796 24596
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 12618 24596 12624 24608
rect 12483 24568 12624 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 12618 24556 12624 24568
rect 12676 24556 12682 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1673 24395 1731 24401
rect 1673 24361 1685 24395
rect 1719 24392 1731 24395
rect 2498 24392 2504 24404
rect 1719 24364 2504 24392
rect 1719 24361 1731 24364
rect 1673 24355 1731 24361
rect 2498 24352 2504 24364
rect 2556 24352 2562 24404
rect 3970 24392 3976 24404
rect 2608 24364 3976 24392
rect 2608 24197 2636 24364
rect 3970 24352 3976 24364
rect 4028 24352 4034 24404
rect 7009 24395 7067 24401
rect 7009 24361 7021 24395
rect 7055 24392 7067 24395
rect 7742 24392 7748 24404
rect 7055 24364 7748 24392
rect 7055 24361 7067 24364
rect 7009 24355 7067 24361
rect 7742 24352 7748 24364
rect 7800 24352 7806 24404
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9732 24364 10149 24392
rect 9732 24352 9738 24364
rect 10137 24361 10149 24364
rect 10183 24392 10195 24395
rect 11054 24392 11060 24404
rect 10183 24364 11060 24392
rect 10183 24361 10195 24364
rect 10137 24355 10195 24361
rect 11054 24352 11060 24364
rect 11112 24352 11118 24404
rect 15654 24392 15660 24404
rect 15615 24364 15660 24392
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 17310 24392 17316 24404
rect 17271 24364 17316 24392
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 21818 24392 21824 24404
rect 21779 24364 21824 24392
rect 21818 24352 21824 24364
rect 21876 24352 21882 24404
rect 22922 24392 22928 24404
rect 22883 24364 22928 24392
rect 22922 24352 22928 24364
rect 22980 24352 22986 24404
rect 24026 24392 24032 24404
rect 23987 24364 24032 24392
rect 24026 24352 24032 24364
rect 24084 24352 24090 24404
rect 2866 24284 2872 24336
rect 2924 24324 2930 24336
rect 3145 24327 3203 24333
rect 3145 24324 3157 24327
rect 2924 24296 3157 24324
rect 2924 24284 2930 24296
rect 3145 24293 3157 24296
rect 3191 24324 3203 24327
rect 3786 24324 3792 24336
rect 3191 24296 3792 24324
rect 3191 24293 3203 24296
rect 3145 24287 3203 24293
rect 3786 24284 3792 24296
rect 3844 24284 3850 24336
rect 3881 24327 3939 24333
rect 3881 24293 3893 24327
rect 3927 24324 3939 24327
rect 4706 24324 4712 24336
rect 3927 24296 4712 24324
rect 3927 24293 3939 24296
rect 3881 24287 3939 24293
rect 4706 24284 4712 24296
rect 4764 24284 4770 24336
rect 7929 24327 7987 24333
rect 7929 24324 7941 24327
rect 4816 24296 7941 24324
rect 3050 24216 3056 24268
rect 3108 24256 3114 24268
rect 4816 24256 4844 24296
rect 7929 24293 7941 24296
rect 7975 24324 7987 24327
rect 8110 24324 8116 24336
rect 7975 24296 8116 24324
rect 7975 24293 7987 24296
rect 7929 24287 7987 24293
rect 8110 24284 8116 24296
rect 8168 24284 8174 24336
rect 9766 24284 9772 24336
rect 9824 24324 9830 24336
rect 9824 24296 11376 24324
rect 9824 24284 9830 24296
rect 11348 24268 11376 24296
rect 4982 24265 4988 24268
rect 4976 24256 4988 24265
rect 3108 24228 4844 24256
rect 4943 24228 4988 24256
rect 3108 24216 3114 24228
rect 4976 24219 4988 24228
rect 4982 24216 4988 24219
rect 5040 24216 5046 24268
rect 6546 24216 6552 24268
rect 6604 24256 6610 24268
rect 7837 24259 7895 24265
rect 7837 24256 7849 24259
rect 6604 24228 7849 24256
rect 6604 24216 6610 24228
rect 7837 24225 7849 24228
rect 7883 24256 7895 24259
rect 9214 24256 9220 24268
rect 7883 24228 9220 24256
rect 7883 24225 7895 24228
rect 7837 24219 7895 24225
rect 9214 24216 9220 24228
rect 9272 24256 9278 24268
rect 10045 24259 10103 24265
rect 10045 24256 10057 24259
rect 9272 24228 10057 24256
rect 9272 24216 9278 24228
rect 10045 24225 10057 24228
rect 10091 24225 10103 24259
rect 11330 24256 11336 24268
rect 11243 24228 11336 24256
rect 10045 24219 10103 24225
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 11606 24265 11612 24268
rect 11600 24256 11612 24265
rect 11567 24228 11612 24256
rect 11600 24219 11612 24228
rect 11606 24216 11612 24219
rect 11664 24216 11670 24268
rect 15470 24256 15476 24268
rect 15431 24228 15476 24256
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 17129 24259 17187 24265
rect 17129 24225 17141 24259
rect 17175 24256 17187 24259
rect 17310 24256 17316 24268
rect 17175 24228 17316 24256
rect 17175 24225 17187 24228
rect 17129 24219 17187 24225
rect 17310 24216 17316 24228
rect 17368 24216 17374 24268
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 21637 24259 21695 24265
rect 21637 24256 21649 24259
rect 21600 24228 21649 24256
rect 21600 24216 21606 24228
rect 21637 24225 21649 24228
rect 21683 24225 21695 24259
rect 22738 24256 22744 24268
rect 22699 24228 22744 24256
rect 21637 24219 21695 24225
rect 22738 24216 22744 24228
rect 22796 24216 22802 24268
rect 23842 24256 23848 24268
rect 23803 24228 23848 24256
rect 23842 24216 23848 24228
rect 23900 24216 23906 24268
rect 2041 24191 2099 24197
rect 2041 24157 2053 24191
rect 2087 24188 2099 24191
rect 2593 24191 2651 24197
rect 2593 24188 2605 24191
rect 2087 24160 2605 24188
rect 2087 24157 2099 24160
rect 2041 24151 2099 24157
rect 2593 24157 2605 24160
rect 2639 24157 2651 24191
rect 2593 24151 2651 24157
rect 2777 24191 2835 24197
rect 2777 24157 2789 24191
rect 2823 24188 2835 24191
rect 2866 24188 2872 24200
rect 2823 24160 2872 24188
rect 2823 24157 2835 24160
rect 2777 24151 2835 24157
rect 2866 24148 2872 24160
rect 2924 24148 2930 24200
rect 4430 24148 4436 24200
rect 4488 24188 4494 24200
rect 4709 24191 4767 24197
rect 4709 24188 4721 24191
rect 4488 24160 4721 24188
rect 4488 24148 4494 24160
rect 4709 24157 4721 24160
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 8021 24191 8079 24197
rect 8021 24157 8033 24191
rect 8067 24157 8079 24191
rect 8021 24151 8079 24157
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24188 9551 24191
rect 9950 24188 9956 24200
rect 9539 24160 9956 24188
rect 9539 24157 9551 24160
rect 9493 24151 9551 24157
rect 7374 24120 7380 24132
rect 7335 24092 7380 24120
rect 7374 24080 7380 24092
rect 7432 24120 7438 24132
rect 8036 24120 8064 24151
rect 9950 24148 9956 24160
rect 10008 24188 10014 24200
rect 10321 24191 10379 24197
rect 10321 24188 10333 24191
rect 10008 24160 10333 24188
rect 10008 24148 10014 24160
rect 10321 24157 10333 24160
rect 10367 24188 10379 24191
rect 10367 24160 10456 24188
rect 10367 24157 10379 24160
rect 10321 24151 10379 24157
rect 7432 24092 8064 24120
rect 7432 24080 7438 24092
rect 2133 24055 2191 24061
rect 2133 24021 2145 24055
rect 2179 24052 2191 24055
rect 2222 24052 2228 24064
rect 2179 24024 2228 24052
rect 2179 24021 2191 24024
rect 2133 24015 2191 24021
rect 2222 24012 2228 24024
rect 2280 24012 2286 24064
rect 4341 24055 4399 24061
rect 4341 24021 4353 24055
rect 4387 24052 4399 24055
rect 4614 24052 4620 24064
rect 4387 24024 4620 24052
rect 4387 24021 4399 24024
rect 4341 24015 4399 24021
rect 4614 24012 4620 24024
rect 4672 24052 4678 24064
rect 6089 24055 6147 24061
rect 6089 24052 6101 24055
rect 4672 24024 6101 24052
rect 4672 24012 4678 24024
rect 6089 24021 6101 24024
rect 6135 24021 6147 24055
rect 7466 24052 7472 24064
rect 7427 24024 7472 24052
rect 6089 24015 6147 24021
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 9677 24055 9735 24061
rect 9677 24021 9689 24055
rect 9723 24052 9735 24055
rect 10134 24052 10140 24064
rect 9723 24024 10140 24052
rect 9723 24021 9735 24024
rect 9677 24015 9735 24021
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 10428 24052 10456 24160
rect 12713 24055 12771 24061
rect 12713 24052 12725 24055
rect 10428 24024 12725 24052
rect 12713 24021 12725 24024
rect 12759 24021 12771 24055
rect 12713 24015 12771 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1673 23851 1731 23857
rect 1673 23817 1685 23851
rect 1719 23848 1731 23851
rect 2406 23848 2412 23860
rect 1719 23820 2412 23848
rect 1719 23817 1731 23820
rect 1673 23811 1731 23817
rect 2406 23808 2412 23820
rect 2464 23808 2470 23860
rect 3878 23808 3884 23860
rect 3936 23848 3942 23860
rect 4341 23851 4399 23857
rect 4341 23848 4353 23851
rect 3936 23820 4353 23848
rect 3936 23808 3942 23820
rect 4341 23817 4353 23820
rect 4387 23817 4399 23851
rect 4341 23811 4399 23817
rect 2133 23647 2191 23653
rect 2133 23613 2145 23647
rect 2179 23613 2191 23647
rect 4356 23644 4384 23811
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 4893 23851 4951 23857
rect 4893 23848 4905 23851
rect 4764 23820 4905 23848
rect 4764 23808 4770 23820
rect 4893 23817 4905 23820
rect 4939 23817 4951 23851
rect 8110 23848 8116 23860
rect 8071 23820 8116 23848
rect 4893 23811 4951 23817
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 9214 23848 9220 23860
rect 9175 23820 9220 23848
rect 9214 23808 9220 23820
rect 9272 23808 9278 23860
rect 9674 23848 9680 23860
rect 9635 23820 9680 23848
rect 9674 23808 9680 23820
rect 9732 23808 9738 23860
rect 10042 23808 10048 23860
rect 10100 23848 10106 23860
rect 11149 23851 11207 23857
rect 11149 23848 11161 23851
rect 10100 23820 11161 23848
rect 10100 23808 10106 23820
rect 11149 23817 11161 23820
rect 11195 23817 11207 23851
rect 11149 23811 11207 23817
rect 11330 23808 11336 23860
rect 11388 23848 11394 23860
rect 11698 23848 11704 23860
rect 11388 23820 11704 23848
rect 11388 23808 11394 23820
rect 11698 23808 11704 23820
rect 11756 23808 11762 23860
rect 16390 23848 16396 23860
rect 16351 23820 16396 23848
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 18598 23848 18604 23860
rect 18559 23820 18604 23848
rect 18598 23808 18604 23820
rect 18656 23808 18662 23860
rect 19705 23851 19763 23857
rect 19705 23817 19717 23851
rect 19751 23848 19763 23851
rect 21358 23848 21364 23860
rect 19751 23820 21364 23848
rect 19751 23817 19763 23820
rect 19705 23811 19763 23817
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 21910 23848 21916 23860
rect 21871 23820 21916 23848
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 20809 23783 20867 23789
rect 20809 23749 20821 23783
rect 20855 23780 20867 23783
rect 21818 23780 21824 23792
rect 20855 23752 21824 23780
rect 20855 23749 20867 23752
rect 20809 23743 20867 23749
rect 21818 23740 21824 23752
rect 21876 23740 21882 23792
rect 23845 23783 23903 23789
rect 23845 23749 23857 23783
rect 23891 23780 23903 23783
rect 25314 23780 25320 23792
rect 23891 23752 25320 23780
rect 23891 23749 23903 23752
rect 23845 23743 23903 23749
rect 25314 23740 25320 23752
rect 25372 23740 25378 23792
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 5350 23712 5356 23724
rect 4847 23684 5356 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 5350 23672 5356 23684
rect 5408 23672 5414 23724
rect 5442 23672 5448 23724
rect 5500 23712 5506 23724
rect 5500 23684 5545 23712
rect 5500 23672 5506 23684
rect 7006 23672 7012 23724
rect 7064 23712 7070 23724
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7064 23684 7665 23712
rect 7064 23672 7070 23684
rect 7653 23681 7665 23684
rect 7699 23681 7711 23715
rect 7653 23675 7711 23681
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23712 8723 23715
rect 8711 23684 9904 23712
rect 8711 23681 8723 23684
rect 8665 23675 8723 23681
rect 5258 23644 5264 23656
rect 4356 23616 5264 23644
rect 2133 23607 2191 23613
rect 2041 23511 2099 23517
rect 2041 23477 2053 23511
rect 2087 23508 2099 23511
rect 2148 23508 2176 23607
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 6822 23604 6828 23656
rect 6880 23644 6886 23656
rect 7466 23644 7472 23656
rect 6880 23616 7472 23644
rect 6880 23604 6886 23616
rect 7466 23604 7472 23616
rect 7524 23604 7530 23656
rect 7561 23647 7619 23653
rect 7561 23613 7573 23647
rect 7607 23644 7619 23647
rect 7742 23644 7748 23656
rect 7607 23616 7748 23644
rect 7607 23613 7619 23616
rect 7561 23607 7619 23613
rect 7742 23604 7748 23616
rect 7800 23604 7806 23656
rect 9490 23604 9496 23656
rect 9548 23644 9554 23656
rect 9766 23644 9772 23656
rect 9548 23616 9772 23644
rect 9548 23604 9554 23616
rect 9766 23604 9772 23616
rect 9824 23604 9830 23656
rect 2406 23585 2412 23588
rect 2400 23576 2412 23585
rect 2367 23548 2412 23576
rect 2400 23539 2412 23548
rect 2464 23576 2470 23588
rect 2958 23576 2964 23588
rect 2464 23548 2964 23576
rect 2406 23536 2412 23539
rect 2464 23536 2470 23548
rect 2958 23536 2964 23548
rect 3016 23536 3022 23588
rect 6638 23576 6644 23588
rect 5920 23548 6644 23576
rect 2682 23508 2688 23520
rect 2087 23480 2688 23508
rect 2087 23477 2099 23480
rect 2041 23471 2099 23477
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 2866 23468 2872 23520
rect 2924 23508 2930 23520
rect 3513 23511 3571 23517
rect 3513 23508 3525 23511
rect 2924 23480 3525 23508
rect 2924 23468 2930 23480
rect 3513 23477 3525 23480
rect 3559 23477 3571 23511
rect 3513 23471 3571 23477
rect 4430 23468 4436 23520
rect 4488 23508 4494 23520
rect 5920 23517 5948 23548
rect 6638 23536 6644 23548
rect 6696 23536 6702 23588
rect 9876 23576 9904 23684
rect 13725 23647 13783 23653
rect 13725 23644 13737 23647
rect 13556 23616 13737 23644
rect 9950 23576 9956 23588
rect 9876 23548 9956 23576
rect 9950 23536 9956 23548
rect 10008 23585 10014 23588
rect 10008 23579 10072 23585
rect 10008 23545 10026 23579
rect 10060 23545 10072 23579
rect 10008 23539 10072 23545
rect 10008 23536 10014 23539
rect 11054 23536 11060 23588
rect 11112 23576 11118 23588
rect 11606 23576 11612 23588
rect 11112 23548 11612 23576
rect 11112 23536 11118 23548
rect 11606 23536 11612 23548
rect 11664 23576 11670 23588
rect 12069 23579 12127 23585
rect 12069 23576 12081 23579
rect 11664 23548 12081 23576
rect 11664 23536 11670 23548
rect 12069 23545 12081 23548
rect 12115 23576 12127 23579
rect 12342 23576 12348 23588
rect 12115 23548 12348 23576
rect 12115 23545 12127 23548
rect 12069 23539 12127 23545
rect 12342 23536 12348 23548
rect 12400 23536 12406 23588
rect 13556 23520 13584 23616
rect 13725 23613 13737 23616
rect 13771 23613 13783 23647
rect 13725 23607 13783 23613
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 18414 23644 18420 23656
rect 16255 23616 16896 23644
rect 18375 23616 18420 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 13814 23536 13820 23588
rect 13872 23576 13878 23588
rect 13970 23579 14028 23585
rect 13970 23576 13982 23579
rect 13872 23548 13982 23576
rect 13872 23536 13878 23548
rect 13970 23545 13982 23548
rect 14016 23545 14028 23579
rect 13970 23539 14028 23545
rect 5905 23511 5963 23517
rect 5905 23508 5917 23511
rect 4488 23480 5917 23508
rect 4488 23468 4494 23480
rect 5905 23477 5917 23480
rect 5951 23477 5963 23511
rect 6546 23508 6552 23520
rect 6507 23480 6552 23508
rect 5905 23471 5963 23477
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 6730 23468 6736 23520
rect 6788 23508 6794 23520
rect 7101 23511 7159 23517
rect 7101 23508 7113 23511
rect 6788 23480 7113 23508
rect 6788 23468 6794 23480
rect 7101 23477 7113 23480
rect 7147 23477 7159 23511
rect 7101 23471 7159 23477
rect 8757 23511 8815 23517
rect 8757 23477 8769 23511
rect 8803 23508 8815 23511
rect 9674 23508 9680 23520
rect 8803 23480 9680 23508
rect 8803 23477 8815 23480
rect 8757 23471 8815 23477
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 12710 23508 12716 23520
rect 12671 23480 12716 23508
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 13538 23508 13544 23520
rect 13499 23480 13544 23508
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 15102 23508 15108 23520
rect 15063 23480 15108 23508
rect 15102 23468 15108 23480
rect 15160 23468 15166 23520
rect 15470 23468 15476 23520
rect 15528 23508 15534 23520
rect 16868 23517 16896 23616
rect 18414 23604 18420 23616
rect 18472 23644 18478 23656
rect 18969 23647 19027 23653
rect 18969 23644 18981 23647
rect 18472 23616 18981 23644
rect 18472 23604 18478 23616
rect 18969 23613 18981 23616
rect 19015 23613 19027 23647
rect 18969 23607 19027 23613
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 19521 23647 19579 23653
rect 19521 23644 19533 23647
rect 19392 23616 19533 23644
rect 19392 23604 19398 23616
rect 19521 23613 19533 23616
rect 19567 23644 19579 23647
rect 20073 23647 20131 23653
rect 20073 23644 20085 23647
rect 19567 23616 20085 23644
rect 19567 23613 19579 23616
rect 19521 23607 19579 23613
rect 20073 23613 20085 23616
rect 20119 23613 20131 23647
rect 20073 23607 20131 23613
rect 20625 23647 20683 23653
rect 20625 23613 20637 23647
rect 20671 23613 20683 23647
rect 20625 23607 20683 23613
rect 19242 23536 19248 23588
rect 19300 23576 19306 23588
rect 20640 23576 20668 23607
rect 21174 23604 21180 23656
rect 21232 23644 21238 23656
rect 21729 23647 21787 23653
rect 21729 23644 21741 23647
rect 21232 23616 21741 23644
rect 21232 23604 21238 23616
rect 21729 23613 21741 23616
rect 21775 23644 21787 23647
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 21775 23616 22293 23644
rect 21775 23613 21787 23616
rect 21729 23607 21787 23613
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 22281 23607 22339 23613
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 23532 23616 23673 23644
rect 23532 23604 23538 23616
rect 23661 23613 23673 23616
rect 23707 23613 23719 23647
rect 23661 23607 23719 23613
rect 21269 23579 21327 23585
rect 21269 23576 21281 23579
rect 19300 23548 21281 23576
rect 19300 23536 19306 23548
rect 21269 23545 21281 23548
rect 21315 23545 21327 23579
rect 23676 23576 23704 23607
rect 23842 23604 23848 23656
rect 23900 23644 23906 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 23900 23616 24593 23644
rect 23900 23604 23906 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24762 23644 24768 23656
rect 24723 23616 24768 23644
rect 24581 23607 24639 23613
rect 24762 23604 24768 23616
rect 24820 23644 24826 23656
rect 25317 23647 25375 23653
rect 25317 23644 25329 23647
rect 24820 23616 25329 23644
rect 24820 23604 24826 23616
rect 25317 23613 25329 23616
rect 25363 23613 25375 23647
rect 25317 23607 25375 23613
rect 24213 23579 24271 23585
rect 24213 23576 24225 23579
rect 23676 23548 24225 23576
rect 21269 23539 21327 23545
rect 24213 23545 24225 23548
rect 24259 23545 24271 23579
rect 24213 23539 24271 23545
rect 15657 23511 15715 23517
rect 15657 23508 15669 23511
rect 15528 23480 15669 23508
rect 15528 23468 15534 23480
rect 15657 23477 15669 23480
rect 15703 23477 15715 23511
rect 15657 23471 15715 23477
rect 16853 23511 16911 23517
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 16942 23508 16948 23520
rect 16899 23480 16948 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 17221 23511 17279 23517
rect 17221 23477 17233 23511
rect 17267 23508 17279 23511
rect 17310 23508 17316 23520
rect 17267 23480 17316 23508
rect 17267 23477 17279 23480
rect 17221 23471 17279 23477
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 21542 23508 21548 23520
rect 21503 23480 21548 23508
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 22738 23508 22744 23520
rect 22699 23480 22744 23508
rect 22738 23468 22744 23480
rect 22796 23468 22802 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2317 23307 2375 23313
rect 2317 23273 2329 23307
rect 2363 23304 2375 23307
rect 2363 23276 2820 23304
rect 2363 23273 2375 23276
rect 2317 23267 2375 23273
rect 2130 23196 2136 23248
rect 2188 23236 2194 23248
rect 2409 23239 2467 23245
rect 2409 23236 2421 23239
rect 2188 23208 2421 23236
rect 2188 23196 2194 23208
rect 2409 23205 2421 23208
rect 2455 23236 2467 23239
rect 2498 23236 2504 23248
rect 2455 23208 2504 23236
rect 2455 23205 2467 23208
rect 2409 23199 2467 23205
rect 2498 23196 2504 23208
rect 2556 23196 2562 23248
rect 2792 23168 2820 23276
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 2961 23307 3019 23313
rect 2961 23304 2973 23307
rect 2924 23276 2973 23304
rect 2924 23264 2930 23276
rect 2961 23273 2973 23276
rect 3007 23273 3019 23307
rect 2961 23267 3019 23273
rect 3881 23307 3939 23313
rect 3881 23273 3893 23307
rect 3927 23304 3939 23307
rect 4525 23307 4583 23313
rect 4525 23304 4537 23307
rect 3927 23276 4537 23304
rect 3927 23273 3939 23276
rect 3881 23267 3939 23273
rect 4525 23273 4537 23276
rect 4571 23304 4583 23307
rect 4982 23304 4988 23316
rect 4571 23276 4988 23304
rect 4571 23273 4583 23276
rect 4525 23267 4583 23273
rect 4982 23264 4988 23276
rect 5040 23264 5046 23316
rect 6641 23307 6699 23313
rect 6641 23273 6653 23307
rect 6687 23304 6699 23307
rect 6822 23304 6828 23316
rect 6687 23276 6828 23304
rect 6687 23273 6699 23276
rect 6641 23267 6699 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 7006 23304 7012 23316
rect 6967 23276 7012 23304
rect 7006 23264 7012 23276
rect 7064 23304 7070 23316
rect 8481 23307 8539 23313
rect 8481 23304 8493 23307
rect 7064 23276 8493 23304
rect 7064 23264 7070 23276
rect 8481 23273 8493 23276
rect 8527 23273 8539 23307
rect 9490 23304 9496 23316
rect 9451 23276 9496 23304
rect 8481 23267 8539 23273
rect 9490 23264 9496 23276
rect 9548 23264 9554 23316
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 13173 23307 13231 23313
rect 13173 23304 13185 23307
rect 12492 23276 13185 23304
rect 12492 23264 12498 23276
rect 13173 23273 13185 23276
rect 13219 23273 13231 23307
rect 13173 23267 13231 23273
rect 15473 23307 15531 23313
rect 15473 23273 15485 23307
rect 15519 23304 15531 23307
rect 16482 23304 16488 23316
rect 15519 23276 16488 23304
rect 15519 23273 15531 23276
rect 15473 23267 15531 23273
rect 16482 23264 16488 23276
rect 16540 23264 16546 23316
rect 16758 23304 16764 23316
rect 16719 23276 16764 23304
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 18049 23307 18107 23313
rect 18049 23273 18061 23307
rect 18095 23304 18107 23307
rect 19334 23304 19340 23316
rect 18095 23276 19340 23304
rect 18095 23273 18107 23276
rect 18049 23267 18107 23273
rect 19334 23264 19340 23276
rect 19392 23264 19398 23316
rect 21085 23307 21143 23313
rect 21085 23273 21097 23307
rect 21131 23304 21143 23307
rect 21542 23304 21548 23316
rect 21131 23276 21548 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 21542 23264 21548 23276
rect 21600 23264 21606 23316
rect 22370 23304 22376 23316
rect 22331 23276 22376 23304
rect 22370 23264 22376 23276
rect 22428 23264 22434 23316
rect 23477 23307 23535 23313
rect 23477 23273 23489 23307
rect 23523 23304 23535 23307
rect 23842 23304 23848 23316
rect 23523 23276 23848 23304
rect 23523 23273 23535 23276
rect 23477 23267 23535 23273
rect 23842 23264 23848 23276
rect 23900 23264 23906 23316
rect 9766 23196 9772 23248
rect 9824 23236 9830 23248
rect 10134 23236 10140 23248
rect 9824 23208 10140 23236
rect 9824 23196 9830 23208
rect 10134 23196 10140 23208
rect 10192 23196 10198 23248
rect 12066 23245 12072 23248
rect 12060 23236 12072 23245
rect 12027 23208 12072 23236
rect 12060 23199 12072 23208
rect 12066 23196 12072 23199
rect 12124 23196 12130 23248
rect 3050 23168 3056 23180
rect 2792 23140 3056 23168
rect 3050 23128 3056 23140
rect 3108 23168 3114 23180
rect 3418 23168 3424 23180
rect 3108 23140 3424 23168
rect 3108 23128 3114 23140
rect 3418 23128 3424 23140
rect 3476 23128 3482 23180
rect 4430 23128 4436 23180
rect 4488 23168 4494 23180
rect 4617 23171 4675 23177
rect 4617 23168 4629 23171
rect 4488 23140 4629 23168
rect 4488 23128 4494 23140
rect 4617 23137 4629 23140
rect 4663 23137 4675 23171
rect 4617 23131 4675 23137
rect 4706 23128 4712 23180
rect 4764 23168 4770 23180
rect 4873 23171 4931 23177
rect 4873 23168 4885 23171
rect 4764 23140 4885 23168
rect 4764 23128 4770 23140
rect 4873 23137 4885 23140
rect 4919 23137 4931 23171
rect 4873 23131 4931 23137
rect 6638 23128 6644 23180
rect 6696 23168 6702 23180
rect 7098 23168 7104 23180
rect 6696 23140 7104 23168
rect 6696 23128 6702 23140
rect 7098 23128 7104 23140
rect 7156 23128 7162 23180
rect 7374 23177 7380 23180
rect 7368 23168 7380 23177
rect 7335 23140 7380 23168
rect 7368 23131 7380 23140
rect 7374 23128 7380 23131
rect 7432 23128 7438 23180
rect 9674 23128 9680 23180
rect 9732 23168 9738 23180
rect 10045 23171 10103 23177
rect 10045 23168 10057 23171
rect 9732 23140 10057 23168
rect 9732 23128 9738 23140
rect 10045 23137 10057 23140
rect 10091 23137 10103 23171
rect 10045 23131 10103 23137
rect 11698 23128 11704 23180
rect 11756 23168 11762 23180
rect 11793 23171 11851 23177
rect 11793 23168 11805 23171
rect 11756 23140 11805 23168
rect 11756 23128 11762 23140
rect 11793 23137 11805 23140
rect 11839 23137 11851 23171
rect 11793 23131 11851 23137
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 15562 23168 15568 23180
rect 15335 23140 15568 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 15562 23128 15568 23140
rect 15620 23128 15626 23180
rect 16574 23168 16580 23180
rect 16535 23140 16580 23168
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 17862 23168 17868 23180
rect 17823 23140 17868 23168
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 18874 23168 18880 23180
rect 18835 23140 18880 23168
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 20714 23128 20720 23180
rect 20772 23168 20778 23180
rect 20901 23171 20959 23177
rect 20901 23168 20913 23171
rect 20772 23140 20913 23168
rect 20772 23128 20778 23140
rect 20901 23137 20913 23140
rect 20947 23137 20959 23171
rect 22186 23168 22192 23180
rect 22147 23140 22192 23168
rect 20901 23131 20959 23137
rect 22186 23128 22192 23140
rect 22244 23128 22250 23180
rect 23290 23168 23296 23180
rect 23251 23140 23296 23168
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23069 2559 23103
rect 2501 23063 2559 23069
rect 2516 23032 2544 23063
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 10229 23103 10287 23109
rect 10229 23100 10241 23103
rect 10192 23072 10241 23100
rect 10192 23060 10198 23072
rect 10229 23069 10241 23072
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 2866 23032 2872 23044
rect 1780 23004 2872 23032
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 1780 22973 1808 23004
rect 2866 22992 2872 23004
rect 2924 22992 2930 23044
rect 19061 23035 19119 23041
rect 19061 23001 19073 23035
rect 19107 23032 19119 23035
rect 19242 23032 19248 23044
rect 19107 23004 19248 23032
rect 19107 23001 19119 23004
rect 19061 22995 19119 23001
rect 19242 22992 19248 23004
rect 19300 22992 19306 23044
rect 1765 22967 1823 22973
rect 1765 22964 1777 22967
rect 1728 22936 1777 22964
rect 1728 22924 1734 22936
rect 1765 22933 1777 22936
rect 1811 22933 1823 22967
rect 1765 22927 1823 22933
rect 1949 22967 2007 22973
rect 1949 22933 1961 22967
rect 1995 22964 2007 22967
rect 2130 22964 2136 22976
rect 1995 22936 2136 22964
rect 1995 22933 2007 22936
rect 1949 22927 2007 22933
rect 2130 22924 2136 22936
rect 2188 22924 2194 22976
rect 5997 22967 6055 22973
rect 5997 22933 6009 22967
rect 6043 22964 6055 22967
rect 6270 22964 6276 22976
rect 6043 22936 6276 22964
rect 6043 22933 6055 22936
rect 5997 22927 6055 22933
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 9677 22967 9735 22973
rect 9677 22933 9689 22967
rect 9723 22964 9735 22967
rect 10042 22964 10048 22976
rect 9723 22936 10048 22964
rect 9723 22933 9735 22936
rect 9677 22927 9735 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 10778 22964 10784 22976
rect 10739 22936 10784 22964
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 13814 22964 13820 22976
rect 13775 22936 13820 22964
rect 13814 22924 13820 22936
rect 13872 22924 13878 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2498 22720 2504 22772
rect 2556 22760 2562 22772
rect 4617 22763 4675 22769
rect 4617 22760 4629 22763
rect 2556 22732 4629 22760
rect 2556 22720 2562 22732
rect 4617 22729 4629 22732
rect 4663 22729 4675 22763
rect 7098 22760 7104 22772
rect 7059 22732 7104 22760
rect 4617 22723 4675 22729
rect 2225 22559 2283 22565
rect 2225 22556 2237 22559
rect 1596 22528 2237 22556
rect 1486 22380 1492 22432
rect 1544 22420 1550 22432
rect 1596 22429 1624 22528
rect 2225 22525 2237 22528
rect 2271 22556 2283 22559
rect 4249 22559 4307 22565
rect 4249 22556 4261 22559
rect 2271 22528 4261 22556
rect 2271 22525 2283 22528
rect 2225 22519 2283 22525
rect 2700 22500 2728 22528
rect 4249 22525 4261 22528
rect 4295 22525 4307 22559
rect 4632 22556 4660 22723
rect 7098 22720 7104 22732
rect 7156 22760 7162 22772
rect 7285 22763 7343 22769
rect 7285 22760 7297 22763
rect 7156 22732 7297 22760
rect 7156 22720 7162 22732
rect 7285 22729 7297 22732
rect 7331 22760 7343 22763
rect 7469 22763 7527 22769
rect 7469 22760 7481 22763
rect 7331 22732 7481 22760
rect 7331 22729 7343 22732
rect 7285 22723 7343 22729
rect 7469 22729 7481 22732
rect 7515 22760 7527 22763
rect 8018 22760 8024 22772
rect 7515 22732 8024 22760
rect 7515 22729 7527 22732
rect 7469 22723 7527 22729
rect 8018 22720 8024 22732
rect 8076 22720 8082 22772
rect 9674 22760 9680 22772
rect 9635 22732 9680 22760
rect 9674 22720 9680 22732
rect 9732 22720 9738 22772
rect 10134 22720 10140 22772
rect 10192 22760 10198 22772
rect 11425 22763 11483 22769
rect 11425 22760 11437 22763
rect 10192 22732 11437 22760
rect 10192 22720 10198 22732
rect 11425 22729 11437 22732
rect 11471 22729 11483 22763
rect 11425 22723 11483 22729
rect 11698 22720 11704 22772
rect 11756 22760 11762 22772
rect 11793 22763 11851 22769
rect 11793 22760 11805 22763
rect 11756 22732 11805 22760
rect 11756 22720 11762 22732
rect 11793 22729 11805 22732
rect 11839 22760 11851 22763
rect 11974 22760 11980 22772
rect 11839 22732 11980 22760
rect 11839 22729 11851 22732
rect 11793 22723 11851 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12066 22720 12072 22772
rect 12124 22760 12130 22772
rect 12161 22763 12219 22769
rect 12161 22760 12173 22763
rect 12124 22732 12173 22760
rect 12124 22720 12130 22732
rect 12161 22729 12173 22732
rect 12207 22729 12219 22763
rect 12161 22723 12219 22729
rect 13814 22720 13820 22772
rect 13872 22760 13878 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 13872 22732 14933 22760
rect 13872 22720 13878 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 16298 22760 16304 22772
rect 16259 22732 16304 22760
rect 14921 22723 14979 22729
rect 16298 22720 16304 22732
rect 16356 22720 16362 22772
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 16758 22760 16764 22772
rect 16632 22732 16764 22760
rect 16632 22720 16638 22732
rect 16758 22720 16764 22732
rect 16816 22760 16822 22772
rect 16945 22763 17003 22769
rect 16945 22760 16957 22763
rect 16816 22732 16957 22760
rect 16816 22720 16822 22732
rect 16945 22729 16957 22732
rect 16991 22729 17003 22763
rect 16945 22723 17003 22729
rect 10413 22695 10471 22701
rect 10413 22661 10425 22695
rect 10459 22661 10471 22695
rect 10413 22655 10471 22661
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 6270 22624 6276 22636
rect 5859 22596 6276 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 6270 22584 6276 22596
rect 6328 22584 6334 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 7374 22624 7380 22636
rect 6687 22596 7380 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 7374 22584 7380 22596
rect 7432 22624 7438 22636
rect 7432 22596 7788 22624
rect 7432 22584 7438 22596
rect 5537 22559 5595 22565
rect 5537 22556 5549 22559
rect 4632 22528 5549 22556
rect 4249 22519 4307 22525
rect 5537 22525 5549 22528
rect 5583 22556 5595 22559
rect 6546 22556 6552 22568
rect 5583 22528 6552 22556
rect 5583 22525 5595 22528
rect 5537 22519 5595 22525
rect 6546 22516 6552 22528
rect 6604 22516 6610 22568
rect 7285 22559 7343 22565
rect 7285 22525 7297 22559
rect 7331 22556 7343 22559
rect 7653 22559 7711 22565
rect 7653 22556 7665 22559
rect 7331 22528 7665 22556
rect 7331 22525 7343 22528
rect 7285 22519 7343 22525
rect 7653 22525 7665 22528
rect 7699 22525 7711 22559
rect 7760 22556 7788 22596
rect 8202 22556 8208 22568
rect 7760 22528 8208 22556
rect 7653 22519 7711 22525
rect 8202 22516 8208 22528
rect 8260 22516 8266 22568
rect 1670 22448 1676 22500
rect 1728 22488 1734 22500
rect 2470 22491 2528 22497
rect 2470 22488 2482 22491
rect 1728 22460 2482 22488
rect 1728 22448 1734 22460
rect 2470 22457 2482 22460
rect 2516 22457 2528 22491
rect 2470 22451 2528 22457
rect 2682 22448 2688 22500
rect 2740 22448 2746 22500
rect 5077 22491 5135 22497
rect 5077 22457 5089 22491
rect 5123 22488 5135 22491
rect 5629 22491 5687 22497
rect 5629 22488 5641 22491
rect 5123 22460 5641 22488
rect 5123 22457 5135 22460
rect 5077 22451 5135 22457
rect 5629 22457 5641 22460
rect 5675 22488 5687 22491
rect 5994 22488 6000 22500
rect 5675 22460 6000 22488
rect 5675 22457 5687 22460
rect 5629 22451 5687 22457
rect 5994 22448 6000 22460
rect 6052 22448 6058 22500
rect 7006 22448 7012 22500
rect 7064 22488 7070 22500
rect 7558 22488 7564 22500
rect 7064 22460 7564 22488
rect 7064 22448 7070 22460
rect 7558 22448 7564 22460
rect 7616 22488 7622 22500
rect 7898 22491 7956 22497
rect 7898 22488 7910 22491
rect 7616 22460 7910 22488
rect 7616 22448 7622 22460
rect 7898 22457 7910 22460
rect 7944 22457 7956 22491
rect 10428 22488 10456 22655
rect 10778 22584 10784 22636
rect 10836 22624 10842 22636
rect 10873 22627 10931 22633
rect 10873 22624 10885 22627
rect 10836 22596 10885 22624
rect 10836 22584 10842 22596
rect 10873 22593 10885 22596
rect 10919 22593 10931 22627
rect 10873 22587 10931 22593
rect 10965 22627 11023 22633
rect 10965 22593 10977 22627
rect 11011 22624 11023 22627
rect 11054 22624 11060 22636
rect 11011 22596 11060 22624
rect 11011 22593 11023 22596
rect 10965 22587 11023 22593
rect 10686 22516 10692 22568
rect 10744 22556 10750 22568
rect 10980 22556 11008 22587
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 13538 22556 13544 22568
rect 10744 22528 11008 22556
rect 13451 22528 13544 22556
rect 10744 22516 10750 22528
rect 13538 22516 13544 22528
rect 13596 22516 13602 22568
rect 15838 22516 15844 22568
rect 15896 22556 15902 22568
rect 16117 22559 16175 22565
rect 16117 22556 16129 22559
rect 15896 22528 16129 22556
rect 15896 22516 15902 22528
rect 16117 22525 16129 22528
rect 16163 22556 16175 22559
rect 16577 22559 16635 22565
rect 16577 22556 16589 22559
rect 16163 22528 16589 22556
rect 16163 22525 16175 22528
rect 16117 22519 16175 22525
rect 16577 22525 16589 22528
rect 16623 22525 16635 22559
rect 16577 22519 16635 22525
rect 10870 22488 10876 22500
rect 10428 22460 10876 22488
rect 7898 22451 7956 22457
rect 10870 22448 10876 22460
rect 10928 22448 10934 22500
rect 12434 22448 12440 22500
rect 12492 22488 12498 22500
rect 13357 22491 13415 22497
rect 13357 22488 13369 22491
rect 12492 22460 12537 22488
rect 12912 22460 13369 22488
rect 12492 22448 12498 22460
rect 1581 22423 1639 22429
rect 1581 22420 1593 22423
rect 1544 22392 1593 22420
rect 1544 22380 1550 22392
rect 1581 22389 1593 22392
rect 1627 22389 1639 22423
rect 1581 22383 1639 22389
rect 2041 22423 2099 22429
rect 2041 22389 2053 22423
rect 2087 22420 2099 22423
rect 2590 22420 2596 22432
rect 2087 22392 2596 22420
rect 2087 22389 2099 22392
rect 2041 22383 2099 22389
rect 2590 22380 2596 22392
rect 2648 22380 2654 22432
rect 2866 22380 2872 22432
rect 2924 22420 2930 22432
rect 3605 22423 3663 22429
rect 3605 22420 3617 22423
rect 2924 22392 3617 22420
rect 2924 22380 2930 22392
rect 3605 22389 3617 22392
rect 3651 22420 3663 22423
rect 3970 22420 3976 22432
rect 3651 22392 3976 22420
rect 3651 22389 3663 22392
rect 3605 22383 3663 22389
rect 3970 22380 3976 22392
rect 4028 22380 4034 22432
rect 5166 22420 5172 22432
rect 5127 22392 5172 22420
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 6270 22420 6276 22432
rect 6231 22392 6276 22420
rect 6270 22380 6276 22392
rect 6328 22380 6334 22432
rect 9030 22420 9036 22432
rect 8991 22392 9036 22420
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 9766 22380 9772 22432
rect 9824 22420 9830 22432
rect 10321 22423 10379 22429
rect 10321 22420 10333 22423
rect 9824 22392 10333 22420
rect 9824 22380 9830 22392
rect 10321 22389 10333 22392
rect 10367 22420 10379 22423
rect 10781 22423 10839 22429
rect 10781 22420 10793 22423
rect 10367 22392 10793 22420
rect 10367 22389 10379 22392
rect 10321 22383 10379 22389
rect 10781 22389 10793 22392
rect 10827 22389 10839 22423
rect 10781 22383 10839 22389
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 12912 22420 12940 22460
rect 13357 22457 13369 22460
rect 13403 22488 13415 22491
rect 13556 22488 13584 22516
rect 13808 22491 13866 22497
rect 13808 22488 13820 22491
rect 13403 22460 13584 22488
rect 13648 22460 13820 22488
rect 13403 22457 13415 22460
rect 13357 22451 13415 22457
rect 13078 22420 13084 22432
rect 12032 22392 12940 22420
rect 12991 22392 13084 22420
rect 12032 22380 12038 22392
rect 13078 22380 13084 22392
rect 13136 22420 13142 22432
rect 13648 22420 13676 22460
rect 13808 22457 13820 22460
rect 13854 22488 13866 22491
rect 14550 22488 14556 22500
rect 13854 22460 14556 22488
rect 13854 22457 13866 22460
rect 13808 22451 13866 22457
rect 14550 22448 14556 22460
rect 14608 22448 14614 22500
rect 15930 22448 15936 22500
rect 15988 22488 15994 22500
rect 17862 22488 17868 22500
rect 15988 22460 17868 22488
rect 15988 22448 15994 22460
rect 17862 22448 17868 22460
rect 17920 22488 17926 22500
rect 18233 22491 18291 22497
rect 18233 22488 18245 22491
rect 17920 22460 18245 22488
rect 17920 22448 17926 22460
rect 18233 22457 18245 22460
rect 18279 22457 18291 22491
rect 18233 22451 18291 22457
rect 15562 22420 15568 22432
rect 13136 22392 13676 22420
rect 15523 22392 15568 22420
rect 13136 22380 13142 22392
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 18874 22420 18880 22432
rect 18835 22392 18880 22420
rect 18874 22380 18880 22392
rect 18932 22380 18938 22432
rect 20714 22380 20720 22432
rect 20772 22420 20778 22432
rect 20901 22423 20959 22429
rect 20901 22420 20913 22423
rect 20772 22392 20913 22420
rect 20772 22380 20778 22392
rect 20901 22389 20913 22392
rect 20947 22389 20959 22423
rect 22186 22420 22192 22432
rect 22147 22392 22192 22420
rect 20901 22383 20959 22389
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 23290 22420 23296 22432
rect 23251 22392 23296 22420
rect 23290 22380 23296 22392
rect 23348 22380 23354 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1670 22216 1676 22228
rect 1631 22188 1676 22216
rect 1670 22176 1676 22188
rect 1728 22176 1734 22228
rect 2130 22216 2136 22228
rect 2091 22188 2136 22216
rect 2130 22176 2136 22188
rect 2188 22216 2194 22228
rect 4706 22216 4712 22228
rect 2188 22188 2728 22216
rect 4667 22188 4712 22216
rect 2188 22176 2194 22188
rect 2700 22080 2728 22188
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 5166 22176 5172 22228
rect 5224 22216 5230 22228
rect 5445 22219 5503 22225
rect 5445 22216 5457 22219
rect 5224 22188 5457 22216
rect 5224 22176 5230 22188
rect 5445 22185 5457 22188
rect 5491 22185 5503 22219
rect 5445 22179 5503 22185
rect 6457 22219 6515 22225
rect 6457 22185 6469 22219
rect 6503 22216 6515 22219
rect 6822 22216 6828 22228
rect 6503 22188 6828 22216
rect 6503 22185 6515 22188
rect 6457 22179 6515 22185
rect 5350 22148 5356 22160
rect 5311 22120 5356 22148
rect 5350 22108 5356 22120
rect 5408 22108 5414 22160
rect 2869 22083 2927 22089
rect 2700 22052 2820 22080
rect 2222 22012 2228 22024
rect 2183 21984 2228 22012
rect 2222 21972 2228 21984
rect 2280 21972 2286 22024
rect 2409 22015 2467 22021
rect 2409 21981 2421 22015
rect 2455 22012 2467 22015
rect 2682 22012 2688 22024
rect 2455 21984 2688 22012
rect 2455 21981 2467 21984
rect 2409 21975 2467 21981
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 2792 22012 2820 22052
rect 2869 22049 2881 22083
rect 2915 22080 2927 22083
rect 3050 22080 3056 22092
rect 2915 22052 3056 22080
rect 2915 22049 2927 22052
rect 2869 22043 2927 22049
rect 3050 22040 3056 22052
rect 3108 22040 3114 22092
rect 5460 22080 5488 22179
rect 6822 22176 6828 22188
rect 6880 22216 6886 22228
rect 6917 22219 6975 22225
rect 6917 22216 6929 22219
rect 6880 22188 6929 22216
rect 6880 22176 6886 22188
rect 6917 22185 6929 22188
rect 6963 22185 6975 22219
rect 7558 22216 7564 22228
rect 7519 22188 7564 22216
rect 6917 22179 6975 22185
rect 7558 22176 7564 22188
rect 7616 22216 7622 22228
rect 7929 22219 7987 22225
rect 7929 22216 7941 22219
rect 7616 22188 7941 22216
rect 7616 22176 7622 22188
rect 7929 22185 7941 22188
rect 7975 22185 7987 22219
rect 8662 22216 8668 22228
rect 8575 22188 8668 22216
rect 7929 22179 7987 22185
rect 8662 22176 8668 22188
rect 8720 22216 8726 22228
rect 9030 22216 9036 22228
rect 8720 22188 9036 22216
rect 8720 22176 8726 22188
rect 9030 22176 9036 22188
rect 9088 22176 9094 22228
rect 9677 22219 9735 22225
rect 9677 22185 9689 22219
rect 9723 22216 9735 22219
rect 9766 22216 9772 22228
rect 9723 22188 9772 22216
rect 9723 22185 9735 22188
rect 9677 22179 9735 22185
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 10689 22219 10747 22225
rect 10689 22185 10701 22219
rect 10735 22216 10747 22219
rect 10778 22216 10784 22228
rect 10735 22188 10784 22216
rect 10735 22185 10747 22188
rect 10689 22179 10747 22185
rect 10778 22176 10784 22188
rect 10836 22176 10842 22228
rect 12710 22176 12716 22228
rect 12768 22216 12774 22228
rect 12897 22219 12955 22225
rect 12897 22216 12909 22219
rect 12768 22188 12909 22216
rect 12768 22176 12774 22188
rect 12897 22185 12909 22188
rect 12943 22185 12955 22219
rect 12897 22179 12955 22185
rect 5997 22083 6055 22089
rect 5997 22080 6009 22083
rect 5460 22052 6009 22080
rect 5997 22049 6009 22052
rect 6043 22049 6055 22083
rect 8110 22080 8116 22092
rect 8071 22052 8116 22080
rect 5997 22043 6055 22049
rect 8110 22040 8116 22052
rect 8168 22040 8174 22092
rect 9493 22083 9551 22089
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9582 22080 9588 22092
rect 9539 22052 9588 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 10505 22083 10563 22089
rect 10505 22049 10517 22083
rect 10551 22080 10563 22083
rect 10686 22080 10692 22092
rect 10551 22052 10692 22080
rect 10551 22049 10563 22052
rect 10505 22043 10563 22049
rect 10686 22040 10692 22052
rect 10744 22040 10750 22092
rect 11054 22080 11060 22092
rect 11015 22052 11060 22080
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 3605 22015 3663 22021
rect 3605 22012 3617 22015
rect 2792 21984 3617 22012
rect 3605 21981 3617 21984
rect 3651 21981 3663 22015
rect 3605 21975 3663 21981
rect 4341 22015 4399 22021
rect 4341 21981 4353 22015
rect 4387 22012 4399 22015
rect 5537 22015 5595 22021
rect 5537 22012 5549 22015
rect 4387 21984 5549 22012
rect 4387 21981 4399 21984
rect 4341 21975 4399 21981
rect 5537 21981 5549 21984
rect 5583 22012 5595 22015
rect 6178 22012 6184 22024
rect 5583 21984 6184 22012
rect 5583 21981 5595 21984
rect 5537 21975 5595 21981
rect 6178 21972 6184 21984
rect 6236 21972 6242 22024
rect 6730 21972 6736 22024
rect 6788 22012 6794 22024
rect 7009 22015 7067 22021
rect 7009 22012 7021 22015
rect 6788 21984 7021 22012
rect 6788 21972 6794 21984
rect 7009 21981 7021 21984
rect 7055 21981 7067 22015
rect 7009 21975 7067 21981
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22012 7251 22015
rect 7834 22012 7840 22024
rect 7239 21984 7840 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 7834 21972 7840 21984
rect 7892 22012 7898 22024
rect 8662 22012 8668 22024
rect 7892 21984 8668 22012
rect 7892 21972 7898 21984
rect 8662 21972 8668 21984
rect 8720 21972 8726 22024
rect 10962 21972 10968 22024
rect 11020 22012 11026 22024
rect 11149 22015 11207 22021
rect 11149 22012 11161 22015
rect 11020 21984 11161 22012
rect 11020 21972 11026 21984
rect 11149 21981 11161 21984
rect 11195 21981 11207 22015
rect 11149 21975 11207 21981
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 22012 11391 22015
rect 12066 22012 12072 22024
rect 11379 21984 12072 22012
rect 11379 21981 11391 21984
rect 11333 21975 11391 21981
rect 10778 21904 10784 21956
rect 10836 21944 10842 21956
rect 11348 21944 11376 21975
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 12989 22015 13047 22021
rect 12989 22012 13001 22015
rect 12676 21984 13001 22012
rect 12676 21972 12682 21984
rect 12989 21981 13001 21984
rect 13035 21981 13047 22015
rect 12989 21975 13047 21981
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 22012 13231 22015
rect 13722 22012 13728 22024
rect 13219 21984 13728 22012
rect 13219 21981 13231 21984
rect 13173 21975 13231 21981
rect 10836 21916 11376 21944
rect 10836 21904 10842 21916
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 13188 21944 13216 21975
rect 13722 21972 13728 21984
rect 13780 21972 13786 22024
rect 12308 21916 13216 21944
rect 12308 21904 12314 21916
rect 1765 21879 1823 21885
rect 1765 21845 1777 21879
rect 1811 21876 1823 21879
rect 2130 21876 2136 21888
rect 1811 21848 2136 21876
rect 1811 21845 1823 21848
rect 1765 21839 1823 21845
rect 2130 21836 2136 21848
rect 2188 21836 2194 21888
rect 3234 21836 3240 21888
rect 3292 21876 3298 21888
rect 3329 21879 3387 21885
rect 3329 21876 3341 21879
rect 3292 21848 3341 21876
rect 3292 21836 3298 21848
rect 3329 21845 3341 21848
rect 3375 21876 3387 21879
rect 3418 21876 3424 21888
rect 3375 21848 3424 21876
rect 3375 21845 3387 21848
rect 3329 21839 3387 21845
rect 3418 21836 3424 21848
rect 3476 21836 3482 21888
rect 4982 21876 4988 21888
rect 4943 21848 4988 21876
rect 4982 21836 4988 21848
rect 5040 21836 5046 21888
rect 6549 21879 6607 21885
rect 6549 21845 6561 21879
rect 6595 21876 6607 21879
rect 6638 21876 6644 21888
rect 6595 21848 6644 21876
rect 6595 21845 6607 21848
rect 6549 21839 6607 21845
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 8297 21879 8355 21885
rect 8297 21845 8309 21879
rect 8343 21876 8355 21879
rect 8386 21876 8392 21888
rect 8343 21848 8392 21876
rect 8343 21845 8355 21848
rect 8297 21839 8355 21845
rect 8386 21836 8392 21848
rect 8444 21836 8450 21888
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 13170 21876 13176 21888
rect 12575 21848 13176 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 13538 21876 13544 21888
rect 13499 21848 13544 21876
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 2038 21672 2044 21684
rect 1999 21644 2044 21672
rect 2038 21632 2044 21644
rect 2096 21632 2102 21684
rect 2409 21675 2467 21681
rect 2409 21641 2421 21675
rect 2455 21672 2467 21675
rect 2682 21672 2688 21684
rect 2455 21644 2688 21672
rect 2455 21641 2467 21644
rect 2409 21635 2467 21641
rect 2682 21632 2688 21644
rect 2740 21632 2746 21684
rect 4341 21675 4399 21681
rect 4341 21641 4353 21675
rect 4387 21672 4399 21675
rect 5350 21672 5356 21684
rect 4387 21644 5356 21672
rect 4387 21641 4399 21644
rect 4341 21635 4399 21641
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 6546 21672 6552 21684
rect 6507 21644 6552 21672
rect 6546 21632 6552 21644
rect 6604 21632 6610 21684
rect 6822 21672 6828 21684
rect 6783 21644 6828 21672
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 7834 21672 7840 21684
rect 7795 21644 7840 21672
rect 7834 21632 7840 21644
rect 7892 21632 7898 21684
rect 11054 21672 11060 21684
rect 11015 21644 11060 21672
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 12250 21672 12256 21684
rect 12211 21644 12256 21672
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 12710 21672 12716 21684
rect 12671 21644 12716 21672
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 14550 21672 14556 21684
rect 14511 21644 14556 21672
rect 14550 21632 14556 21644
rect 14608 21632 14614 21684
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21536 3203 21539
rect 3694 21536 3700 21548
rect 3191 21508 3700 21536
rect 3191 21505 3203 21508
rect 3145 21499 3203 21505
rect 3694 21496 3700 21508
rect 3752 21496 3758 21548
rect 3789 21539 3847 21545
rect 3789 21505 3801 21539
rect 3835 21505 3847 21539
rect 5718 21536 5724 21548
rect 5679 21508 5724 21536
rect 3789 21499 3847 21505
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 2038 21468 2044 21480
rect 1443 21440 2044 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2038 21428 2044 21440
rect 2096 21428 2102 21480
rect 3804 21468 3832 21499
rect 5718 21496 5724 21508
rect 5776 21496 5782 21548
rect 6564 21536 6592 21632
rect 10781 21607 10839 21613
rect 10781 21573 10793 21607
rect 10827 21604 10839 21607
rect 10962 21604 10968 21616
rect 10827 21576 10968 21604
rect 10827 21573 10839 21576
rect 10781 21567 10839 21573
rect 10962 21564 10968 21576
rect 11020 21564 11026 21616
rect 11885 21607 11943 21613
rect 11885 21573 11897 21607
rect 11931 21604 11943 21607
rect 12618 21604 12624 21616
rect 11931 21576 12624 21604
rect 11931 21573 11943 21576
rect 11885 21567 11943 21573
rect 12618 21564 12624 21576
rect 12676 21564 12682 21616
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 6564 21508 7297 21536
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7466 21536 7472 21548
rect 7427 21508 7472 21536
rect 7285 21499 7343 21505
rect 7466 21496 7472 21508
rect 7524 21496 7530 21548
rect 11790 21496 11796 21548
rect 11848 21536 11854 21548
rect 11848 21508 13308 21536
rect 11848 21496 11854 21508
rect 2884 21440 3832 21468
rect 5077 21471 5135 21477
rect 2884 21344 2912 21440
rect 5077 21437 5089 21471
rect 5123 21468 5135 21471
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 5123 21440 5641 21468
rect 5123 21437 5135 21440
rect 5077 21431 5135 21437
rect 5629 21437 5641 21440
rect 5675 21468 5687 21471
rect 5994 21468 6000 21480
rect 5675 21440 6000 21468
rect 5675 21437 5687 21440
rect 5629 21431 5687 21437
rect 5994 21428 6000 21440
rect 6052 21428 6058 21480
rect 6273 21471 6331 21477
rect 6273 21437 6285 21471
rect 6319 21468 6331 21471
rect 6914 21468 6920 21480
rect 6319 21440 6920 21468
rect 6319 21437 6331 21440
rect 6273 21431 6331 21437
rect 6914 21428 6920 21440
rect 6972 21468 6978 21480
rect 7193 21471 7251 21477
rect 7193 21468 7205 21471
rect 6972 21440 7205 21468
rect 6972 21428 6978 21440
rect 7193 21437 7205 21440
rect 7239 21437 7251 21471
rect 8573 21471 8631 21477
rect 8573 21468 8585 21471
rect 7193 21431 7251 21437
rect 8404 21440 8585 21468
rect 3418 21360 3424 21412
rect 3476 21400 3482 21412
rect 3605 21403 3663 21409
rect 3605 21400 3617 21403
rect 3476 21372 3617 21400
rect 3476 21360 3482 21372
rect 3605 21369 3617 21372
rect 3651 21400 3663 21403
rect 4709 21403 4767 21409
rect 4709 21400 4721 21403
rect 3651 21372 4721 21400
rect 3651 21369 3663 21372
rect 3605 21363 3663 21369
rect 4709 21369 4721 21372
rect 4755 21400 4767 21403
rect 8404 21400 8432 21440
rect 8573 21437 8585 21440
rect 8619 21437 8631 21471
rect 8573 21431 8631 21437
rect 8662 21428 8668 21480
rect 8720 21468 8726 21480
rect 8829 21471 8887 21477
rect 8829 21468 8841 21471
rect 8720 21440 8841 21468
rect 8720 21428 8726 21440
rect 8829 21437 8841 21440
rect 8875 21437 8887 21471
rect 13173 21471 13231 21477
rect 13173 21468 13185 21471
rect 8829 21431 8887 21437
rect 13004 21440 13185 21468
rect 9490 21400 9496 21412
rect 4755 21372 5580 21400
rect 4755 21369 4767 21372
rect 4709 21363 4767 21369
rect 5552 21344 5580 21372
rect 8404 21372 9496 21400
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 2038 21332 2044 21344
rect 1912 21304 2044 21332
rect 1912 21292 1918 21304
rect 2038 21292 2044 21304
rect 2096 21292 2102 21344
rect 2777 21335 2835 21341
rect 2777 21301 2789 21335
rect 2823 21332 2835 21335
rect 2866 21332 2872 21344
rect 2823 21304 2872 21332
rect 2823 21301 2835 21304
rect 2777 21295 2835 21301
rect 2866 21292 2872 21304
rect 2924 21292 2930 21344
rect 3234 21332 3240 21344
rect 3195 21304 3240 21332
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 5169 21335 5227 21341
rect 5169 21301 5181 21335
rect 5215 21332 5227 21335
rect 5258 21332 5264 21344
rect 5215 21304 5264 21332
rect 5215 21301 5227 21304
rect 5169 21295 5227 21301
rect 5258 21292 5264 21304
rect 5316 21292 5322 21344
rect 5534 21332 5540 21344
rect 5495 21304 5540 21332
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 8018 21292 8024 21344
rect 8076 21332 8082 21344
rect 8404 21341 8432 21372
rect 9490 21360 9496 21372
rect 9548 21360 9554 21412
rect 8389 21335 8447 21341
rect 8389 21332 8401 21335
rect 8076 21304 8401 21332
rect 8076 21292 8082 21304
rect 8389 21301 8401 21304
rect 8435 21301 8447 21335
rect 9950 21332 9956 21344
rect 9911 21304 9956 21332
rect 8389 21295 8447 21301
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 11330 21332 11336 21344
rect 11291 21304 11336 21332
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 13004 21341 13032 21440
rect 13173 21437 13185 21440
rect 13219 21437 13231 21471
rect 13173 21431 13231 21437
rect 13280 21400 13308 21508
rect 13440 21403 13498 21409
rect 13440 21400 13452 21403
rect 13280 21372 13452 21400
rect 13440 21369 13452 21372
rect 13486 21400 13498 21403
rect 13538 21400 13544 21412
rect 13486 21372 13544 21400
rect 13486 21369 13498 21372
rect 13440 21363 13498 21369
rect 13538 21360 13544 21372
rect 13596 21400 13602 21412
rect 14090 21400 14096 21412
rect 13596 21372 14096 21400
rect 13596 21360 13602 21372
rect 14090 21360 14096 21372
rect 14148 21360 14154 21412
rect 12989 21335 13047 21341
rect 12989 21332 13001 21335
rect 12768 21304 13001 21332
rect 12768 21292 12774 21304
rect 12989 21301 13001 21304
rect 13035 21301 13047 21335
rect 12989 21295 13047 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 3421 21131 3479 21137
rect 3421 21128 3433 21131
rect 2280 21100 3433 21128
rect 2280 21088 2286 21100
rect 3421 21097 3433 21100
rect 3467 21097 3479 21131
rect 3421 21091 3479 21097
rect 6457 21131 6515 21137
rect 6457 21097 6469 21131
rect 6503 21128 6515 21131
rect 6730 21128 6736 21140
rect 6503 21100 6736 21128
rect 6503 21097 6515 21100
rect 6457 21091 6515 21097
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 9950 21088 9956 21140
rect 10008 21128 10014 21140
rect 10321 21131 10379 21137
rect 10321 21128 10333 21131
rect 10008 21100 10333 21128
rect 10008 21088 10014 21100
rect 10321 21097 10333 21100
rect 10367 21097 10379 21131
rect 10778 21128 10784 21140
rect 10739 21100 10784 21128
rect 10321 21091 10379 21097
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11330 21088 11336 21140
rect 11388 21128 11394 21140
rect 11517 21131 11575 21137
rect 11517 21128 11529 21131
rect 11388 21100 11529 21128
rect 11388 21088 11394 21100
rect 11517 21097 11529 21100
rect 11563 21097 11575 21131
rect 14090 21128 14096 21140
rect 14051 21100 14096 21128
rect 11517 21091 11575 21097
rect 14090 21088 14096 21100
rect 14148 21088 14154 21140
rect 1486 21020 1492 21072
rect 1544 21060 1550 21072
rect 1946 21060 1952 21072
rect 1544 21032 1952 21060
rect 1544 21020 1550 21032
rect 1946 21020 1952 21032
rect 2004 21020 2010 21072
rect 6270 21020 6276 21072
rect 6328 21060 6334 21072
rect 6816 21063 6874 21069
rect 6816 21060 6828 21063
rect 6328 21032 6828 21060
rect 6328 21020 6334 21032
rect 6816 21029 6828 21032
rect 6862 21060 6874 21063
rect 6914 21060 6920 21072
rect 6862 21032 6920 21060
rect 6862 21029 6874 21032
rect 6816 21023 6874 21029
rect 6914 21020 6920 21032
rect 6972 21020 6978 21072
rect 12980 21063 13038 21069
rect 12980 21029 12992 21063
rect 13026 21060 13038 21063
rect 13078 21060 13084 21072
rect 13026 21032 13084 21060
rect 13026 21029 13038 21032
rect 12980 21023 13038 21029
rect 13078 21020 13084 21032
rect 13136 21020 13142 21072
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 3142 20992 3148 21004
rect 2547 20964 3148 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 4332 20995 4390 21001
rect 4332 20992 4344 20995
rect 4028 20964 4344 20992
rect 4028 20952 4034 20964
rect 4332 20961 4344 20964
rect 4378 20992 4390 20995
rect 4378 20964 5488 20992
rect 4378 20961 4390 20964
rect 4332 20955 4390 20961
rect 5460 20936 5488 20964
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 9732 20964 9777 20992
rect 9732 20952 9738 20964
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 2682 20856 2688 20868
rect 2643 20828 2688 20856
rect 2682 20816 2688 20828
rect 2740 20816 2746 20868
rect 2222 20748 2228 20800
rect 2280 20788 2286 20800
rect 2317 20791 2375 20797
rect 2317 20788 2329 20791
rect 2280 20760 2329 20788
rect 2280 20748 2286 20760
rect 2317 20757 2329 20760
rect 2363 20757 2375 20791
rect 3786 20788 3792 20800
rect 3747 20760 3792 20788
rect 2317 20751 2375 20757
rect 3786 20748 3792 20760
rect 3844 20748 3850 20800
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 4080 20788 4108 20887
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 5644 20896 6561 20924
rect 5644 20856 5672 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 5000 20828 5672 20856
rect 5000 20788 5028 20828
rect 5718 20816 5724 20868
rect 5776 20816 5782 20868
rect 4028 20760 5028 20788
rect 4028 20748 4034 20760
rect 5074 20748 5080 20800
rect 5132 20788 5138 20800
rect 5445 20791 5503 20797
rect 5445 20788 5457 20791
rect 5132 20760 5457 20788
rect 5132 20748 5138 20760
rect 5445 20757 5457 20760
rect 5491 20788 5503 20791
rect 5736 20788 5764 20816
rect 5997 20791 6055 20797
rect 5997 20788 6009 20791
rect 5491 20760 6009 20788
rect 5491 20757 5503 20760
rect 5445 20751 5503 20757
rect 5997 20757 6009 20760
rect 6043 20757 6055 20791
rect 6564 20788 6592 20887
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 11609 20927 11667 20933
rect 11609 20924 11621 20927
rect 11112 20896 11621 20924
rect 11112 20884 11118 20896
rect 11609 20893 11621 20896
rect 11655 20893 11667 20927
rect 11790 20924 11796 20936
rect 11751 20896 11796 20924
rect 11609 20887 11667 20893
rect 7650 20816 7656 20868
rect 7708 20856 7714 20868
rect 8110 20856 8116 20868
rect 7708 20828 8116 20856
rect 7708 20816 7714 20828
rect 8110 20816 8116 20828
rect 8168 20856 8174 20868
rect 8849 20859 8907 20865
rect 8849 20856 8861 20859
rect 8168 20828 8861 20856
rect 8168 20816 8174 20828
rect 8849 20825 8861 20828
rect 8895 20825 8907 20859
rect 11624 20856 11652 20887
rect 11790 20884 11796 20896
rect 11848 20884 11854 20936
rect 11974 20884 11980 20936
rect 12032 20924 12038 20936
rect 12710 20924 12716 20936
rect 12032 20896 12716 20924
rect 12032 20884 12038 20896
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 12342 20856 12348 20868
rect 11624 20828 12348 20856
rect 8849 20819 8907 20825
rect 12342 20816 12348 20828
rect 12400 20816 12406 20868
rect 6730 20788 6736 20800
rect 6564 20760 6736 20788
rect 5997 20751 6055 20757
rect 6730 20748 6736 20760
rect 6788 20748 6794 20800
rect 7834 20748 7840 20800
rect 7892 20788 7898 20800
rect 7929 20791 7987 20797
rect 7929 20788 7941 20791
rect 7892 20760 7941 20788
rect 7892 20748 7898 20760
rect 7929 20757 7941 20760
rect 7975 20757 7987 20791
rect 8570 20788 8576 20800
rect 8531 20760 8576 20788
rect 7929 20751 7987 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 9861 20791 9919 20797
rect 9861 20757 9873 20791
rect 9907 20788 9919 20791
rect 10134 20788 10140 20800
rect 9907 20760 10140 20788
rect 9907 20757 9919 20760
rect 9861 20751 9919 20757
rect 10134 20748 10140 20760
rect 10192 20748 10198 20800
rect 11149 20791 11207 20797
rect 11149 20757 11161 20791
rect 11195 20788 11207 20791
rect 11698 20788 11704 20800
rect 11195 20760 11704 20788
rect 11195 20757 11207 20760
rect 11149 20751 11207 20757
rect 11698 20748 11704 20760
rect 11756 20748 11762 20800
rect 12526 20788 12532 20800
rect 12487 20760 12532 20788
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1394 20544 1400 20596
rect 1452 20584 1458 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1452 20556 1593 20584
rect 1452 20544 1458 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 3329 20587 3387 20593
rect 3329 20584 3341 20587
rect 3016 20556 3341 20584
rect 3016 20544 3022 20556
rect 3329 20553 3341 20556
rect 3375 20553 3387 20587
rect 3970 20584 3976 20596
rect 3931 20556 3976 20584
rect 3329 20547 3387 20553
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 5534 20584 5540 20596
rect 5495 20556 5540 20584
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 6086 20544 6092 20596
rect 6144 20584 6150 20596
rect 6181 20587 6239 20593
rect 6181 20584 6193 20587
rect 6144 20556 6193 20584
rect 6144 20544 6150 20556
rect 6181 20553 6193 20556
rect 6227 20553 6239 20587
rect 6181 20547 6239 20553
rect 1946 20448 1952 20460
rect 1907 20420 1952 20448
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 4890 20408 4896 20460
rect 4948 20448 4954 20460
rect 4985 20451 5043 20457
rect 4985 20448 4997 20451
rect 4948 20420 4997 20448
rect 4948 20408 4954 20420
rect 4985 20417 4997 20420
rect 5031 20417 5043 20451
rect 4985 20411 5043 20417
rect 2222 20389 2228 20392
rect 2216 20380 2228 20389
rect 2183 20352 2228 20380
rect 2216 20343 2228 20352
rect 2222 20340 2228 20343
rect 2280 20340 2286 20392
rect 4798 20380 4804 20392
rect 4759 20352 4804 20380
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 6196 20380 6224 20547
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7285 20587 7343 20593
rect 7285 20584 7297 20587
rect 6972 20556 7297 20584
rect 6972 20544 6978 20556
rect 7285 20553 7297 20556
rect 7331 20553 7343 20587
rect 7285 20547 7343 20553
rect 9861 20587 9919 20593
rect 9861 20553 9873 20587
rect 9907 20584 9919 20587
rect 11054 20584 11060 20596
rect 9907 20556 11060 20584
rect 9907 20553 9919 20556
rect 9861 20547 9919 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 11330 20584 11336 20596
rect 11291 20556 11336 20584
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 11885 20587 11943 20593
rect 11885 20553 11897 20587
rect 11931 20584 11943 20587
rect 11974 20584 11980 20596
rect 11931 20556 11980 20584
rect 11931 20553 11943 20556
rect 11885 20547 11943 20553
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 13814 20584 13820 20596
rect 12492 20556 12537 20584
rect 13775 20556 13820 20584
rect 12492 20544 12498 20556
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 9398 20476 9404 20528
rect 9456 20516 9462 20528
rect 9950 20516 9956 20528
rect 9456 20488 9956 20516
rect 9456 20476 9462 20488
rect 9950 20476 9956 20488
rect 10008 20516 10014 20528
rect 10008 20488 10916 20516
rect 10008 20476 10014 20488
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20448 10287 20451
rect 10778 20448 10784 20460
rect 10275 20420 10784 20448
rect 10275 20417 10287 20420
rect 10229 20411 10287 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 10888 20457 10916 20488
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 12860 20488 12940 20516
rect 12860 20476 12866 20488
rect 12912 20457 12940 20488
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20448 12311 20451
rect 12897 20451 12955 20457
rect 12897 20448 12909 20451
rect 12299 20420 12909 20448
rect 12299 20417 12311 20420
rect 12253 20411 12311 20417
rect 12897 20417 12909 20420
rect 12943 20417 12955 20451
rect 13078 20448 13084 20460
rect 13039 20420 13084 20448
rect 12897 20411 12955 20417
rect 13078 20408 13084 20420
rect 13136 20408 13142 20460
rect 14550 20448 14556 20460
rect 14511 20420 14556 20448
rect 14550 20408 14556 20420
rect 14608 20448 14614 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14608 20420 15025 20448
rect 14608 20408 14614 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 8110 20389 8116 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6196 20352 6837 20380
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20349 7895 20383
rect 8104 20380 8116 20389
rect 8071 20352 8116 20380
rect 7837 20343 7895 20349
rect 8104 20343 8116 20352
rect 1946 20272 1952 20324
rect 2004 20312 2010 20324
rect 3970 20312 3976 20324
rect 2004 20284 3976 20312
rect 2004 20272 2010 20284
rect 3970 20272 3976 20284
rect 4028 20272 4034 20324
rect 4062 20272 4068 20324
rect 4120 20312 4126 20324
rect 4341 20315 4399 20321
rect 4341 20312 4353 20315
rect 4120 20284 4353 20312
rect 4120 20272 4126 20284
rect 4341 20281 4353 20284
rect 4387 20312 4399 20315
rect 4893 20315 4951 20321
rect 4893 20312 4905 20315
rect 4387 20284 4905 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 4893 20281 4905 20284
rect 4939 20312 4951 20315
rect 5442 20312 5448 20324
rect 4939 20284 5448 20312
rect 4939 20281 4951 20284
rect 4893 20275 4951 20281
rect 5442 20272 5448 20284
rect 5500 20272 5506 20324
rect 7653 20315 7711 20321
rect 7653 20312 7665 20315
rect 6748 20284 7665 20312
rect 6748 20256 6776 20284
rect 7653 20281 7665 20284
rect 7699 20312 7711 20315
rect 7852 20312 7880 20343
rect 8110 20340 8116 20343
rect 8168 20340 8174 20392
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 12584 20352 12817 20380
rect 12584 20340 12590 20352
rect 12805 20349 12817 20352
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 13872 20352 14473 20380
rect 13872 20340 13878 20352
rect 14461 20349 14473 20352
rect 14507 20349 14519 20383
rect 14461 20343 14519 20349
rect 8018 20312 8024 20324
rect 7699 20284 8024 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 8018 20272 8024 20284
rect 8076 20272 8082 20324
rect 10686 20312 10692 20324
rect 10599 20284 10692 20312
rect 10686 20272 10692 20284
rect 10744 20312 10750 20324
rect 13449 20315 13507 20321
rect 13449 20312 13461 20315
rect 10744 20284 13461 20312
rect 10744 20272 10750 20284
rect 13449 20281 13461 20284
rect 13495 20312 13507 20315
rect 14369 20315 14427 20321
rect 14369 20312 14381 20315
rect 13495 20284 14381 20312
rect 13495 20281 13507 20284
rect 13449 20275 13507 20281
rect 14369 20281 14381 20284
rect 14415 20281 14427 20315
rect 14369 20275 14427 20281
rect 4430 20244 4436 20256
rect 4391 20216 4436 20244
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 6641 20247 6699 20253
rect 6641 20213 6653 20247
rect 6687 20244 6699 20247
rect 6730 20244 6736 20256
rect 6687 20216 6736 20244
rect 6687 20213 6699 20216
rect 6641 20207 6699 20213
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 7006 20244 7012 20256
rect 6967 20216 7012 20244
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 9214 20244 9220 20256
rect 9175 20216 9220 20244
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10321 20247 10379 20253
rect 10321 20244 10333 20247
rect 9824 20216 10333 20244
rect 9824 20204 9830 20216
rect 10321 20213 10333 20216
rect 10367 20213 10379 20247
rect 13998 20244 14004 20256
rect 13959 20216 14004 20244
rect 10321 20207 10379 20213
rect 13998 20204 14004 20216
rect 14056 20204 14062 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2222 20000 2228 20052
rect 2280 20040 2286 20052
rect 2590 20040 2596 20052
rect 2280 20012 2596 20040
rect 2280 20000 2286 20012
rect 2590 20000 2596 20012
rect 2648 20040 2654 20052
rect 2869 20043 2927 20049
rect 2869 20040 2881 20043
rect 2648 20012 2881 20040
rect 2648 20000 2654 20012
rect 2869 20009 2881 20012
rect 2915 20009 2927 20043
rect 2869 20003 2927 20009
rect 3234 20000 3240 20052
rect 3292 20040 3298 20052
rect 3421 20043 3479 20049
rect 3421 20040 3433 20043
rect 3292 20012 3433 20040
rect 3292 20000 3298 20012
rect 3421 20009 3433 20012
rect 3467 20009 3479 20043
rect 3421 20003 3479 20009
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 4798 20040 4804 20052
rect 4571 20012 4804 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 4798 20000 4804 20012
rect 4856 20040 4862 20052
rect 5353 20043 5411 20049
rect 5353 20040 5365 20043
rect 4856 20012 5365 20040
rect 4856 20000 4862 20012
rect 5353 20009 5365 20012
rect 5399 20009 5411 20043
rect 5353 20003 5411 20009
rect 5442 20000 5448 20052
rect 5500 20040 5506 20052
rect 8021 20043 8079 20049
rect 5500 20012 5545 20040
rect 5500 20000 5506 20012
rect 8021 20009 8033 20043
rect 8067 20040 8079 20043
rect 8110 20040 8116 20052
rect 8067 20012 8116 20040
rect 8067 20009 8079 20012
rect 8021 20003 8079 20009
rect 8110 20000 8116 20012
rect 8168 20040 8174 20052
rect 8294 20040 8300 20052
rect 8168 20012 8300 20040
rect 8168 20000 8174 20012
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 10413 20043 10471 20049
rect 10413 20009 10425 20043
rect 10459 20040 10471 20043
rect 10686 20040 10692 20052
rect 10459 20012 10692 20040
rect 10459 20009 10471 20012
rect 10413 20003 10471 20009
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 11790 20040 11796 20052
rect 11751 20012 11796 20040
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12253 20043 12311 20049
rect 12253 20009 12265 20043
rect 12299 20040 12311 20043
rect 13078 20040 13084 20052
rect 12299 20012 13084 20040
rect 12299 20009 12311 20012
rect 12253 20003 12311 20009
rect 13078 20000 13084 20012
rect 13136 20040 13142 20052
rect 13725 20043 13783 20049
rect 13725 20040 13737 20043
rect 13136 20012 13737 20040
rect 13136 20000 13142 20012
rect 13725 20009 13737 20012
rect 13771 20040 13783 20043
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 13771 20012 14289 20040
rect 13771 20009 13783 20012
rect 13725 20003 13783 20009
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 1670 19972 1676 19984
rect 1504 19944 1676 19972
rect 1504 19913 1532 19944
rect 1670 19932 1676 19944
rect 1728 19972 1734 19984
rect 1946 19972 1952 19984
rect 1728 19944 1952 19972
rect 1728 19932 1734 19944
rect 1946 19932 1952 19944
rect 2004 19932 2010 19984
rect 6178 19932 6184 19984
rect 6236 19972 6242 19984
rect 6886 19975 6944 19981
rect 6886 19972 6898 19975
rect 6236 19944 6898 19972
rect 6236 19932 6242 19944
rect 6886 19941 6898 19944
rect 6932 19972 6944 19975
rect 7834 19972 7840 19984
rect 6932 19944 7840 19972
rect 6932 19941 6944 19944
rect 6886 19935 6944 19941
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 1489 19907 1547 19913
rect 1489 19873 1501 19907
rect 1535 19873 1547 19907
rect 1489 19867 1547 19873
rect 1756 19907 1814 19913
rect 1756 19873 1768 19907
rect 1802 19904 1814 19907
rect 2958 19904 2964 19916
rect 1802 19876 2964 19904
rect 1802 19873 1814 19876
rect 1756 19867 1814 19873
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 6730 19904 6736 19916
rect 6687 19876 6736 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 9677 19907 9735 19913
rect 9677 19873 9689 19907
rect 9723 19904 9735 19907
rect 9858 19904 9864 19916
rect 9723 19876 9864 19904
rect 9723 19873 9735 19876
rect 9677 19867 9735 19873
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11149 19907 11207 19913
rect 11149 19904 11161 19907
rect 11112 19876 11161 19904
rect 11112 19864 11118 19876
rect 11149 19873 11161 19876
rect 11195 19873 11207 19907
rect 11149 19867 11207 19873
rect 11974 19864 11980 19916
rect 12032 19904 12038 19916
rect 12342 19904 12348 19916
rect 12032 19876 12348 19904
rect 12032 19864 12038 19876
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12618 19913 12624 19916
rect 12612 19904 12624 19913
rect 12579 19876 12624 19904
rect 12612 19867 12624 19876
rect 12618 19864 12624 19867
rect 12676 19864 12682 19916
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19805 5595 19839
rect 11238 19836 11244 19848
rect 11199 19808 11244 19836
rect 5537 19799 5595 19805
rect 5074 19728 5080 19780
rect 5132 19768 5138 19780
rect 5552 19768 5580 19799
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11422 19836 11428 19848
rect 11383 19808 11428 19836
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 15286 19836 15292 19848
rect 15247 19808 15292 19836
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 5132 19740 5580 19768
rect 5132 19728 5138 19740
rect 9674 19728 9680 19780
rect 9732 19728 9738 19780
rect 3142 19660 3148 19712
rect 3200 19700 3206 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3200 19672 3801 19700
rect 3200 19660 3206 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 4890 19700 4896 19712
rect 4851 19672 4896 19700
rect 3789 19663 3847 19669
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 4985 19703 5043 19709
rect 4985 19669 4997 19703
rect 5031 19700 5043 19703
rect 5166 19700 5172 19712
rect 5031 19672 5172 19700
rect 5031 19669 5043 19672
rect 4985 19663 5043 19669
rect 5166 19660 5172 19672
rect 5224 19700 5230 19712
rect 5997 19703 6055 19709
rect 5997 19700 6009 19703
rect 5224 19672 6009 19700
rect 5224 19660 5230 19672
rect 5997 19669 6009 19672
rect 6043 19669 6055 19703
rect 5997 19663 6055 19669
rect 9306 19660 9312 19712
rect 9364 19700 9370 19712
rect 9401 19703 9459 19709
rect 9401 19700 9413 19703
rect 9364 19672 9413 19700
rect 9364 19660 9370 19672
rect 9401 19669 9413 19672
rect 9447 19700 9459 19703
rect 9692 19700 9720 19728
rect 9447 19672 9720 19700
rect 9861 19703 9919 19709
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 9861 19669 9873 19703
rect 9907 19700 9919 19703
rect 10134 19700 10140 19712
rect 9907 19672 10140 19700
rect 9907 19669 9919 19672
rect 9861 19663 9919 19669
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 10778 19700 10784 19712
rect 10739 19672 10784 19700
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2590 19496 2596 19508
rect 2551 19468 2596 19496
rect 2590 19456 2596 19468
rect 2648 19456 2654 19508
rect 2958 19496 2964 19508
rect 2919 19468 2964 19496
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 3142 19496 3148 19508
rect 3103 19468 3148 19496
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 4709 19499 4767 19505
rect 4709 19465 4721 19499
rect 4755 19496 4767 19499
rect 4798 19496 4804 19508
rect 4755 19468 4804 19496
rect 4755 19465 4767 19468
rect 4709 19459 4767 19465
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 10042 19496 10048 19508
rect 9824 19468 10048 19496
rect 9824 19456 9830 19468
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 11422 19496 11428 19508
rect 11335 19468 11428 19496
rect 11422 19456 11428 19468
rect 11480 19496 11486 19508
rect 11885 19499 11943 19505
rect 11885 19496 11897 19499
rect 11480 19468 11897 19496
rect 11480 19456 11486 19468
rect 11885 19465 11897 19468
rect 11931 19496 11943 19499
rect 12618 19496 12624 19508
rect 11931 19468 12624 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 12618 19456 12624 19468
rect 12676 19496 12682 19508
rect 13817 19499 13875 19505
rect 13817 19496 13829 19499
rect 12676 19468 13829 19496
rect 12676 19456 12682 19468
rect 13817 19465 13829 19468
rect 13863 19465 13875 19499
rect 13817 19459 13875 19465
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 2608 19360 2636 19456
rect 2976 19428 3004 19456
rect 2976 19400 3740 19428
rect 2271 19332 2636 19360
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 3234 19320 3240 19372
rect 3292 19360 3298 19372
rect 3712 19369 3740 19400
rect 3605 19363 3663 19369
rect 3605 19360 3617 19363
rect 3292 19332 3617 19360
rect 3292 19320 3298 19332
rect 3605 19329 3617 19332
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 4430 19360 4436 19372
rect 3697 19323 3755 19329
rect 4080 19332 4436 19360
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 3142 19292 3148 19304
rect 2087 19264 3148 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 3510 19292 3516 19304
rect 3423 19264 3516 19292
rect 3510 19252 3516 19264
rect 3568 19292 3574 19304
rect 4080 19292 4108 19332
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 5350 19360 5356 19372
rect 5000 19332 5356 19360
rect 5000 19292 5028 19332
rect 5350 19320 5356 19332
rect 5408 19320 5414 19372
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8159 19332 8248 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 5166 19292 5172 19304
rect 3568 19264 4108 19292
rect 4356 19264 5028 19292
rect 5127 19264 5172 19292
rect 3568 19252 3574 19264
rect 2406 19224 2412 19236
rect 1596 19196 2412 19224
rect 1596 19165 1624 19196
rect 2406 19184 2412 19196
rect 2464 19184 2470 19236
rect 4356 19168 4384 19264
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5258 19252 5264 19304
rect 5316 19292 5322 19304
rect 5316 19264 5361 19292
rect 5316 19252 5322 19264
rect 5534 19252 5540 19304
rect 5592 19292 5598 19304
rect 5813 19295 5871 19301
rect 5813 19292 5825 19295
rect 5592 19264 5825 19292
rect 5592 19252 5598 19264
rect 5813 19261 5825 19264
rect 5859 19261 5871 19295
rect 6178 19292 6184 19304
rect 6139 19264 6184 19292
rect 5813 19255 5871 19261
rect 6178 19252 6184 19264
rect 6236 19252 6242 19304
rect 7377 19295 7435 19301
rect 7377 19261 7389 19295
rect 7423 19292 7435 19295
rect 7926 19292 7932 19304
rect 7423 19264 7932 19292
rect 7423 19261 7435 19264
rect 7377 19255 7435 19261
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8220 19292 8248 19332
rect 10042 19320 10048 19372
rect 10100 19360 10106 19372
rect 10778 19360 10784 19372
rect 10100 19332 10784 19360
rect 10100 19320 10106 19332
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19978 19360 19984 19372
rect 19484 19332 19984 19360
rect 19484 19320 19490 19332
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 20898 19360 20904 19372
rect 20772 19332 20904 19360
rect 20772 19320 20778 19332
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 8938 19292 8944 19304
rect 8220 19264 8616 19292
rect 8851 19264 8944 19292
rect 8588 19233 8616 19264
rect 8938 19252 8944 19264
rect 8996 19292 9002 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8996 19264 9045 19292
rect 8996 19252 9002 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12299 19264 12449 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12437 19261 12449 19264
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14148 19264 14933 19292
rect 14148 19252 14154 19264
rect 14921 19261 14933 19264
rect 14967 19292 14979 19295
rect 15381 19295 15439 19301
rect 15381 19292 15393 19295
rect 14967 19264 15393 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 15381 19261 15393 19264
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 8573 19227 8631 19233
rect 8573 19193 8585 19227
rect 8619 19224 8631 19227
rect 8619 19196 9168 19224
rect 8619 19193 8631 19196
rect 8573 19187 8631 19193
rect 1581 19159 1639 19165
rect 1581 19125 1593 19159
rect 1627 19125 1639 19159
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1581 19119 1639 19125
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 4338 19156 4344 19168
rect 4299 19128 4344 19156
rect 4338 19116 4344 19128
rect 4396 19116 4402 19168
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 6822 19156 6828 19168
rect 6687 19128 6828 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7466 19156 7472 19168
rect 7427 19128 7472 19156
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7616 19128 7849 19156
rect 7616 19116 7622 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 9140 19156 9168 19196
rect 9214 19184 9220 19236
rect 9272 19233 9278 19236
rect 9272 19227 9336 19233
rect 9272 19193 9290 19227
rect 9324 19193 9336 19227
rect 9272 19187 9336 19193
rect 9272 19184 9278 19187
rect 9858 19184 9864 19236
rect 9916 19224 9922 19236
rect 10226 19224 10232 19236
rect 9916 19196 10232 19224
rect 9916 19184 9922 19196
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 12710 19233 12716 19236
rect 12704 19224 12716 19233
rect 12671 19196 12716 19224
rect 12704 19187 12716 19196
rect 12710 19184 12716 19187
rect 12768 19184 12774 19236
rect 10413 19159 10471 19165
rect 10413 19156 10425 19159
rect 9140 19128 10425 19156
rect 7837 19119 7895 19125
rect 10413 19125 10425 19128
rect 10459 19156 10471 19159
rect 10778 19156 10784 19168
rect 10459 19128 10784 19156
rect 10459 19125 10471 19128
rect 10413 19119 10471 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11054 19156 11060 19168
rect 11015 19128 11060 19156
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 15102 19156 15108 19168
rect 15063 19128 15108 19156
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15896 19128 15945 19156
rect 15896 19116 15902 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1670 18952 1676 18964
rect 1631 18924 1676 18952
rect 1670 18912 1676 18924
rect 1728 18912 1734 18964
rect 2958 18912 2964 18964
rect 3016 18952 3022 18964
rect 3145 18955 3203 18961
rect 3145 18952 3157 18955
rect 3016 18924 3157 18952
rect 3016 18912 3022 18924
rect 3145 18921 3157 18924
rect 3191 18921 3203 18955
rect 3510 18952 3516 18964
rect 3471 18924 3516 18952
rect 3145 18915 3203 18921
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 5258 18952 5264 18964
rect 4755 18924 5264 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 7650 18952 7656 18964
rect 7611 18924 7656 18952
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 9125 18955 9183 18961
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 9214 18952 9220 18964
rect 9171 18924 9220 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 10413 18955 10471 18961
rect 10413 18921 10425 18955
rect 10459 18952 10471 18955
rect 11238 18952 11244 18964
rect 10459 18924 11244 18952
rect 10459 18921 10471 18924
rect 10413 18915 10471 18921
rect 11238 18912 11244 18924
rect 11296 18952 11302 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 11296 18924 13001 18952
rect 11296 18912 11302 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 12989 18915 13047 18921
rect 13354 18912 13360 18964
rect 13412 18952 13418 18964
rect 13449 18955 13507 18961
rect 13449 18952 13461 18955
rect 13412 18924 13461 18952
rect 13412 18912 13418 18924
rect 13449 18921 13461 18924
rect 13495 18921 13507 18955
rect 13449 18915 13507 18921
rect 5350 18844 5356 18896
rect 5408 18893 5414 18896
rect 5408 18887 5472 18893
rect 5408 18853 5426 18887
rect 5460 18853 5472 18887
rect 5408 18847 5472 18853
rect 5408 18844 5414 18847
rect 5534 18844 5540 18896
rect 5592 18844 5598 18896
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 9401 18887 9459 18893
rect 9401 18884 9413 18887
rect 7524 18856 9413 18884
rect 7524 18844 7530 18856
rect 9401 18853 9413 18856
rect 9447 18884 9459 18887
rect 9766 18884 9772 18896
rect 9447 18856 9772 18884
rect 9447 18853 9459 18856
rect 9401 18847 9459 18853
rect 9766 18844 9772 18856
rect 9824 18844 9830 18896
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 2133 18819 2191 18825
rect 2133 18816 2145 18819
rect 1452 18788 2145 18816
rect 1452 18776 1458 18788
rect 2133 18785 2145 18788
rect 2179 18785 2191 18819
rect 4062 18816 4068 18828
rect 4023 18788 4068 18816
rect 2133 18779 2191 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18816 5227 18819
rect 5552 18816 5580 18844
rect 5215 18788 5580 18816
rect 7193 18819 7251 18825
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 7650 18816 7656 18828
rect 7239 18788 7656 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 7650 18776 7656 18788
rect 7708 18816 7714 18828
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7708 18788 8033 18816
rect 7708 18776 7714 18788
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8110 18776 8116 18828
rect 8168 18816 8174 18828
rect 10778 18825 10784 18828
rect 10772 18816 10784 18825
rect 8168 18788 8213 18816
rect 10739 18788 10784 18816
rect 8168 18776 8174 18788
rect 10772 18779 10784 18788
rect 10778 18776 10784 18779
rect 10836 18776 10842 18828
rect 13354 18816 13360 18828
rect 13315 18788 13360 18816
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 2222 18748 2228 18760
rect 2183 18720 2228 18748
rect 2222 18708 2228 18720
rect 2280 18708 2286 18760
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 2958 18748 2964 18760
rect 2372 18720 2964 18748
rect 2372 18708 2378 18720
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 7558 18748 7564 18760
rect 7519 18720 7564 18748
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 9214 18748 9220 18760
rect 8343 18720 9220 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 9214 18708 9220 18720
rect 9272 18708 9278 18760
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18717 13599 18751
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 13541 18711 13599 18717
rect 1765 18615 1823 18621
rect 1765 18581 1777 18615
rect 1811 18612 1823 18615
rect 1946 18612 1952 18624
rect 1811 18584 1952 18612
rect 1811 18581 1823 18584
rect 1765 18575 1823 18581
rect 1946 18572 1952 18584
rect 2004 18612 2010 18624
rect 2682 18612 2688 18624
rect 2004 18584 2688 18612
rect 2004 18572 2010 18584
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 2866 18612 2872 18624
rect 2827 18584 2872 18612
rect 2866 18572 2872 18584
rect 2924 18572 2930 18624
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 5077 18615 5135 18621
rect 5077 18581 5089 18615
rect 5123 18612 5135 18615
rect 5166 18612 5172 18624
rect 5123 18584 5172 18612
rect 5123 18581 5135 18584
rect 5077 18575 5135 18581
rect 5166 18572 5172 18584
rect 5224 18572 5230 18624
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 6914 18612 6920 18624
rect 6595 18584 6920 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 9950 18612 9956 18624
rect 9911 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10520 18612 10548 18711
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 12710 18680 12716 18692
rect 12308 18652 12716 18680
rect 12308 18640 12314 18652
rect 12710 18640 12716 18652
rect 12768 18680 12774 18692
rect 12897 18683 12955 18689
rect 12897 18680 12909 18683
rect 12768 18652 12909 18680
rect 12768 18640 12774 18652
rect 12897 18649 12909 18652
rect 12943 18680 12955 18683
rect 13556 18680 13584 18711
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 16298 18748 16304 18760
rect 16259 18720 16304 18748
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 12943 18652 13584 18680
rect 12943 18649 12955 18652
rect 12897 18643 12955 18649
rect 10686 18612 10692 18624
rect 10520 18584 10692 18612
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 11790 18572 11796 18624
rect 11848 18612 11854 18624
rect 11885 18615 11943 18621
rect 11885 18612 11897 18615
rect 11848 18584 11897 18612
rect 11848 18572 11854 18584
rect 11885 18581 11897 18584
rect 11931 18581 11943 18615
rect 12526 18612 12532 18624
rect 12439 18584 12532 18612
rect 11885 18575 11943 18581
rect 12526 18572 12532 18584
rect 12584 18612 12590 18624
rect 13630 18612 13636 18624
rect 12584 18584 13636 18612
rect 12584 18572 12590 18584
rect 13630 18572 13636 18584
rect 13688 18612 13694 18624
rect 14001 18615 14059 18621
rect 14001 18612 14013 18615
rect 13688 18584 14013 18612
rect 13688 18572 13694 18584
rect 14001 18581 14013 18584
rect 14047 18581 14059 18615
rect 14001 18575 14059 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 2041 18411 2099 18417
rect 2041 18408 2053 18411
rect 1728 18380 2053 18408
rect 1728 18368 1734 18380
rect 2041 18377 2053 18380
rect 2087 18377 2099 18411
rect 2041 18371 2099 18377
rect 2056 18272 2084 18371
rect 2958 18368 2964 18420
rect 3016 18408 3022 18420
rect 3605 18411 3663 18417
rect 3605 18408 3617 18411
rect 3016 18380 3617 18408
rect 3016 18368 3022 18380
rect 3605 18377 3617 18380
rect 3651 18377 3663 18411
rect 3605 18371 3663 18377
rect 4249 18411 4307 18417
rect 4249 18377 4261 18411
rect 4295 18408 4307 18411
rect 4338 18408 4344 18420
rect 4295 18380 4344 18408
rect 4295 18377 4307 18380
rect 4249 18371 4307 18377
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 8202 18408 8208 18420
rect 8163 18380 8208 18408
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 9306 18408 9312 18420
rect 9267 18380 9312 18408
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 11425 18411 11483 18417
rect 11425 18408 11437 18411
rect 10836 18380 11437 18408
rect 10836 18368 10842 18380
rect 11425 18377 11437 18380
rect 11471 18377 11483 18411
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 11425 18371 11483 18377
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 13354 18408 13360 18420
rect 13315 18380 13360 18408
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 23845 18411 23903 18417
rect 23845 18377 23857 18411
rect 23891 18408 23903 18411
rect 24762 18408 24768 18420
rect 23891 18380 24768 18408
rect 23891 18377 23903 18380
rect 23845 18371 23903 18377
rect 24762 18368 24768 18380
rect 24820 18368 24826 18420
rect 8849 18343 8907 18349
rect 8849 18309 8861 18343
rect 8895 18340 8907 18343
rect 9214 18340 9220 18352
rect 8895 18312 9220 18340
rect 8895 18309 8907 18312
rect 8849 18303 8907 18309
rect 9214 18300 9220 18312
rect 9272 18300 9278 18352
rect 11882 18340 11888 18352
rect 9600 18312 11888 18340
rect 2225 18275 2283 18281
rect 2225 18272 2237 18275
rect 2056 18244 2237 18272
rect 2225 18241 2237 18244
rect 2271 18241 2283 18275
rect 5350 18272 5356 18284
rect 5311 18244 5356 18272
rect 2225 18235 2283 18241
rect 5350 18232 5356 18244
rect 5408 18272 5414 18284
rect 6086 18272 6092 18284
rect 5408 18244 6092 18272
rect 5408 18232 5414 18244
rect 6086 18232 6092 18244
rect 6144 18232 6150 18284
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18272 9183 18275
rect 9600 18272 9628 18312
rect 9766 18272 9772 18284
rect 9171 18244 9628 18272
rect 9727 18244 9772 18272
rect 9171 18241 9183 18244
rect 9125 18235 9183 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 9968 18281 9996 18312
rect 11882 18300 11888 18312
rect 11940 18300 11946 18352
rect 13081 18343 13139 18349
rect 13081 18309 13093 18343
rect 13127 18340 13139 18343
rect 13262 18340 13268 18352
rect 13127 18312 13268 18340
rect 13127 18309 13139 18312
rect 13081 18303 13139 18309
rect 13262 18300 13268 18312
rect 13320 18300 13326 18352
rect 14918 18340 14924 18352
rect 14879 18312 14924 18340
rect 14918 18300 14924 18312
rect 14976 18300 14982 18352
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 11054 18232 11060 18284
rect 11112 18272 11118 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 11112 18244 12449 18272
rect 11112 18232 11118 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 2492 18207 2550 18213
rect 2492 18173 2504 18207
rect 2538 18204 2550 18207
rect 2866 18204 2872 18216
rect 2538 18176 2872 18204
rect 2538 18173 2550 18176
rect 2492 18167 2550 18173
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 5074 18204 5080 18216
rect 4663 18176 5080 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 5592 18176 5825 18204
rect 5592 18164 5598 18176
rect 5813 18173 5825 18176
rect 5859 18204 5871 18207
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 5859 18176 6653 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 6641 18173 6653 18176
rect 6687 18204 6699 18207
rect 6822 18204 6828 18216
rect 6687 18176 6828 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 6822 18164 6828 18176
rect 6880 18204 6886 18216
rect 8938 18204 8944 18216
rect 6880 18176 8944 18204
rect 6880 18164 6886 18176
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 9674 18204 9680 18216
rect 9635 18176 9680 18204
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 10962 18204 10968 18216
rect 10919 18176 10968 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 10962 18164 10968 18176
rect 11020 18204 11026 18216
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 11020 18176 11805 18204
rect 11020 18164 11026 18176
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 13630 18204 13636 18216
rect 13587 18176 13636 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 16301 18207 16359 18213
rect 16301 18173 16313 18207
rect 16347 18204 16359 18207
rect 23658 18204 23664 18216
rect 16347 18176 16988 18204
rect 23619 18176 23664 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 4982 18096 4988 18148
rect 5040 18136 5046 18148
rect 5169 18139 5227 18145
rect 5169 18136 5181 18139
rect 5040 18108 5181 18136
rect 5040 18096 5046 18108
rect 5169 18105 5181 18108
rect 5215 18105 5227 18139
rect 5169 18099 5227 18105
rect 6914 18096 6920 18148
rect 6972 18136 6978 18148
rect 13814 18145 13820 18148
rect 7070 18139 7128 18145
rect 7070 18136 7082 18139
rect 6972 18108 7082 18136
rect 6972 18096 6978 18108
rect 7070 18105 7082 18108
rect 7116 18105 7128 18139
rect 13808 18136 13820 18145
rect 13775 18108 13820 18136
rect 7070 18099 7128 18105
rect 13808 18099 13820 18108
rect 13814 18096 13820 18099
rect 13872 18096 13878 18148
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 1673 18071 1731 18077
rect 1673 18068 1685 18071
rect 1452 18040 1685 18068
rect 1452 18028 1458 18040
rect 1673 18037 1685 18040
rect 1719 18037 1731 18071
rect 4706 18068 4712 18080
rect 4667 18040 4712 18068
rect 1673 18031 1731 18037
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 10597 18071 10655 18077
rect 10597 18037 10609 18071
rect 10643 18068 10655 18071
rect 10686 18068 10692 18080
rect 10643 18040 10692 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11054 18068 11060 18080
rect 11015 18040 11060 18068
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 16482 18068 16488 18080
rect 16443 18040 16488 18068
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 16960 18077 16988 18176
rect 23658 18164 23664 18176
rect 23716 18204 23722 18216
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 23716 18176 24133 18204
rect 23716 18164 23722 18176
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 24121 18167 24179 18173
rect 16945 18071 17003 18077
rect 16945 18037 16957 18071
rect 16991 18068 17003 18071
rect 17034 18068 17040 18080
rect 16991 18040 17040 18068
rect 16991 18037 17003 18040
rect 16945 18031 17003 18037
rect 17034 18028 17040 18040
rect 17092 18028 17098 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2222 17864 2228 17876
rect 2183 17836 2228 17864
rect 2222 17824 2228 17836
rect 2280 17864 2286 17876
rect 2317 17867 2375 17873
rect 2317 17864 2329 17867
rect 2280 17836 2329 17864
rect 2280 17824 2286 17836
rect 2317 17833 2329 17836
rect 2363 17833 2375 17867
rect 2317 17827 2375 17833
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 2832 17836 3341 17864
rect 2832 17824 2838 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 3329 17827 3387 17833
rect 3789 17867 3847 17873
rect 3789 17833 3801 17867
rect 3835 17864 3847 17867
rect 3878 17864 3884 17876
rect 3835 17836 3884 17864
rect 3835 17833 3847 17836
rect 3789 17827 3847 17833
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4249 17867 4307 17873
rect 4249 17864 4261 17867
rect 4120 17836 4261 17864
rect 4120 17824 4126 17836
rect 4249 17833 4261 17836
rect 4295 17833 4307 17867
rect 5534 17864 5540 17876
rect 4249 17827 4307 17833
rect 4724 17836 5540 17864
rect 2038 17756 2044 17808
rect 2096 17796 2102 17808
rect 4430 17796 4436 17808
rect 2096 17768 4436 17796
rect 2096 17756 2102 17768
rect 4430 17756 4436 17768
rect 4488 17756 4494 17808
rect 1857 17731 1915 17737
rect 1857 17697 1869 17731
rect 1903 17728 1915 17731
rect 2314 17728 2320 17740
rect 1903 17700 2320 17728
rect 1903 17697 1915 17700
rect 1857 17691 1915 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 2685 17731 2743 17737
rect 2685 17728 2697 17731
rect 2485 17700 2697 17728
rect 2222 17620 2228 17672
rect 2280 17660 2286 17672
rect 2485 17660 2513 17700
rect 2685 17697 2697 17700
rect 2731 17697 2743 17731
rect 2685 17691 2743 17697
rect 4614 17688 4620 17740
rect 4672 17728 4678 17740
rect 4724 17737 4752 17836
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 6086 17864 6092 17876
rect 6047 17836 6092 17864
rect 6086 17824 6092 17836
rect 6144 17824 6150 17876
rect 7650 17864 7656 17876
rect 7611 17836 7656 17864
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 9401 17867 9459 17873
rect 9401 17833 9413 17867
rect 9447 17864 9459 17867
rect 9582 17864 9588 17876
rect 9447 17836 9588 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 11977 17867 12035 17873
rect 11977 17833 11989 17867
rect 12023 17864 12035 17867
rect 12250 17864 12256 17876
rect 12023 17836 12256 17864
rect 12023 17833 12035 17836
rect 11977 17827 12035 17833
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 13446 17864 13452 17876
rect 13407 17836 13452 17864
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 17034 17864 17040 17876
rect 16995 17836 17040 17864
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 5166 17756 5172 17808
rect 5224 17756 5230 17808
rect 7561 17799 7619 17805
rect 7561 17765 7573 17799
rect 7607 17796 7619 17799
rect 8110 17796 8116 17808
rect 7607 17768 8116 17796
rect 7607 17765 7619 17768
rect 7561 17759 7619 17765
rect 8110 17756 8116 17768
rect 8168 17756 8174 17808
rect 8202 17756 8208 17808
rect 8260 17796 8266 17808
rect 8757 17799 8815 17805
rect 8757 17796 8769 17799
rect 8260 17768 8769 17796
rect 8260 17756 8266 17768
rect 8757 17765 8769 17768
rect 8803 17796 8815 17799
rect 9490 17796 9496 17808
rect 8803 17768 9496 17796
rect 8803 17765 8815 17768
rect 8757 17759 8815 17765
rect 9490 17756 9496 17768
rect 9548 17756 9554 17808
rect 10778 17756 10784 17808
rect 10836 17805 10842 17808
rect 10836 17799 10900 17805
rect 10836 17765 10854 17799
rect 10888 17765 10900 17799
rect 10836 17759 10900 17765
rect 10836 17756 10842 17759
rect 4709 17731 4767 17737
rect 4709 17728 4721 17731
rect 4672 17700 4721 17728
rect 4672 17688 4678 17700
rect 4709 17697 4721 17700
rect 4755 17697 4767 17731
rect 4709 17691 4767 17697
rect 4976 17731 5034 17737
rect 4976 17697 4988 17731
rect 5022 17728 5034 17731
rect 5184 17728 5212 17756
rect 5350 17728 5356 17740
rect 5022 17700 5356 17728
rect 5022 17697 5034 17700
rect 4976 17691 5034 17697
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 8018 17728 8024 17740
rect 7979 17700 8024 17728
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 10597 17731 10655 17737
rect 10597 17697 10609 17731
rect 10643 17728 10655 17731
rect 10686 17728 10692 17740
rect 10643 17700 10692 17728
rect 10643 17697 10655 17700
rect 10597 17691 10655 17697
rect 10686 17688 10692 17700
rect 10744 17728 10750 17740
rect 11146 17728 11152 17740
rect 10744 17700 11152 17728
rect 10744 17688 10750 17700
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17697 16911 17731
rect 17862 17728 17868 17740
rect 17823 17700 17868 17728
rect 16853 17691 16911 17697
rect 2280 17632 2513 17660
rect 2280 17620 2286 17632
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 2958 17660 2964 17672
rect 2832 17632 2877 17660
rect 2919 17632 2964 17660
rect 2832 17620 2838 17632
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 8110 17660 8116 17672
rect 8071 17632 8116 17660
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 8294 17660 8300 17672
rect 8255 17632 8300 17660
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 13538 17660 13544 17672
rect 13499 17632 13544 17660
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13722 17620 13728 17632
rect 13780 17660 13786 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13780 17632 14105 17660
rect 13780 17620 13786 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 15378 17620 15384 17672
rect 15436 17660 15442 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15436 17632 15761 17660
rect 15436 17620 15442 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 15896 17632 15941 17660
rect 15896 17620 15902 17632
rect 2038 17552 2044 17604
rect 2096 17592 2102 17604
rect 2976 17592 3004 17620
rect 13078 17592 13084 17604
rect 2096 17564 3004 17592
rect 13039 17564 13084 17592
rect 2096 17552 2102 17564
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 15289 17595 15347 17601
rect 15289 17561 15301 17595
rect 15335 17592 15347 17595
rect 16868 17592 16896 17691
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 17218 17592 17224 17604
rect 15335 17564 17224 17592
rect 15335 17561 15347 17564
rect 15289 17555 15347 17561
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 6914 17524 6920 17536
rect 6875 17496 6920 17524
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 9732 17496 9873 17524
rect 9732 17484 9738 17496
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 9861 17487 9919 17493
rect 12897 17527 12955 17533
rect 12897 17493 12909 17527
rect 12943 17524 12955 17527
rect 12986 17524 12992 17536
rect 12943 17496 12992 17524
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 18049 17527 18107 17533
rect 18049 17524 18061 17527
rect 18012 17496 18061 17524
rect 18012 17484 18018 17496
rect 18049 17493 18061 17496
rect 18095 17493 18107 17527
rect 18049 17487 18107 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 2038 17320 2044 17332
rect 1999 17292 2044 17320
rect 2038 17280 2044 17292
rect 2096 17280 2102 17332
rect 2222 17320 2228 17332
rect 2135 17292 2228 17320
rect 2222 17280 2228 17292
rect 2280 17320 2286 17332
rect 2317 17323 2375 17329
rect 2317 17320 2329 17323
rect 2280 17292 2329 17320
rect 2280 17280 2286 17292
rect 2317 17289 2329 17292
rect 2363 17289 2375 17323
rect 3510 17320 3516 17332
rect 3471 17292 3516 17320
rect 2317 17283 2375 17289
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4249 17323 4307 17329
rect 4249 17320 4261 17323
rect 4212 17292 4261 17320
rect 4212 17280 4218 17292
rect 4249 17289 4261 17292
rect 4295 17289 4307 17323
rect 4249 17283 4307 17289
rect 5353 17323 5411 17329
rect 5353 17289 5365 17323
rect 5399 17320 5411 17323
rect 5534 17320 5540 17332
rect 5399 17292 5540 17320
rect 5399 17289 5411 17292
rect 5353 17283 5411 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 7558 17320 7564 17332
rect 7519 17292 7564 17320
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 8128 17292 10517 17320
rect 2498 17212 2504 17264
rect 2556 17252 2562 17264
rect 2685 17255 2743 17261
rect 2685 17252 2697 17255
rect 2556 17224 2697 17252
rect 2556 17212 2562 17224
rect 2685 17221 2697 17224
rect 2731 17221 2743 17255
rect 2685 17215 2743 17221
rect 2774 17212 2780 17264
rect 2832 17252 2838 17264
rect 3145 17255 3203 17261
rect 3145 17252 3157 17255
rect 2832 17224 3157 17252
rect 2832 17212 2838 17224
rect 3145 17221 3157 17224
rect 3191 17252 3203 17255
rect 5442 17252 5448 17264
rect 3191 17224 5448 17252
rect 3191 17221 3203 17224
rect 3145 17215 3203 17221
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 3878 17184 3884 17196
rect 1412 17156 3884 17184
rect 1412 17125 1440 17156
rect 3878 17144 3884 17156
rect 3936 17144 3942 17196
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4203 17156 4813 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 4801 17153 4813 17156
rect 4847 17184 4859 17187
rect 6914 17184 6920 17196
rect 4847 17156 6920 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 8128 17193 8156 17292
rect 10505 17289 10517 17292
rect 10551 17320 10563 17323
rect 10778 17320 10784 17332
rect 10551 17292 10784 17320
rect 10551 17289 10563 17292
rect 10505 17283 10563 17289
rect 10778 17280 10784 17292
rect 10836 17320 10842 17332
rect 11425 17323 11483 17329
rect 11425 17320 11437 17323
rect 10836 17292 11437 17320
rect 10836 17280 10842 17292
rect 11425 17289 11437 17292
rect 11471 17289 11483 17323
rect 11425 17283 11483 17289
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 13722 17320 13728 17332
rect 12299 17292 13728 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 13722 17280 13728 17292
rect 13780 17320 13786 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 13780 17292 14197 17320
rect 13780 17280 13786 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 14829 17323 14887 17329
rect 14829 17289 14841 17323
rect 14875 17320 14887 17323
rect 15654 17320 15660 17332
rect 14875 17292 15660 17320
rect 14875 17289 14887 17292
rect 14829 17283 14887 17289
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 17218 17320 17224 17332
rect 17179 17292 17224 17320
rect 17218 17280 17224 17292
rect 17276 17280 17282 17332
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 18509 17323 18567 17329
rect 18509 17320 18521 17323
rect 17920 17292 18521 17320
rect 17920 17280 17926 17292
rect 18509 17289 18521 17292
rect 18555 17289 18567 17323
rect 18509 17283 18567 17289
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 8573 17255 8631 17261
rect 8573 17252 8585 17255
rect 8352 17224 8585 17252
rect 8352 17212 8358 17224
rect 8573 17221 8585 17224
rect 8619 17221 8631 17255
rect 8938 17252 8944 17264
rect 8899 17224 8944 17252
rect 8573 17215 8631 17221
rect 8938 17212 8944 17224
rect 8996 17252 9002 17264
rect 8996 17224 9168 17252
rect 8996 17212 9002 17224
rect 9140 17193 9168 17224
rect 19334 17212 19340 17264
rect 19392 17252 19398 17264
rect 20254 17252 20260 17264
rect 19392 17224 20260 17252
rect 19392 17212 19398 17224
rect 20254 17212 20260 17224
rect 20312 17212 20318 17264
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17184 7159 17187
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 7147 17156 8125 17184
rect 7147 17153 7159 17156
rect 7101 17147 7159 17153
rect 8113 17153 8125 17156
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17153 9183 17187
rect 18046 17184 18052 17196
rect 18007 17156 18052 17184
rect 9125 17147 9183 17153
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 3510 17116 3516 17128
rect 2547 17088 3516 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17116 4675 17119
rect 4706 17116 4712 17128
rect 4663 17088 4712 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 7926 17116 7932 17128
rect 7887 17088 7932 17116
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17116 8079 17119
rect 8202 17116 8208 17128
rect 8067 17088 8208 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 9398 17125 9404 17128
rect 9392 17116 9404 17125
rect 9359 17088 9404 17116
rect 9392 17079 9404 17088
rect 9398 17076 9404 17079
rect 9456 17076 9462 17128
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17085 12863 17119
rect 12805 17079 12863 17085
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 15556 17119 15614 17125
rect 15335 17088 15424 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 4982 17008 4988 17060
rect 5040 17048 5046 17060
rect 5997 17051 6055 17057
rect 5997 17048 6009 17051
rect 5040 17020 6009 17048
rect 5040 17008 5046 17020
rect 5997 17017 6009 17020
rect 6043 17017 6055 17051
rect 5997 17011 6055 17017
rect 2225 16983 2283 16989
rect 2225 16949 2237 16983
rect 2271 16980 2283 16983
rect 3050 16980 3056 16992
rect 2271 16952 3056 16980
rect 2271 16949 2283 16952
rect 2225 16943 2283 16949
rect 3050 16940 3056 16952
rect 3108 16940 3114 16992
rect 4709 16983 4767 16989
rect 4709 16949 4721 16983
rect 4755 16980 4767 16983
rect 4798 16980 4804 16992
rect 4755 16952 4804 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 5629 16983 5687 16989
rect 5629 16980 5641 16983
rect 5408 16952 5641 16980
rect 5408 16940 5414 16952
rect 5629 16949 5641 16952
rect 5675 16949 5687 16983
rect 6546 16980 6552 16992
rect 6507 16952 6552 16980
rect 5629 16943 5687 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 11146 16980 11152 16992
rect 11059 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16980 11210 16992
rect 12713 16983 12771 16989
rect 12713 16980 12725 16983
rect 11204 16952 12725 16980
rect 11204 16940 11210 16952
rect 12713 16949 12725 16952
rect 12759 16980 12771 16983
rect 12820 16980 12848 17079
rect 13078 17057 13084 17060
rect 13072 17048 13084 17057
rect 13039 17020 13084 17048
rect 13072 17011 13084 17020
rect 13078 17008 13084 17011
rect 13136 17008 13142 17060
rect 13630 16980 13636 16992
rect 12759 16952 13636 16980
rect 12759 16949 12771 16952
rect 12713 16943 12771 16949
rect 13630 16940 13636 16952
rect 13688 16980 13694 16992
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 13688 16952 15209 16980
rect 13688 16940 13694 16952
rect 15197 16949 15209 16952
rect 15243 16980 15255 16983
rect 15396 16980 15424 17088
rect 15556 17085 15568 17119
rect 15602 17116 15614 17119
rect 15838 17116 15844 17128
rect 15602 17088 15844 17116
rect 15602 17085 15614 17088
rect 15556 17079 15614 17085
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 16206 16980 16212 16992
rect 15243 16952 16212 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 16669 16983 16727 16989
rect 16669 16980 16681 16983
rect 16632 16952 16681 16980
rect 16632 16940 16638 16952
rect 16669 16949 16681 16952
rect 16715 16949 16727 16983
rect 16669 16943 16727 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1394 16776 1400 16788
rect 1355 16748 1400 16776
rect 1394 16736 1400 16748
rect 1452 16736 1458 16788
rect 2317 16779 2375 16785
rect 2317 16745 2329 16779
rect 2363 16776 2375 16779
rect 2682 16776 2688 16788
rect 2363 16748 2688 16776
rect 2363 16745 2375 16748
rect 2317 16739 2375 16745
rect 2682 16736 2688 16748
rect 2740 16776 2746 16788
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2740 16748 2881 16776
rect 2740 16736 2746 16748
rect 2869 16745 2881 16748
rect 2915 16745 2927 16779
rect 2869 16739 2927 16745
rect 3881 16779 3939 16785
rect 3881 16745 3893 16779
rect 3927 16776 3939 16779
rect 4706 16776 4712 16788
rect 3927 16748 4712 16776
rect 3927 16745 3939 16748
rect 3881 16739 3939 16745
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 5169 16779 5227 16785
rect 5169 16745 5181 16779
rect 5215 16776 5227 16779
rect 5442 16776 5448 16788
rect 5215 16748 5448 16776
rect 5215 16745 5227 16748
rect 5169 16739 5227 16745
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 7984 16748 8033 16776
rect 7984 16736 7990 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 9217 16779 9275 16785
rect 9217 16745 9229 16779
rect 9263 16776 9275 16779
rect 9398 16776 9404 16788
rect 9263 16748 9404 16776
rect 9263 16745 9275 16748
rect 9217 16739 9275 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9732 16748 9873 16776
rect 9732 16736 9738 16748
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 11422 16776 11428 16788
rect 11383 16748 11428 16776
rect 9861 16739 9919 16745
rect 11422 16736 11428 16748
rect 11480 16736 11486 16788
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16776 12035 16779
rect 13538 16776 13544 16788
rect 12023 16748 13544 16776
rect 12023 16745 12035 16748
rect 11977 16739 12035 16745
rect 13538 16736 13544 16748
rect 13596 16776 13602 16788
rect 13817 16779 13875 16785
rect 13817 16776 13829 16779
rect 13596 16748 13829 16776
rect 13596 16736 13602 16748
rect 13817 16745 13829 16748
rect 13863 16745 13875 16779
rect 14274 16776 14280 16788
rect 14235 16748 14280 16776
rect 13817 16739 13875 16745
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 15470 16776 15476 16788
rect 15431 16748 15476 16776
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 15838 16776 15844 16788
rect 15799 16748 15844 16776
rect 15838 16736 15844 16748
rect 15896 16776 15902 16788
rect 16117 16779 16175 16785
rect 16117 16776 16129 16779
rect 15896 16748 16129 16776
rect 15896 16736 15902 16748
rect 16117 16745 16129 16748
rect 16163 16745 16175 16779
rect 16117 16739 16175 16745
rect 19337 16779 19395 16785
rect 19337 16745 19349 16779
rect 19383 16776 19395 16779
rect 19426 16776 19432 16788
rect 19383 16748 19432 16776
rect 19383 16745 19395 16748
rect 19337 16739 19395 16745
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 4341 16711 4399 16717
rect 4341 16677 4353 16711
rect 4387 16708 4399 16711
rect 4798 16708 4804 16720
rect 4387 16680 4804 16708
rect 4387 16677 4399 16680
rect 4341 16671 4399 16677
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 4890 16668 4896 16720
rect 4948 16708 4954 16720
rect 7006 16708 7012 16720
rect 4948 16680 7012 16708
rect 4948 16668 4954 16680
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 7374 16668 7380 16720
rect 7432 16708 7438 16720
rect 8110 16708 8116 16720
rect 7432 16680 8116 16708
rect 7432 16668 7438 16680
rect 8110 16668 8116 16680
rect 8168 16708 8174 16720
rect 8481 16711 8539 16717
rect 8481 16708 8493 16711
rect 8168 16680 8493 16708
rect 8168 16668 8174 16680
rect 8481 16677 8493 16680
rect 8527 16677 8539 16711
rect 8481 16671 8539 16677
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 4982 16640 4988 16652
rect 2832 16612 2877 16640
rect 4724 16612 4988 16640
rect 2832 16600 2838 16612
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3099 16544 3556 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 1949 16439 2007 16445
rect 1949 16405 1961 16439
rect 1995 16436 2007 16439
rect 2222 16436 2228 16448
rect 1995 16408 2228 16436
rect 1995 16405 2007 16408
rect 1949 16399 2007 16405
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 2406 16436 2412 16448
rect 2367 16408 2412 16436
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 3528 16445 3556 16544
rect 4724 16513 4752 16612
rect 4982 16600 4988 16612
rect 5040 16600 5046 16652
rect 5074 16600 5080 16652
rect 5132 16640 5138 16652
rect 6362 16640 6368 16652
rect 5132 16612 5177 16640
rect 6323 16612 6368 16640
rect 5132 16600 5138 16612
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 6822 16640 6828 16652
rect 6783 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16640 7803 16643
rect 8018 16640 8024 16652
rect 7791 16612 8024 16640
rect 7791 16609 7803 16612
rect 7745 16603 7803 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8386 16640 8392 16652
rect 8347 16612 8392 16640
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 5350 16572 5356 16584
rect 5311 16544 5356 16572
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 6914 16572 6920 16584
rect 6875 16544 6920 16572
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 8665 16575 8723 16581
rect 8665 16541 8677 16575
rect 8711 16572 8723 16575
rect 9398 16572 9404 16584
rect 8711 16544 9404 16572
rect 8711 16541 8723 16544
rect 8665 16535 8723 16541
rect 4709 16507 4767 16513
rect 4709 16473 4721 16507
rect 4755 16473 4767 16507
rect 4709 16467 4767 16473
rect 6546 16464 6552 16516
rect 6604 16504 6610 16516
rect 7024 16504 7052 16535
rect 9398 16532 9404 16544
rect 9456 16532 9462 16584
rect 9692 16572 9720 16603
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 9824 16612 10609 16640
rect 9824 16600 9830 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10781 16643 10839 16649
rect 10781 16609 10793 16643
rect 10827 16640 10839 16643
rect 11440 16640 11468 16736
rect 13446 16708 13452 16720
rect 13407 16680 13452 16708
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 13722 16668 13728 16720
rect 13780 16708 13786 16720
rect 15105 16711 15163 16717
rect 15105 16708 15117 16711
rect 13780 16680 15117 16708
rect 13780 16668 13786 16680
rect 15105 16677 15117 16680
rect 15151 16708 15163 16711
rect 15378 16708 15384 16720
rect 15151 16680 15384 16708
rect 15151 16677 15163 16680
rect 15105 16671 15163 16677
rect 15378 16668 15384 16680
rect 15436 16668 15442 16720
rect 16850 16668 16856 16720
rect 16908 16717 16914 16720
rect 16908 16711 16972 16717
rect 16908 16677 16926 16711
rect 16960 16677 16972 16711
rect 16908 16671 16972 16677
rect 16908 16668 16914 16671
rect 10827 16612 11468 16640
rect 10827 16609 10839 16612
rect 10781 16603 10839 16609
rect 12250 16600 12256 16652
rect 12308 16640 12314 16652
rect 12345 16643 12403 16649
rect 12345 16640 12357 16643
rect 12308 16612 12357 16640
rect 12308 16600 12314 16612
rect 12345 16609 12357 16612
rect 12391 16609 12403 16643
rect 13078 16640 13084 16652
rect 12345 16603 12403 16609
rect 12636 16612 13084 16640
rect 10686 16572 10692 16584
rect 9692 16544 10692 16572
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12636 16581 12664 16612
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16640 14151 16643
rect 14182 16640 14188 16652
rect 14139 16612 14188 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14642 16600 14648 16652
rect 14700 16640 14706 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 14700 16612 15301 16640
rect 14700 16600 14706 16612
rect 15289 16609 15301 16612
rect 15335 16640 15347 16643
rect 16114 16640 16120 16652
rect 15335 16612 16120 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 19150 16640 19156 16652
rect 19111 16612 19156 16640
rect 19150 16600 19156 16612
rect 19208 16640 19214 16652
rect 19208 16612 19288 16640
rect 19208 16600 19214 16612
rect 12621 16575 12679 16581
rect 12492 16544 12537 16572
rect 12492 16532 12498 16544
rect 12621 16541 12633 16575
rect 12667 16541 12679 16575
rect 12621 16535 12679 16541
rect 6604 16476 7052 16504
rect 6604 16464 6610 16476
rect 12342 16464 12348 16516
rect 12400 16504 12406 16516
rect 12636 16504 12664 16535
rect 16206 16532 16212 16584
rect 16264 16572 16270 16584
rect 16669 16575 16727 16581
rect 16669 16572 16681 16575
rect 16264 16544 16681 16572
rect 16264 16532 16270 16544
rect 16669 16541 16681 16544
rect 16715 16541 16727 16575
rect 19260 16572 19288 16612
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22462 16640 22468 16652
rect 22152 16612 22468 16640
rect 22152 16600 22158 16612
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 19886 16572 19892 16584
rect 19260 16544 19892 16572
rect 16669 16535 16727 16541
rect 19886 16532 19892 16544
rect 19944 16532 19950 16584
rect 12400 16476 12664 16504
rect 12400 16464 12406 16476
rect 3513 16439 3571 16445
rect 3513 16405 3525 16439
rect 3559 16436 3571 16439
rect 3878 16436 3884 16448
rect 3559 16408 3884 16436
rect 3559 16405 3571 16408
rect 3513 16399 3571 16405
rect 3878 16396 3884 16408
rect 3936 16396 3942 16448
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 5721 16439 5779 16445
rect 5721 16436 5733 16439
rect 5316 16408 5733 16436
rect 5316 16396 5322 16408
rect 5721 16405 5733 16408
rect 5767 16405 5779 16439
rect 6454 16436 6460 16448
rect 6415 16408 6460 16436
rect 5721 16399 5779 16405
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 9950 16396 9956 16448
rect 10008 16436 10014 16448
rect 10229 16439 10287 16445
rect 10229 16436 10241 16439
rect 10008 16408 10241 16436
rect 10008 16396 10014 16408
rect 10229 16405 10241 16408
rect 10275 16405 10287 16439
rect 10962 16436 10968 16448
rect 10923 16408 10968 16436
rect 10229 16399 10287 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 13170 16436 13176 16448
rect 13131 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 15378 16436 15384 16448
rect 14792 16408 15384 16436
rect 14792 16396 14798 16408
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 18046 16436 18052 16448
rect 18007 16408 18052 16436
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 3142 16192 3148 16244
rect 3200 16232 3206 16244
rect 4709 16235 4767 16241
rect 4709 16232 4721 16235
rect 3200 16204 4721 16232
rect 3200 16192 3206 16204
rect 4709 16201 4721 16204
rect 4755 16232 4767 16235
rect 5074 16232 5080 16244
rect 4755 16204 5080 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5408 16204 6193 16232
rect 5408 16192 5414 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 6270 16192 6276 16244
rect 6328 16232 6334 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6328 16204 6561 16232
rect 6328 16192 6334 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 6549 16195 6607 16201
rect 4433 16167 4491 16173
rect 4433 16133 4445 16167
rect 4479 16164 4491 16167
rect 5442 16164 5448 16176
rect 4479 16136 5448 16164
rect 4479 16133 4491 16136
rect 4433 16127 4491 16133
rect 5442 16124 5448 16136
rect 5500 16124 5506 16176
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16096 2286 16108
rect 2866 16096 2872 16108
rect 2280 16068 2872 16096
rect 2280 16056 2286 16068
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 3878 16096 3884 16108
rect 3839 16068 3884 16096
rect 3878 16056 3884 16068
rect 3936 16056 3942 16108
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5316 16068 5733 16096
rect 5316 16056 5322 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 6564 16096 6592 16195
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7432 16204 8033 16232
rect 7432 16192 7438 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9398 16232 9404 16244
rect 9079 16204 9404 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 11606 16232 11612 16244
rect 11567 16204 11612 16232
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 13081 16235 13139 16241
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13722 16232 13728 16244
rect 13127 16204 13728 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 16025 16235 16083 16241
rect 16025 16232 16037 16235
rect 15896 16204 16037 16232
rect 15896 16192 15902 16204
rect 16025 16201 16037 16204
rect 16071 16201 16083 16235
rect 19886 16232 19892 16244
rect 19847 16204 19892 16232
rect 16025 16195 16083 16201
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 20622 16232 20628 16244
rect 20583 16204 20628 16232
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 6822 16124 6828 16176
rect 6880 16164 6886 16176
rect 6917 16167 6975 16173
rect 6917 16164 6929 16167
rect 6880 16136 6929 16164
rect 6880 16124 6886 16136
rect 6917 16133 6929 16136
rect 6963 16164 6975 16167
rect 8938 16164 8944 16176
rect 6963 16136 8944 16164
rect 6963 16133 6975 16136
rect 6917 16127 6975 16133
rect 8938 16124 8944 16136
rect 8996 16124 9002 16176
rect 7374 16096 7380 16108
rect 6564 16068 7380 16096
rect 5721 16059 5779 16065
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16096 7619 16099
rect 7834 16096 7840 16108
rect 7607 16068 7840 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 8481 16099 8539 16105
rect 8481 16096 8493 16099
rect 8444 16068 8493 16096
rect 8444 16056 8450 16068
rect 8481 16065 8493 16068
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 10042 16096 10048 16108
rect 9447 16068 10048 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13228 16068 13553 16096
rect 13228 16056 13234 16068
rect 13541 16065 13553 16068
rect 13587 16096 13599 16099
rect 13630 16096 13636 16108
rect 13587 16068 13636 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 13771 16068 14228 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 2038 16028 2044 16040
rect 1999 16000 2044 16028
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 3602 16028 3608 16040
rect 3563 16000 3608 16028
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 4614 15988 4620 16040
rect 4672 16028 4678 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 4672 16000 5641 16028
rect 4672 15988 4678 16000
rect 5629 15997 5641 16000
rect 5675 16028 5687 16031
rect 6454 16028 6460 16040
rect 5675 16000 6460 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 10980 16000 11069 16028
rect 2130 15960 2136 15972
rect 2091 15932 2136 15960
rect 2130 15920 2136 15932
rect 2188 15920 2194 15972
rect 2682 15920 2688 15972
rect 2740 15960 2746 15972
rect 3145 15963 3203 15969
rect 3145 15960 3157 15963
rect 2740 15932 3157 15960
rect 2740 15920 2746 15932
rect 3145 15929 3157 15932
rect 3191 15960 3203 15963
rect 3191 15932 3740 15960
rect 3191 15929 3203 15932
rect 3145 15923 3203 15929
rect 3712 15904 3740 15932
rect 9214 15920 9220 15972
rect 9272 15960 9278 15972
rect 9861 15963 9919 15969
rect 9861 15960 9873 15963
rect 9272 15932 9873 15960
rect 9272 15920 9278 15932
rect 9861 15929 9873 15932
rect 9907 15929 9919 15963
rect 9861 15923 9919 15929
rect 10980 15904 11008 16000
rect 11057 15997 11069 16000
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 11606 15920 11612 15972
rect 11664 15960 11670 15972
rect 12434 15960 12440 15972
rect 11664 15932 12440 15960
rect 11664 15920 11670 15932
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 14200 15969 14228 16068
rect 14642 16028 14648 16040
rect 14603 16000 14648 16028
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 14918 16037 14924 16040
rect 14912 16028 14924 16037
rect 14844 16000 14924 16028
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 12912 15932 13461 15960
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2774 15852 2780 15904
rect 2832 15892 2838 15904
rect 3237 15895 3295 15901
rect 2832 15864 2877 15892
rect 2832 15852 2838 15864
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 3326 15892 3332 15904
rect 3283 15864 3332 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 3694 15892 3700 15904
rect 3655 15864 3700 15892
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5537 15895 5595 15901
rect 5537 15861 5549 15895
rect 5583 15892 5595 15895
rect 5994 15892 6000 15904
rect 5583 15864 6000 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 7285 15895 7343 15901
rect 7285 15892 7297 15895
rect 7064 15864 7297 15892
rect 7064 15852 7070 15864
rect 7285 15861 7297 15864
rect 7331 15861 7343 15895
rect 9490 15892 9496 15904
rect 9451 15864 9496 15892
rect 7285 15855 7343 15861
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 10597 15895 10655 15901
rect 10008 15864 10053 15892
rect 10008 15852 10014 15864
rect 10597 15861 10609 15895
rect 10643 15892 10655 15895
rect 10686 15892 10692 15904
rect 10643 15864 10692 15892
rect 10643 15861 10655 15864
rect 10597 15855 10655 15861
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 10962 15892 10968 15904
rect 10923 15864 10968 15892
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11238 15892 11244 15904
rect 11199 15864 11244 15892
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 12069 15895 12127 15901
rect 12069 15861 12081 15895
rect 12115 15892 12127 15895
rect 12250 15892 12256 15904
rect 12115 15864 12256 15892
rect 12115 15861 12127 15864
rect 12069 15855 12127 15861
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 12912 15901 12940 15932
rect 13449 15929 13461 15932
rect 13495 15929 13507 15963
rect 13449 15923 13507 15929
rect 14185 15963 14243 15969
rect 14185 15929 14197 15963
rect 14231 15960 14243 15963
rect 14844 15960 14872 16000
rect 14912 15991 14924 16000
rect 14918 15988 14924 15991
rect 14976 15988 14982 16040
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 18046 15988 18052 16000
rect 18104 16028 18110 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18104 16000 18521 16028
rect 18104 15988 18110 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 19058 16028 19064 16040
rect 19019 16000 19064 16028
rect 18509 15991 18567 15997
rect 19058 15988 19064 16000
rect 19116 16028 19122 16040
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 19116 16000 19533 16028
rect 19116 15988 19122 16000
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 20438 16028 20444 16040
rect 20399 16000 20444 16028
rect 19521 15991 19579 15997
rect 20438 15988 20444 16000
rect 20496 16028 20502 16040
rect 20993 16031 21051 16037
rect 20993 16028 21005 16031
rect 20496 16000 21005 16028
rect 20496 15988 20502 16000
rect 20993 15997 21005 16000
rect 21039 15997 21051 16031
rect 20993 15991 21051 15997
rect 14231 15932 14872 15960
rect 14231 15929 14243 15932
rect 14185 15923 14243 15929
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12676 15864 12909 15892
rect 12676 15852 12682 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 14553 15895 14611 15901
rect 14553 15861 14565 15895
rect 14599 15892 14611 15895
rect 14642 15892 14648 15904
rect 14599 15864 14648 15892
rect 14599 15861 14611 15864
rect 14553 15855 14611 15861
rect 14642 15852 14648 15864
rect 14700 15892 14706 15904
rect 16206 15892 16212 15904
rect 14700 15864 16212 15892
rect 14700 15852 14706 15864
rect 16206 15852 16212 15864
rect 16264 15892 16270 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16264 15864 16681 15892
rect 16264 15852 16270 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17037 15895 17095 15901
rect 17037 15892 17049 15895
rect 16908 15864 17049 15892
rect 16908 15852 16914 15864
rect 17037 15861 17049 15864
rect 17083 15861 17095 15895
rect 18230 15892 18236 15904
rect 18191 15864 18236 15892
rect 17037 15855 17095 15861
rect 18230 15852 18236 15864
rect 18288 15852 18294 15904
rect 19242 15892 19248 15904
rect 19203 15864 19248 15892
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2866 15688 2872 15700
rect 2827 15660 2872 15688
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 3513 15691 3571 15697
rect 3513 15657 3525 15691
rect 3559 15688 3571 15691
rect 3602 15688 3608 15700
rect 3559 15660 3608 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 3602 15648 3608 15660
rect 3660 15648 3666 15700
rect 4614 15688 4620 15700
rect 4575 15660 4620 15688
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 6972 15660 7205 15688
rect 6972 15648 6978 15660
rect 7193 15657 7205 15660
rect 7239 15657 7251 15691
rect 7193 15651 7251 15657
rect 8297 15691 8355 15697
rect 8297 15657 8309 15691
rect 8343 15688 8355 15691
rect 8386 15688 8392 15700
rect 8343 15660 8392 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 4154 15580 4160 15632
rect 4212 15620 4218 15632
rect 4522 15620 4528 15632
rect 4212 15592 4528 15620
rect 4212 15580 4218 15592
rect 4522 15580 4528 15592
rect 4580 15620 4586 15632
rect 7006 15620 7012 15632
rect 4580 15592 7012 15620
rect 4580 15580 4586 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 7208 15620 7236 15651
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 8938 15688 8944 15700
rect 8899 15660 8944 15688
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 12342 15688 12348 15700
rect 12303 15660 12348 15688
rect 12342 15648 12348 15660
rect 12400 15648 12406 15700
rect 14182 15688 14188 15700
rect 14143 15660 14188 15688
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 14918 15688 14924 15700
rect 14783 15660 14924 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15473 15691 15531 15697
rect 15473 15657 15485 15691
rect 15519 15688 15531 15691
rect 15562 15688 15568 15700
rect 15519 15660 15568 15688
rect 15519 15657 15531 15660
rect 15473 15651 15531 15657
rect 15562 15648 15568 15660
rect 15620 15648 15626 15700
rect 16114 15688 16120 15700
rect 16075 15660 16120 15688
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 16850 15648 16856 15700
rect 16908 15688 16914 15700
rect 17773 15691 17831 15697
rect 17773 15688 17785 15691
rect 16908 15660 17785 15688
rect 16908 15648 16914 15660
rect 17773 15657 17785 15660
rect 17819 15657 17831 15691
rect 17773 15651 17831 15657
rect 8573 15623 8631 15629
rect 8573 15620 8585 15623
rect 7208 15592 8585 15620
rect 8573 15589 8585 15592
rect 8619 15589 8631 15623
rect 8573 15583 8631 15589
rect 10042 15580 10048 15632
rect 10100 15620 10106 15632
rect 10566 15623 10624 15629
rect 10566 15620 10578 15623
rect 10100 15592 10578 15620
rect 10100 15580 10106 15592
rect 10566 15589 10578 15592
rect 10612 15620 10624 15623
rect 10870 15620 10876 15632
rect 10612 15592 10876 15620
rect 10612 15589 10624 15592
rect 10566 15583 10624 15589
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 13173 15623 13231 15629
rect 13173 15589 13185 15623
rect 13219 15620 13231 15623
rect 13354 15620 13360 15632
rect 13219 15592 13360 15620
rect 13219 15589 13231 15592
rect 13173 15583 13231 15589
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 1762 15561 1768 15564
rect 1756 15515 1768 15561
rect 1820 15552 1826 15564
rect 4706 15552 4712 15564
rect 1820 15524 1856 15552
rect 4667 15524 4712 15552
rect 1762 15512 1768 15515
rect 1820 15512 1826 15524
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 4976 15555 5034 15561
rect 4976 15521 4988 15555
rect 5022 15552 5034 15555
rect 5258 15552 5264 15564
rect 5022 15524 5264 15552
rect 5022 15521 5034 15524
rect 4976 15515 5034 15521
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 7558 15552 7564 15564
rect 7519 15524 7564 15552
rect 7558 15512 7564 15524
rect 7616 15552 7622 15564
rect 8294 15552 8300 15564
rect 7616 15524 8300 15552
rect 7616 15512 7622 15524
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15552 15350 15564
rect 15749 15555 15807 15561
rect 15749 15552 15761 15555
rect 15344 15524 15761 15552
rect 15344 15512 15350 15524
rect 15749 15521 15761 15524
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 16660 15555 16718 15561
rect 16660 15521 16672 15555
rect 16706 15552 16718 15555
rect 17402 15552 17408 15564
rect 16706 15524 17408 15552
rect 16706 15521 16718 15524
rect 16660 15515 16718 15521
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 1489 15487 1547 15493
rect 1489 15453 1501 15487
rect 1535 15453 1547 15487
rect 1489 15447 1547 15453
rect 1504 15348 1532 15447
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7653 15487 7711 15493
rect 7653 15484 7665 15487
rect 7340 15456 7665 15484
rect 7340 15444 7346 15456
rect 7653 15453 7665 15456
rect 7699 15453 7711 15487
rect 7834 15484 7840 15496
rect 7795 15456 7840 15484
rect 7653 15447 7711 15453
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 13265 15487 13323 15493
rect 13265 15484 13277 15487
rect 12492 15456 13277 15484
rect 12492 15444 12498 15456
rect 13265 15453 13277 15456
rect 13311 15453 13323 15487
rect 13265 15447 13323 15453
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 12802 15416 12808 15428
rect 12763 15388 12808 15416
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 13170 15376 13176 15428
rect 13228 15416 13234 15428
rect 13372 15416 13400 15447
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 16393 15487 16451 15493
rect 16393 15484 16405 15487
rect 16264 15456 16405 15484
rect 16264 15444 16270 15456
rect 16393 15453 16405 15456
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 13228 15388 13400 15416
rect 13228 15376 13234 15388
rect 1670 15348 1676 15360
rect 1504 15320 1676 15348
rect 1670 15308 1676 15320
rect 1728 15308 1734 15360
rect 3878 15348 3884 15360
rect 3791 15320 3884 15348
rect 3878 15308 3884 15320
rect 3936 15348 3942 15360
rect 4614 15348 4620 15360
rect 3936 15320 4620 15348
rect 3936 15308 3942 15320
rect 4614 15308 4620 15320
rect 4672 15348 4678 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 4672 15320 6101 15348
rect 4672 15308 4678 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 9214 15308 9220 15360
rect 9272 15348 9278 15360
rect 9401 15351 9459 15357
rect 9401 15348 9413 15351
rect 9272 15320 9413 15348
rect 9272 15308 9278 15320
rect 9401 15317 9413 15320
rect 9447 15317 9459 15351
rect 9401 15311 9459 15317
rect 9953 15351 10011 15357
rect 9953 15317 9965 15351
rect 9999 15348 10011 15351
rect 10042 15348 10048 15360
rect 9999 15320 10048 15348
rect 9999 15317 10011 15320
rect 9953 15311 10011 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 11698 15348 11704 15360
rect 11659 15320 11704 15348
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 1581 15147 1639 15153
rect 1581 15144 1593 15147
rect 1544 15116 1593 15144
rect 1544 15104 1550 15116
rect 1581 15113 1593 15116
rect 1627 15113 1639 15147
rect 1581 15107 1639 15113
rect 2409 15147 2467 15153
rect 2409 15113 2421 15147
rect 2455 15144 2467 15147
rect 3142 15144 3148 15156
rect 2455 15116 3148 15144
rect 2455 15113 2467 15116
rect 2409 15107 2467 15113
rect 3142 15104 3148 15116
rect 3200 15104 3206 15156
rect 4706 15104 4712 15156
rect 4764 15144 4770 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 4764 15116 4813 15144
rect 4764 15104 4770 15116
rect 4801 15113 4813 15116
rect 4847 15144 4859 15147
rect 4847 15116 5764 15144
rect 4847 15113 4859 15116
rect 4801 15107 4859 15113
rect 4249 15079 4307 15085
rect 4249 15045 4261 15079
rect 4295 15076 4307 15079
rect 4982 15076 4988 15088
rect 4295 15048 4988 15076
rect 4295 15045 4307 15048
rect 4249 15039 4307 15045
rect 4982 15036 4988 15048
rect 5040 15036 5046 15088
rect 5736 15076 5764 15116
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 6604 15116 8217 15144
rect 6604 15104 6610 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8757 15147 8815 15153
rect 8757 15144 8769 15147
rect 8352 15116 8769 15144
rect 8352 15104 8358 15116
rect 8757 15113 8769 15116
rect 8803 15144 8815 15147
rect 9030 15144 9036 15156
rect 8803 15116 9036 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 10928 15116 11161 15144
rect 10928 15104 10934 15116
rect 11149 15113 11161 15116
rect 11195 15113 11207 15147
rect 11149 15107 11207 15113
rect 12253 15147 12311 15153
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 12342 15144 12348 15156
rect 12299 15116 12348 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 17402 15144 17408 15156
rect 17363 15116 17408 15144
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 20438 15144 20444 15156
rect 19659 15116 20444 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 6457 15079 6515 15085
rect 6457 15076 6469 15079
rect 5736 15048 6469 15076
rect 6457 15045 6469 15048
rect 6503 15076 6515 15079
rect 6641 15079 6699 15085
rect 6641 15076 6653 15079
rect 6503 15048 6653 15076
rect 6503 15045 6515 15048
rect 6457 15039 6515 15045
rect 6641 15045 6653 15048
rect 6687 15045 6699 15079
rect 6641 15039 6699 15045
rect 6273 15011 6331 15017
rect 6273 14977 6285 15011
rect 6319 15008 6331 15011
rect 6362 15008 6368 15020
rect 6319 14980 6368 15008
rect 6319 14977 6331 14980
rect 6273 14971 6331 14977
rect 6362 14968 6368 14980
rect 6420 15008 6426 15020
rect 6420 14980 6960 15008
rect 6420 14968 6426 14980
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 2682 14940 2688 14952
rect 1443 14912 2688 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 3142 14949 3148 14952
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14909 2927 14943
rect 3136 14940 3148 14949
rect 3055 14912 3148 14940
rect 2869 14903 2927 14909
rect 3136 14903 3148 14912
rect 3200 14940 3206 14952
rect 3878 14940 3884 14952
rect 3200 14912 3884 14940
rect 1670 14832 1676 14884
rect 1728 14872 1734 14884
rect 2041 14875 2099 14881
rect 2041 14872 2053 14875
rect 1728 14844 2053 14872
rect 1728 14832 1734 14844
rect 2041 14841 2053 14844
rect 2087 14872 2099 14875
rect 2777 14875 2835 14881
rect 2777 14872 2789 14875
rect 2087 14844 2789 14872
rect 2087 14841 2099 14844
rect 2041 14835 2099 14841
rect 2777 14841 2789 14844
rect 2823 14872 2835 14875
rect 2884 14872 2912 14903
rect 3142 14900 3148 14903
rect 3200 14900 3206 14912
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5442 14940 5448 14952
rect 5399 14912 5448 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 6454 14940 6460 14952
rect 6367 14912 6460 14940
rect 6454 14900 6460 14912
rect 6512 14940 6518 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6512 14912 6837 14940
rect 6512 14900 6518 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6932 14940 6960 14980
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16908 14980 16957 15008
rect 16908 14968 16914 14980
rect 16945 14977 16957 14980
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 7092 14943 7150 14949
rect 7092 14940 7104 14943
rect 6932 14912 7104 14940
rect 6825 14903 6883 14909
rect 7092 14909 7104 14912
rect 7138 14940 7150 14943
rect 7834 14940 7840 14952
rect 7138 14912 7840 14940
rect 7138 14909 7150 14912
rect 7092 14903 7150 14909
rect 4706 14872 4712 14884
rect 2823 14844 4712 14872
rect 2823 14841 2835 14844
rect 2777 14835 2835 14841
rect 4706 14832 4712 14844
rect 4764 14832 4770 14884
rect 6840 14872 6868 14903
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10318 14940 10324 14952
rect 9815 14912 10324 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 8938 14872 8944 14884
rect 6840 14844 8944 14872
rect 8938 14832 8944 14844
rect 8996 14872 9002 14884
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 8996 14844 9229 14872
rect 8996 14832 9002 14844
rect 9217 14841 9229 14844
rect 9263 14841 9275 14875
rect 9217 14835 9275 14841
rect 5258 14804 5264 14816
rect 5219 14776 5264 14804
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 9232 14804 9260 14835
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 9232 14776 9689 14804
rect 9677 14773 9689 14776
rect 9723 14804 9735 14807
rect 9784 14804 9812 14903
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14940 13875 14943
rect 13906 14940 13912 14952
rect 13863 14912 13912 14940
rect 13863 14909 13875 14912
rect 13817 14903 13875 14909
rect 13906 14900 13912 14912
rect 13964 14940 13970 14952
rect 19426 14940 19432 14952
rect 13964 14912 15516 14940
rect 19387 14912 19432 14940
rect 13964 14900 13970 14912
rect 10042 14881 10048 14884
rect 10036 14872 10048 14881
rect 9955 14844 10048 14872
rect 10036 14835 10048 14844
rect 10100 14872 10106 14884
rect 10686 14872 10692 14884
rect 10100 14844 10692 14872
rect 10042 14832 10048 14835
rect 10100 14832 10106 14844
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 12805 14875 12863 14881
rect 12805 14841 12817 14875
rect 12851 14872 12863 14875
rect 13170 14872 13176 14884
rect 12851 14844 13176 14872
rect 12851 14841 12863 14844
rect 12805 14835 12863 14841
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 13998 14832 14004 14884
rect 14056 14872 14062 14884
rect 14154 14875 14212 14881
rect 14154 14872 14166 14875
rect 14056 14844 14166 14872
rect 14056 14832 14062 14844
rect 14154 14841 14166 14844
rect 14200 14841 14212 14875
rect 14154 14835 14212 14841
rect 15488 14816 15516 14912
rect 19426 14900 19432 14912
rect 19484 14940 19490 14952
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19484 14912 19901 14940
rect 19484 14900 19490 14912
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 19889 14903 19947 14909
rect 15933 14875 15991 14881
rect 15933 14841 15945 14875
rect 15979 14872 15991 14875
rect 16758 14872 16764 14884
rect 15979 14844 16764 14872
rect 15979 14841 15991 14844
rect 15933 14835 15991 14841
rect 16758 14832 16764 14844
rect 16816 14832 16822 14884
rect 11882 14804 11888 14816
rect 9723 14776 11888 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 12894 14804 12900 14816
rect 12855 14776 12900 14804
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13354 14804 13360 14816
rect 13315 14776 13360 14804
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 15286 14804 15292 14816
rect 15247 14776 15292 14804
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 16206 14804 16212 14816
rect 15528 14776 16212 14804
rect 15528 14764 15534 14776
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16390 14804 16396 14816
rect 16351 14776 16396 14804
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 16540 14776 16865 14804
rect 16540 14764 16546 14776
rect 16853 14773 16865 14776
rect 16899 14804 16911 14807
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 16899 14776 17785 14804
rect 16899 14773 16911 14776
rect 16853 14767 16911 14773
rect 17773 14773 17785 14776
rect 17819 14773 17831 14807
rect 17773 14767 17831 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1762 14560 1768 14612
rect 1820 14600 1826 14612
rect 1857 14603 1915 14609
rect 1857 14600 1869 14603
rect 1820 14572 1869 14600
rect 1820 14560 1826 14572
rect 1857 14569 1869 14572
rect 1903 14569 1915 14603
rect 1857 14563 1915 14569
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 1872 14396 1900 14563
rect 2130 14560 2136 14612
rect 2188 14600 2194 14612
rect 2409 14603 2467 14609
rect 2409 14600 2421 14603
rect 2188 14572 2421 14600
rect 2188 14560 2194 14572
rect 2409 14569 2421 14572
rect 2455 14569 2467 14603
rect 2409 14563 2467 14569
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 4430 14600 4436 14612
rect 2740 14572 3924 14600
rect 4391 14572 4436 14600
rect 2740 14560 2746 14572
rect 2777 14535 2835 14541
rect 2777 14501 2789 14535
rect 2823 14532 2835 14535
rect 3326 14532 3332 14544
rect 2823 14504 3332 14532
rect 2823 14501 2835 14504
rect 2777 14495 2835 14501
rect 3326 14492 3332 14504
rect 3384 14532 3390 14544
rect 3786 14532 3792 14544
rect 3384 14504 3792 14532
rect 3384 14492 3390 14504
rect 3786 14492 3792 14504
rect 3844 14492 3850 14544
rect 3896 14541 3924 14572
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 4580 14572 4625 14600
rect 4580 14560 4586 14572
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 5316 14572 7481 14600
rect 5316 14560 5322 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 10042 14600 10048 14612
rect 10003 14572 10048 14600
rect 7469 14563 7527 14569
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10781 14603 10839 14609
rect 10781 14569 10793 14603
rect 10827 14600 10839 14603
rect 10870 14600 10876 14612
rect 10827 14572 10876 14600
rect 10827 14569 10839 14572
rect 10781 14563 10839 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 13998 14600 14004 14612
rect 13959 14572 14004 14600
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 15378 14600 15384 14612
rect 15335 14572 15384 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 16816 14572 16865 14600
rect 16816 14560 16822 14572
rect 16853 14569 16865 14572
rect 16899 14569 16911 14603
rect 16853 14563 16911 14569
rect 3881 14535 3939 14541
rect 3881 14501 3893 14535
rect 3927 14532 3939 14535
rect 4890 14532 4896 14544
rect 3927 14504 4896 14532
rect 3927 14501 3939 14504
rect 3881 14495 3939 14501
rect 4890 14492 4896 14504
rect 4948 14492 4954 14544
rect 6356 14535 6414 14541
rect 6356 14501 6368 14535
rect 6402 14532 6414 14535
rect 6546 14532 6552 14544
rect 6402 14504 6552 14532
rect 6402 14501 6414 14504
rect 6356 14495 6414 14501
rect 6546 14492 6552 14504
rect 6604 14492 6610 14544
rect 12066 14541 12072 14544
rect 12060 14532 12072 14541
rect 12027 14504 12072 14532
rect 12060 14495 12072 14504
rect 12066 14492 12072 14495
rect 12124 14492 12130 14544
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 16298 14532 16304 14544
rect 15252 14504 16304 14532
rect 15252 14492 15258 14504
rect 16298 14492 16304 14504
rect 16356 14492 16362 14544
rect 2869 14467 2927 14473
rect 2869 14433 2881 14467
rect 2915 14464 2927 14467
rect 3234 14464 3240 14476
rect 2915 14436 3240 14464
rect 2915 14433 2927 14436
rect 2869 14427 2927 14433
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 6086 14424 6092 14476
rect 6144 14473 6150 14476
rect 6144 14464 6154 14473
rect 8386 14464 8392 14476
rect 6144 14436 6189 14464
rect 8347 14436 8392 14464
rect 6144 14427 6154 14436
rect 6144 14424 6150 14427
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 10318 14464 10324 14476
rect 10183 14436 10324 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14464 11851 14467
rect 11882 14464 11888 14476
rect 11839 14436 11888 14464
rect 11839 14433 11851 14436
rect 11793 14427 11851 14433
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 16850 14464 16856 14476
rect 16807 14436 16856 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 1872 14368 3065 14396
rect 3053 14365 3065 14368
rect 3099 14396 3111 14399
rect 3142 14396 3148 14408
rect 3099 14368 3148 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3142 14356 3148 14368
rect 3200 14396 3206 14408
rect 4614 14396 4620 14408
rect 3200 14368 4200 14396
rect 4575 14368 4620 14396
rect 3200 14356 3206 14368
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 4065 14331 4123 14337
rect 4065 14328 4077 14331
rect 3292 14300 4077 14328
rect 3292 14288 3298 14300
rect 4065 14297 4077 14300
rect 4111 14297 4123 14331
rect 4065 14291 4123 14297
rect 2317 14263 2375 14269
rect 2317 14229 2329 14263
rect 2363 14260 2375 14263
rect 2498 14260 2504 14272
rect 2363 14232 2504 14260
rect 2363 14229 2375 14232
rect 2317 14223 2375 14229
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 3418 14260 3424 14272
rect 3379 14232 3424 14260
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 4172 14260 4200 14368
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 8570 14396 8576 14408
rect 8531 14368 8576 14396
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 10229 14359 10287 14365
rect 15028 14368 15761 14396
rect 9217 14331 9275 14337
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 9582 14328 9588 14340
rect 9263 14300 9588 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 9582 14288 9588 14300
rect 9640 14328 9646 14340
rect 10244 14328 10272 14359
rect 9640 14300 10272 14328
rect 9640 14288 9646 14300
rect 4982 14260 4988 14272
rect 4172 14232 4988 14260
rect 4982 14220 4988 14232
rect 5040 14260 5046 14272
rect 5077 14263 5135 14269
rect 5077 14260 5089 14263
rect 5040 14232 5089 14260
rect 5040 14220 5046 14232
rect 5077 14229 5089 14232
rect 5123 14229 5135 14263
rect 5442 14260 5448 14272
rect 5403 14232 5448 14260
rect 5077 14223 5135 14229
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5997 14263 6055 14269
rect 5997 14229 6009 14263
rect 6043 14260 6055 14263
rect 6362 14260 6368 14272
rect 6043 14232 6368 14260
rect 6043 14229 6055 14232
rect 5997 14223 6055 14229
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 7340 14232 8033 14260
rect 7340 14220 7346 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 9674 14260 9680 14272
rect 9635 14232 9680 14260
rect 8021 14223 8079 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 13170 14260 13176 14272
rect 13131 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13998 14220 14004 14272
rect 14056 14260 14062 14272
rect 15028 14269 15056 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 15856 14328 15884 14359
rect 15620 14300 15884 14328
rect 15620 14288 15626 14300
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14056 14232 15025 14260
rect 14056 14220 14062 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 4338 14056 4344 14068
rect 4299 14028 4344 14056
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 4488 14028 5365 14056
rect 4488 14016 4494 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 6178 14056 6184 14068
rect 6091 14028 6184 14056
rect 5353 14019 5411 14025
rect 4157 13991 4215 13997
rect 4157 13957 4169 13991
rect 4203 13988 4215 13991
rect 4522 13988 4528 14000
rect 4203 13960 4528 13988
rect 4203 13957 4215 13960
rect 4157 13951 4215 13957
rect 4522 13948 4528 13960
rect 4580 13948 4586 14000
rect 5368 13988 5396 14019
rect 6178 14016 6184 14028
rect 6236 14056 6242 14068
rect 6362 14056 6368 14068
rect 6236 14028 6368 14056
rect 6236 14016 6242 14028
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7377 14059 7435 14065
rect 7377 14056 7389 14059
rect 6972 14028 7389 14056
rect 6972 14016 6978 14028
rect 7377 14025 7389 14028
rect 7423 14025 7435 14059
rect 8938 14056 8944 14068
rect 8899 14028 8944 14056
rect 7377 14019 7435 14025
rect 7009 13991 7067 13997
rect 7009 13988 7021 13991
rect 5368 13960 7021 13988
rect 7009 13957 7021 13960
rect 7055 13957 7067 13991
rect 7009 13951 7067 13957
rect 2498 13920 2504 13932
rect 1412 13892 2504 13920
rect 1412 13861 1440 13892
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 2958 13920 2964 13932
rect 2731 13892 2964 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2958 13880 2964 13892
rect 3016 13920 3022 13932
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 3016 13892 3249 13920
rect 3016 13880 3022 13892
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3418 13920 3424 13932
rect 3379 13892 3424 13920
rect 3237 13883 3295 13889
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 4982 13920 4988 13932
rect 4943 13892 4988 13920
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 4798 13852 4804 13864
rect 4759 13824 4804 13852
rect 1397 13815 1455 13821
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 7024 13852 7052 13951
rect 7392 13920 7420 14019
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 10042 14016 10048 14068
rect 10100 14056 10106 14068
rect 11422 14056 11428 14068
rect 10100 14028 11428 14056
rect 10100 14016 10106 14028
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 12124 14028 12173 14056
rect 12124 14016 12130 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 14090 14016 14096 14068
rect 14148 14056 14154 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 14148 14028 15209 14056
rect 14148 14016 14154 14028
rect 8956 13988 8984 14016
rect 15028 14000 15056 14028
rect 15197 14025 15209 14028
rect 15243 14056 15255 14059
rect 15562 14056 15568 14068
rect 15243 14028 15568 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 15712 14028 15761 14056
rect 15712 14016 15718 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 15749 14019 15807 14025
rect 16301 14059 16359 14065
rect 16301 14025 16313 14059
rect 16347 14056 16359 14059
rect 16482 14056 16488 14068
rect 16347 14028 16488 14056
rect 16347 14025 16359 14028
rect 16301 14019 16359 14025
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 8956 13960 9168 13988
rect 8021 13923 8079 13929
rect 8021 13920 8033 13923
rect 7392 13892 8033 13920
rect 8021 13889 8033 13892
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 9140 13929 9168 13960
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 11149 13991 11207 13997
rect 11149 13988 11161 13991
rect 10376 13960 11161 13988
rect 10376 13948 10382 13960
rect 11149 13957 11161 13960
rect 11195 13988 11207 13991
rect 12710 13988 12716 14000
rect 11195 13960 12716 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 15010 13948 15016 14000
rect 15068 13948 15074 14000
rect 8205 13923 8263 13929
rect 8205 13920 8217 13923
rect 8168 13892 8217 13920
rect 8168 13880 8174 13892
rect 8205 13889 8217 13892
rect 8251 13920 8263 13923
rect 9125 13923 9183 13929
rect 8251 13892 9076 13920
rect 8251 13889 8263 13892
rect 8205 13883 8263 13889
rect 7466 13852 7472 13864
rect 7024 13824 7472 13852
rect 7466 13812 7472 13824
rect 7524 13852 7530 13864
rect 7929 13855 7987 13861
rect 7929 13852 7941 13855
rect 7524 13824 7941 13852
rect 7524 13812 7530 13824
rect 7929 13821 7941 13824
rect 7975 13821 7987 13855
rect 7929 13815 7987 13821
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8352 13824 8585 13852
rect 8352 13812 8358 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 2317 13787 2375 13793
rect 2317 13753 2329 13787
rect 2363 13784 2375 13787
rect 3145 13787 3203 13793
rect 3145 13784 3157 13787
rect 2363 13756 3157 13784
rect 2363 13753 2375 13756
rect 2317 13747 2375 13753
rect 3145 13753 3157 13756
rect 3191 13784 3203 13787
rect 4062 13784 4068 13796
rect 3191 13756 4068 13784
rect 3191 13753 3203 13756
rect 3145 13747 3203 13753
rect 4062 13744 4068 13756
rect 4120 13744 4126 13796
rect 9048 13784 9076 13892
rect 9125 13889 9137 13923
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 13354 13920 13360 13932
rect 12483 13892 13360 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 16356 13892 16773 13920
rect 16356 13880 16362 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13920 17003 13923
rect 17034 13920 17040 13932
rect 16991 13892 17040 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 17034 13880 17040 13892
rect 17092 13920 17098 13932
rect 17420 13920 17448 14016
rect 17092 13892 17448 13920
rect 17092 13880 17098 13892
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13504 13824 13737 13852
rect 13504 13812 13510 13824
rect 13725 13821 13737 13824
rect 13771 13852 13783 13855
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13771 13824 13829 13852
rect 13771 13821 13783 13824
rect 13725 13815 13783 13821
rect 13817 13821 13829 13824
rect 13863 13852 13875 13855
rect 13906 13852 13912 13864
rect 13863 13824 13912 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 9392 13787 9450 13793
rect 9392 13784 9404 13787
rect 9048 13756 9404 13784
rect 9392 13753 9404 13756
rect 9438 13784 9450 13787
rect 9582 13784 9588 13796
rect 9438 13756 9588 13784
rect 9438 13753 9450 13756
rect 9392 13747 9450 13753
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 13357 13787 13415 13793
rect 13357 13753 13369 13787
rect 13403 13784 13415 13787
rect 14084 13787 14142 13793
rect 14084 13784 14096 13787
rect 13403 13756 14096 13784
rect 13403 13753 13415 13756
rect 13357 13747 13415 13753
rect 14084 13753 14096 13756
rect 14130 13784 14142 13787
rect 14642 13784 14648 13796
rect 14130 13756 14648 13784
rect 14130 13753 14142 13756
rect 14084 13747 14142 13753
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 2777 13719 2835 13725
rect 2777 13716 2789 13719
rect 2648 13688 2789 13716
rect 2648 13676 2654 13688
rect 2777 13685 2789 13688
rect 2823 13685 2835 13719
rect 4706 13716 4712 13728
rect 4667 13688 4712 13716
rect 2777 13679 2835 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 5534 13676 5540 13728
rect 5592 13716 5598 13728
rect 5721 13719 5779 13725
rect 5721 13716 5733 13719
rect 5592 13688 5733 13716
rect 5592 13676 5598 13688
rect 5721 13685 5733 13688
rect 5767 13685 5779 13719
rect 7558 13716 7564 13728
rect 7519 13688 7564 13716
rect 5721 13679 5779 13685
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10686 13716 10692 13728
rect 10551 13688 10692 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 11882 13716 11888 13728
rect 11843 13688 11888 13716
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 16114 13716 16120 13728
rect 16075 13688 16120 13716
rect 16114 13676 16120 13688
rect 16172 13716 16178 13728
rect 16669 13719 16727 13725
rect 16669 13716 16681 13719
rect 16172 13688 16681 13716
rect 16172 13676 16178 13688
rect 16669 13685 16681 13688
rect 16715 13685 16727 13719
rect 16669 13679 16727 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 842 13472 848 13524
rect 900 13512 906 13524
rect 3142 13512 3148 13524
rect 900 13484 3004 13512
rect 3103 13484 3148 13512
rect 900 13472 906 13484
rect 2501 13447 2559 13453
rect 2501 13413 2513 13447
rect 2547 13444 2559 13447
rect 2590 13444 2596 13456
rect 2547 13416 2596 13444
rect 2547 13413 2559 13416
rect 2501 13407 2559 13413
rect 2590 13404 2596 13416
rect 2648 13404 2654 13456
rect 2976 13444 3004 13484
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 3878 13512 3884 13524
rect 3839 13484 3884 13512
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4304 13484 4445 13512
rect 4304 13472 4310 13484
rect 4433 13481 4445 13484
rect 4479 13481 4491 13515
rect 4433 13475 4491 13481
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 5077 13515 5135 13521
rect 5077 13512 5089 13515
rect 4764 13484 5089 13512
rect 4764 13472 4770 13484
rect 5077 13481 5089 13484
rect 5123 13481 5135 13515
rect 5077 13475 5135 13481
rect 5905 13515 5963 13521
rect 5905 13481 5917 13515
rect 5951 13512 5963 13515
rect 5994 13512 6000 13524
rect 5951 13484 6000 13512
rect 5951 13481 5963 13484
rect 5905 13475 5963 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6270 13512 6276 13524
rect 6231 13484 6276 13512
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 7650 13512 7656 13524
rect 7611 13484 7656 13512
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 8110 13512 8116 13524
rect 8071 13484 8116 13512
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 9950 13512 9956 13524
rect 9723 13484 9956 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 10134 13512 10140 13524
rect 10095 13484 10140 13512
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14001 13515 14059 13521
rect 14001 13512 14013 13515
rect 13872 13484 14013 13512
rect 13872 13472 13878 13484
rect 14001 13481 14013 13484
rect 14047 13481 14059 13515
rect 15010 13512 15016 13524
rect 14971 13484 15016 13512
rect 14001 13475 14059 13481
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 16945 13515 17003 13521
rect 16945 13481 16957 13515
rect 16991 13512 17003 13515
rect 17034 13512 17040 13524
rect 16991 13484 17040 13512
rect 16991 13481 17003 13484
rect 16945 13475 17003 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 19426 13512 19432 13524
rect 19387 13484 19432 13512
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 21085 13515 21143 13521
rect 21085 13481 21097 13515
rect 21131 13512 21143 13515
rect 21174 13512 21180 13524
rect 21131 13484 21180 13512
rect 21131 13481 21143 13484
rect 21085 13475 21143 13481
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 4525 13447 4583 13453
rect 4525 13444 4537 13447
rect 2976 13416 4537 13444
rect 4525 13413 4537 13416
rect 4571 13444 4583 13447
rect 4614 13444 4620 13456
rect 4571 13416 4620 13444
rect 4571 13413 4583 13416
rect 4525 13407 4583 13413
rect 4614 13404 4620 13416
rect 4672 13444 4678 13456
rect 7098 13444 7104 13456
rect 4672 13416 7104 13444
rect 4672 13404 4678 13416
rect 7098 13404 7104 13416
rect 7156 13444 7162 13456
rect 7282 13444 7288 13456
rect 7156 13416 7288 13444
rect 7156 13404 7162 13416
rect 7282 13404 7288 13416
rect 7340 13404 7346 13456
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 5813 13379 5871 13385
rect 2004 13348 2728 13376
rect 2004 13336 2010 13348
rect 2700 13317 2728 13348
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 7469 13379 7527 13385
rect 5859 13348 6592 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 6564 13320 6592 13348
rect 7469 13345 7481 13379
rect 7515 13376 7527 13379
rect 7834 13376 7840 13388
rect 7515 13348 7840 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8754 13336 8760 13388
rect 8812 13376 8818 13388
rect 9674 13376 9680 13388
rect 8812 13348 9680 13376
rect 8812 13336 8818 13348
rect 9674 13336 9680 13348
rect 9732 13376 9738 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9732 13348 10057 13376
rect 9732 13336 9738 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 12233 13379 12291 13385
rect 12233 13376 12245 13379
rect 11572 13348 12245 13376
rect 11572 13336 11578 13348
rect 12233 13345 12245 13348
rect 12279 13376 12291 13379
rect 13170 13376 13176 13388
rect 12279 13348 13176 13376
rect 12279 13345 12291 13348
rect 12233 13339 12291 13345
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 15832 13379 15890 13385
rect 15832 13345 15844 13379
rect 15878 13376 15890 13379
rect 16206 13376 16212 13388
rect 15878 13348 16212 13376
rect 15878 13345 15890 13348
rect 15832 13339 15890 13345
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 18138 13336 18144 13388
rect 18196 13376 18202 13388
rect 18305 13379 18363 13385
rect 18305 13376 18317 13379
rect 18196 13348 18317 13376
rect 18196 13336 18202 13348
rect 18305 13345 18317 13348
rect 18351 13345 18363 13379
rect 18305 13339 18363 13345
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20864 13348 20913 13376
rect 20864 13336 20870 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 2608 13240 2636 13271
rect 2608 13212 3924 13240
rect 3896 13184 3924 13212
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 4632 13240 4660 13271
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 6236 13280 6377 13308
rect 6236 13268 6242 13280
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 6546 13308 6552 13320
rect 6507 13280 6552 13308
rect 6365 13271 6423 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 8570 13308 8576 13320
rect 8531 13280 8576 13308
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 10226 13308 10232 13320
rect 10187 13280 10232 13308
rect 10226 13268 10232 13280
rect 10284 13308 10290 13320
rect 10686 13308 10692 13320
rect 10284 13280 10692 13308
rect 10284 13268 10290 13280
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11940 13280 11989 13308
rect 11940 13268 11946 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 15562 13308 15568 13320
rect 15523 13280 15568 13308
rect 11977 13271 12035 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 18012 13280 18061 13308
rect 18012 13268 18018 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 4028 13212 4660 13240
rect 4028 13200 4034 13212
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 2222 13172 2228 13184
rect 2179 13144 2228 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 3878 13132 3884 13184
rect 3936 13172 3942 13184
rect 4065 13175 4123 13181
rect 4065 13172 4077 13175
rect 3936 13144 4077 13172
rect 3936 13132 3942 13144
rect 4065 13141 4077 13144
rect 4111 13141 4123 13175
rect 7006 13172 7012 13184
rect 6967 13144 7012 13172
rect 4065 13135 4123 13141
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7282 13172 7288 13184
rect 7243 13144 7288 13172
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 9493 13175 9551 13181
rect 9493 13141 9505 13175
rect 9539 13172 9551 13175
rect 9582 13172 9588 13184
rect 9539 13144 9588 13172
rect 9539 13141 9551 13144
rect 9493 13135 9551 13141
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 13354 13172 13360 13184
rect 13315 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 3970 12968 3976 12980
rect 3568 12940 3976 12968
rect 3568 12928 3574 12940
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4580 12940 4997 12968
rect 4580 12928 4586 12940
rect 4985 12937 4997 12940
rect 5031 12968 5043 12971
rect 5031 12940 5672 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 4614 12900 4620 12912
rect 4575 12872 4620 12900
rect 4614 12860 4620 12872
rect 4672 12900 4678 12912
rect 5074 12900 5080 12912
rect 4672 12872 5080 12900
rect 4672 12860 4678 12872
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 5644 12900 5672 12940
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 6328 12940 6561 12968
rect 6328 12928 6334 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 6549 12931 6607 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9214 12968 9220 12980
rect 9175 12940 9220 12968
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10192 12940 10609 12968
rect 10192 12928 10198 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 11514 12968 11520 12980
rect 11475 12940 11520 12968
rect 10597 12931 10655 12937
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12158 12968 12164 12980
rect 12119 12940 12164 12968
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13998 12968 14004 12980
rect 12492 12940 12537 12968
rect 13959 12940 14004 12968
rect 12492 12928 12498 12940
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 15988 12940 16405 12968
rect 15988 12928 15994 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 16393 12931 16451 12937
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 22002 12968 22008 12980
rect 21315 12940 22008 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 22465 12971 22523 12977
rect 22465 12937 22477 12971
rect 22511 12968 22523 12971
rect 23382 12968 23388 12980
rect 22511 12940 23388 12968
rect 22511 12937 22523 12940
rect 22465 12931 22523 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 6822 12900 6828 12912
rect 5644 12872 6828 12900
rect 2590 12832 2596 12844
rect 2551 12804 2596 12832
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 5644 12841 5672 12872
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5810 12832 5816 12844
rect 5771 12804 5816 12832
rect 5629 12795 5687 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7064 12804 7389 12832
rect 7064 12792 7070 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9364 12804 9781 12832
rect 9364 12792 9370 12804
rect 9769 12801 9781 12804
rect 9815 12832 9827 12835
rect 10226 12832 10232 12844
rect 9815 12804 10232 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 12526 12792 12532 12844
rect 12584 12832 12590 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12584 12804 12909 12832
rect 12584 12792 12590 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 13078 12832 13084 12844
rect 13039 12804 13084 12832
rect 12897 12795 12955 12801
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12832 13599 12835
rect 14642 12832 14648 12844
rect 13587 12804 14648 12832
rect 13587 12801 13599 12804
rect 13541 12795 13599 12801
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 17034 12832 17040 12844
rect 16995 12804 17040 12832
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1578 12764 1584 12776
rect 1443 12736 1584 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 2130 12764 2136 12776
rect 2043 12736 2136 12764
rect 2130 12724 2136 12736
rect 2188 12764 2194 12776
rect 2849 12767 2907 12773
rect 2849 12764 2861 12767
rect 2188 12736 2861 12764
rect 2188 12724 2194 12736
rect 2849 12733 2861 12736
rect 2895 12733 2907 12767
rect 2849 12727 2907 12733
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 4522 12764 4528 12776
rect 3384 12736 4528 12764
rect 3384 12724 3390 12736
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12764 5595 12767
rect 5718 12764 5724 12776
rect 5583 12736 5724 12764
rect 5583 12733 5595 12736
rect 5537 12727 5595 12733
rect 5718 12724 5724 12736
rect 5776 12764 5782 12776
rect 6362 12764 6368 12776
rect 5776 12736 6368 12764
rect 5776 12724 5782 12736
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 9674 12764 9680 12776
rect 8435 12736 9680 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12216 12736 12817 12764
rect 12216 12724 12222 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 13872 12736 14473 12764
rect 13872 12724 13878 12736
rect 14461 12733 14473 12736
rect 14507 12733 14519 12767
rect 14461 12727 14519 12733
rect 18138 12724 18144 12776
rect 18196 12764 18202 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18196 12736 18889 12764
rect 18196 12724 18202 12736
rect 18877 12733 18889 12736
rect 18923 12733 18935 12767
rect 18877 12727 18935 12733
rect 20806 12724 20812 12776
rect 20864 12764 20870 12776
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 20864 12736 20913 12764
rect 20864 12724 20870 12736
rect 20901 12733 20913 12736
rect 20947 12733 20959 12767
rect 21082 12764 21088 12776
rect 20995 12736 21088 12764
rect 20901 12727 20959 12733
rect 21082 12724 21088 12736
rect 21140 12764 21146 12776
rect 21545 12767 21603 12773
rect 21545 12764 21557 12767
rect 21140 12736 21557 12764
rect 21140 12724 21146 12736
rect 21545 12733 21557 12736
rect 21591 12733 21603 12767
rect 22278 12764 22284 12776
rect 22239 12736 22284 12764
rect 21545 12727 21603 12733
rect 22278 12724 22284 12736
rect 22336 12764 22342 12776
rect 22741 12767 22799 12773
rect 22741 12764 22753 12767
rect 22336 12736 22753 12764
rect 22336 12724 22342 12736
rect 22741 12733 22753 12736
rect 22787 12733 22799 12767
rect 22741 12727 22799 12733
rect 7282 12696 7288 12708
rect 5184 12668 7288 12696
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2590 12628 2596 12640
rect 2547 12600 2596 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2590 12588 2596 12600
rect 2648 12628 2654 12640
rect 2958 12628 2964 12640
rect 2648 12600 2964 12628
rect 2648 12588 2654 12600
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 5184 12637 5212 12668
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 9125 12699 9183 12705
rect 9125 12665 9137 12699
rect 9171 12696 9183 12699
rect 9585 12699 9643 12705
rect 9585 12696 9597 12699
rect 9171 12668 9597 12696
rect 9171 12665 9183 12668
rect 9125 12659 9183 12665
rect 9585 12665 9597 12668
rect 9631 12696 9643 12699
rect 10781 12699 10839 12705
rect 10781 12696 10793 12699
rect 9631 12668 10793 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 10781 12665 10793 12668
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 13909 12699 13967 12705
rect 13909 12665 13921 12699
rect 13955 12696 13967 12699
rect 14366 12696 14372 12708
rect 13955 12668 14372 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 14366 12656 14372 12668
rect 14424 12656 14430 12708
rect 15289 12699 15347 12705
rect 15289 12665 15301 12699
rect 15335 12696 15347 12699
rect 16206 12696 16212 12708
rect 15335 12668 16212 12696
rect 15335 12665 15347 12668
rect 15289 12659 15347 12665
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 16301 12699 16359 12705
rect 16301 12665 16313 12699
rect 16347 12696 16359 12699
rect 16761 12699 16819 12705
rect 16761 12696 16773 12699
rect 16347 12668 16773 12696
rect 16347 12665 16359 12668
rect 16301 12659 16359 12665
rect 16761 12665 16773 12668
rect 16807 12696 16819 12699
rect 18049 12699 18107 12705
rect 18049 12696 18061 12699
rect 16807 12668 18061 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 18049 12665 18061 12668
rect 18095 12665 18107 12699
rect 18049 12659 18107 12665
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12597 5227 12631
rect 6178 12628 6184 12640
rect 6139 12600 6184 12628
rect 5169 12591 5227 12597
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7190 12628 7196 12640
rect 7151 12600 7196 12628
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 7834 12628 7840 12640
rect 7795 12600 7840 12628
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 15657 12631 15715 12637
rect 15657 12628 15669 12631
rect 15620 12600 15669 12628
rect 15620 12588 15626 12600
rect 15657 12597 15669 12600
rect 15703 12628 15715 12631
rect 15930 12628 15936 12640
rect 15703 12600 15936 12628
rect 15703 12597 15715 12600
rect 15657 12591 15715 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16482 12588 16488 12640
rect 16540 12628 16546 12640
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 16540 12600 16865 12628
rect 16540 12588 16546 12600
rect 16853 12597 16865 12600
rect 16899 12628 16911 12631
rect 17405 12631 17463 12637
rect 17405 12628 17417 12631
rect 16899 12600 17417 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17405 12597 17417 12600
rect 17451 12597 17463 12631
rect 17405 12591 17463 12597
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18509 12631 18567 12637
rect 18509 12628 18521 12631
rect 18012 12600 18521 12628
rect 18012 12588 18018 12600
rect 18509 12597 18521 12600
rect 18555 12597 18567 12631
rect 18509 12591 18567 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3234 12424 3240 12436
rect 3195 12396 3240 12424
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 3970 12424 3976 12436
rect 3927 12396 3976 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 2869 12359 2927 12365
rect 2869 12356 2881 12359
rect 2832 12328 2881 12356
rect 2832 12316 2838 12328
rect 2869 12325 2881 12328
rect 2915 12356 2927 12359
rect 3896 12356 3924 12387
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4246 12424 4252 12436
rect 4207 12396 4252 12424
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4617 12427 4675 12433
rect 4617 12424 4629 12427
rect 4396 12396 4629 12424
rect 4396 12384 4402 12396
rect 4617 12393 4629 12396
rect 4663 12393 4675 12427
rect 6822 12424 6828 12436
rect 6783 12396 6828 12424
rect 4617 12387 4675 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 9306 12424 9312 12436
rect 9267 12396 9312 12424
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 11238 12424 11244 12436
rect 11199 12396 11244 12424
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11609 12427 11667 12433
rect 11609 12393 11621 12427
rect 11655 12424 11667 12427
rect 11698 12424 11704 12436
rect 11655 12396 11704 12424
rect 11655 12393 11667 12396
rect 11609 12387 11667 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12526 12424 12532 12436
rect 12487 12396 12532 12424
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 12897 12427 12955 12433
rect 12897 12393 12909 12427
rect 12943 12424 12955 12427
rect 13078 12424 13084 12436
rect 12943 12396 13084 12424
rect 12943 12393 12955 12396
rect 12897 12387 12955 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13357 12427 13415 12433
rect 13357 12393 13369 12427
rect 13403 12424 13415 12427
rect 13446 12424 13452 12436
rect 13403 12396 13452 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 15841 12427 15899 12433
rect 15841 12393 15853 12427
rect 15887 12393 15899 12427
rect 16390 12424 16396 12436
rect 16351 12396 16396 12424
rect 15841 12387 15899 12393
rect 2915 12328 3924 12356
rect 2915 12325 2927 12328
rect 2869 12319 2927 12325
rect 5534 12316 5540 12368
rect 5592 12356 5598 12368
rect 5690 12359 5748 12365
rect 5690 12356 5702 12359
rect 5592 12328 5702 12356
rect 5592 12316 5598 12328
rect 5690 12325 5702 12328
rect 5736 12356 5748 12359
rect 5810 12356 5816 12368
rect 5736 12328 5816 12356
rect 5736 12325 5748 12328
rect 5690 12319 5748 12325
rect 5810 12316 5816 12328
rect 5868 12316 5874 12368
rect 8570 12316 8576 12368
rect 8628 12316 8634 12368
rect 10134 12356 10140 12368
rect 10095 12328 10140 12356
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 15856 12356 15884 12387
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 21913 12427 21971 12433
rect 21913 12393 21925 12427
rect 21959 12424 21971 12427
rect 22738 12424 22744 12436
rect 21959 12396 22744 12424
rect 21959 12393 21971 12396
rect 21913 12387 21971 12393
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 16666 12356 16672 12368
rect 15856 12328 16672 12356
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 16936 12359 16994 12365
rect 16936 12325 16948 12359
rect 16982 12356 16994 12359
rect 17126 12356 17132 12368
rect 16982 12328 17132 12356
rect 16982 12325 16994 12328
rect 16936 12319 16994 12325
rect 17126 12316 17132 12328
rect 17184 12316 17190 12368
rect 2130 12288 2136 12300
rect 2091 12260 2136 12288
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2222 12248 2228 12300
rect 2280 12288 2286 12300
rect 2682 12288 2688 12300
rect 2280 12260 2688 12288
rect 2280 12248 2286 12260
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4154 12288 4160 12300
rect 4111 12260 4160 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 5258 12288 5264 12300
rect 5219 12260 5264 12288
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 6454 12288 6460 12300
rect 5491 12260 6460 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 6454 12248 6460 12260
rect 6512 12248 6518 12300
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 8260 12260 8309 12288
rect 8260 12248 8266 12260
rect 8297 12257 8309 12260
rect 8343 12288 8355 12291
rect 8588 12288 8616 12316
rect 8343 12260 8616 12288
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 10008 12260 10057 12288
rect 10008 12248 10014 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11572 12260 11713 12288
rect 11572 12248 11578 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 14001 12291 14059 12297
rect 14001 12288 14013 12291
rect 13136 12260 14013 12288
rect 13136 12248 13142 12260
rect 14001 12257 14013 12260
rect 14047 12257 14059 12291
rect 14001 12251 14059 12257
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15528 12260 15669 12288
rect 15528 12248 15534 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 21726 12288 21732 12300
rect 21687 12260 21732 12288
rect 15657 12251 15715 12257
rect 21726 12248 21732 12260
rect 21784 12248 21790 12300
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2590 12220 2596 12232
rect 2455 12192 2596 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10778 12220 10784 12232
rect 10367 12192 10784 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12152 1731 12155
rect 2038 12152 2044 12164
rect 1719 12124 2044 12152
rect 1719 12121 1731 12124
rect 1673 12115 1731 12121
rect 2038 12112 2044 12124
rect 2096 12112 2102 12164
rect 7742 12152 7748 12164
rect 7703 12124 7748 12152
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 10336 12152 10364 12183
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11790 12220 11796 12232
rect 11751 12192 11796 12220
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13814 12220 13820 12232
rect 12768 12192 13820 12220
rect 12768 12180 12774 12192
rect 13814 12180 13820 12192
rect 13872 12220 13878 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13872 12192 14105 12220
rect 13872 12180 13878 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14642 12220 14648 12232
rect 14323 12192 14648 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15930 12220 15936 12232
rect 15344 12192 15936 12220
rect 15344 12180 15350 12192
rect 15930 12180 15936 12192
rect 15988 12220 15994 12232
rect 16666 12220 16672 12232
rect 15988 12192 16672 12220
rect 15988 12180 15994 12192
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 9732 12124 10364 12152
rect 9732 12112 9738 12124
rect 17954 12112 17960 12164
rect 18012 12152 18018 12164
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 18012 12124 18061 12152
rect 18012 12112 18018 12124
rect 18049 12121 18061 12124
rect 18095 12121 18107 12155
rect 18049 12115 18107 12121
rect 1762 12084 1768 12096
rect 1723 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 7469 12087 7527 12093
rect 7469 12053 7481 12087
rect 7515 12084 7527 12087
rect 7558 12084 7564 12096
rect 7515 12056 7564 12084
rect 7515 12053 7527 12056
rect 7469 12047 7527 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 7926 12084 7932 12096
rect 7887 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 13630 12084 13636 12096
rect 13591 12056 13636 12084
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 15470 12084 15476 12096
rect 15431 12056 15476 12084
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 1636 11852 4077 11880
rect 1636 11840 1642 11852
rect 4065 11849 4077 11852
rect 4111 11880 4123 11883
rect 4154 11880 4160 11892
rect 4111 11852 4160 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5166 11880 5172 11892
rect 5127 11852 5172 11880
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 6273 11883 6331 11889
rect 6273 11880 6285 11883
rect 6236 11852 6285 11880
rect 6236 11840 6242 11852
rect 6273 11849 6285 11852
rect 6319 11880 6331 11883
rect 6454 11880 6460 11892
rect 6319 11852 6460 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 6454 11840 6460 11852
rect 6512 11880 6518 11892
rect 8297 11883 8355 11889
rect 8297 11880 8309 11883
rect 6512 11852 8309 11880
rect 6512 11840 6518 11852
rect 8297 11849 8309 11852
rect 8343 11849 8355 11883
rect 8297 11843 8355 11849
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 7837 11815 7895 11821
rect 7837 11812 7849 11815
rect 7156 11784 7849 11812
rect 7156 11772 7162 11784
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5534 11744 5540 11756
rect 4755 11716 5540 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5534 11704 5540 11716
rect 5592 11744 5598 11756
rect 7300 11753 7328 11784
rect 7837 11781 7849 11784
rect 7883 11781 7895 11815
rect 7837 11775 7895 11781
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 5592 11716 5733 11744
rect 5592 11704 5598 11716
rect 5721 11713 5733 11716
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11744 7343 11747
rect 7469 11747 7527 11753
rect 7331 11716 7365 11744
rect 7331 11713 7343 11716
rect 7285 11707 7343 11713
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 7558 11744 7564 11756
rect 7515 11716 7564 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 8312 11744 8340 11843
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10781 11883 10839 11889
rect 10781 11880 10793 11883
rect 10192 11852 10793 11880
rect 10192 11840 10198 11852
rect 10781 11849 10793 11852
rect 10827 11849 10839 11883
rect 11238 11880 11244 11892
rect 11151 11852 11244 11880
rect 10781 11843 10839 11849
rect 11238 11840 11244 11852
rect 11296 11880 11302 11892
rect 11790 11880 11796 11892
rect 11296 11852 11796 11880
rect 11296 11840 11302 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12710 11880 12716 11892
rect 12671 11852 12716 11880
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 16025 11883 16083 11889
rect 16025 11849 16037 11883
rect 16071 11880 16083 11883
rect 16482 11880 16488 11892
rect 16071 11852 16488 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 17129 11883 17187 11889
rect 17129 11880 17141 11883
rect 16724 11852 17141 11880
rect 16724 11840 16730 11852
rect 17129 11849 17141 11852
rect 17175 11880 17187 11883
rect 17862 11880 17868 11892
rect 17175 11852 17868 11880
rect 17175 11849 17187 11852
rect 17129 11843 17187 11849
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18046 11880 18052 11892
rect 18007 11852 18052 11880
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8312 11716 8493 11744
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 16298 11744 16304 11756
rect 15611 11716 16304 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 16298 11704 16304 11716
rect 16356 11744 16362 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 16356 11716 16497 11744
rect 16356 11704 16362 11716
rect 16485 11713 16497 11716
rect 16531 11713 16543 11747
rect 16485 11707 16543 11713
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11744 16727 11747
rect 17126 11744 17132 11756
rect 16715 11716 17132 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 1946 11676 1952 11688
rect 1859 11648 1952 11676
rect 1946 11636 1952 11648
rect 2004 11676 2010 11688
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 2004 11648 2053 11676
rect 2004 11636 2010 11648
rect 2041 11645 2053 11648
rect 2087 11645 2099 11679
rect 2041 11639 2099 11645
rect 2308 11679 2366 11685
rect 2308 11645 2320 11679
rect 2354 11676 2366 11679
rect 2774 11676 2780 11688
rect 2354 11648 2780 11676
rect 2354 11645 2366 11648
rect 2308 11639 2366 11645
rect 2056 11608 2084 11639
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 8570 11636 8576 11688
rect 8628 11676 8634 11688
rect 8737 11679 8795 11685
rect 8737 11676 8749 11679
rect 8628 11648 8749 11676
rect 8628 11636 8634 11648
rect 8737 11645 8749 11648
rect 8783 11645 8795 11679
rect 8737 11639 8795 11645
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11676 13323 11679
rect 13354 11676 13360 11688
rect 13311 11648 13360 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 18506 11676 18512 11688
rect 18467 11648 18512 11676
rect 18506 11636 18512 11648
rect 18564 11676 18570 11688
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 18564 11648 19073 11676
rect 18564 11636 18570 11648
rect 19061 11645 19073 11648
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 2958 11608 2964 11620
rect 2056 11580 2964 11608
rect 2958 11568 2964 11580
rect 3016 11568 3022 11620
rect 3694 11568 3700 11620
rect 3752 11608 3758 11620
rect 4985 11611 5043 11617
rect 4985 11608 4997 11611
rect 3752 11580 4997 11608
rect 3752 11568 3758 11580
rect 4985 11577 4997 11580
rect 5031 11608 5043 11611
rect 5629 11611 5687 11617
rect 5629 11608 5641 11611
rect 5031 11580 5641 11608
rect 5031 11577 5043 11580
rect 4985 11571 5043 11577
rect 5629 11577 5641 11580
rect 5675 11577 5687 11611
rect 6546 11608 6552 11620
rect 6507 11580 6552 11608
rect 5629 11571 5687 11577
rect 6546 11568 6552 11580
rect 6604 11608 6610 11620
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 6604 11580 7205 11608
rect 6604 11568 6610 11580
rect 7193 11577 7205 11580
rect 7239 11577 7251 11611
rect 7193 11571 7251 11577
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 9950 11608 9956 11620
rect 9732 11580 9956 11608
rect 9732 11568 9738 11580
rect 9950 11568 9956 11580
rect 10008 11608 10014 11620
rect 10413 11611 10471 11617
rect 10413 11608 10425 11611
rect 10008 11580 10425 11608
rect 10008 11568 10014 11580
rect 10413 11577 10425 11580
rect 10459 11577 10471 11611
rect 10413 11571 10471 11577
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11514 11608 11520 11620
rect 11112 11580 11520 11608
rect 11112 11568 11118 11580
rect 11514 11568 11520 11580
rect 11572 11608 11578 11620
rect 13538 11617 13544 11620
rect 12161 11611 12219 11617
rect 12161 11608 12173 11611
rect 11572 11580 12173 11608
rect 11572 11568 11578 11580
rect 12161 11577 12173 11580
rect 12207 11577 12219 11611
rect 13532 11608 13544 11617
rect 13499 11580 13544 11608
rect 12161 11571 12219 11577
rect 13532 11571 13544 11580
rect 13538 11568 13544 11571
rect 13596 11568 13602 11620
rect 16574 11568 16580 11620
rect 16632 11608 16638 11620
rect 17773 11611 17831 11617
rect 17773 11608 17785 11611
rect 16632 11580 17785 11608
rect 16632 11568 16638 11580
rect 17773 11577 17785 11580
rect 17819 11608 17831 11611
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 17819 11580 18429 11608
rect 17819 11577 17831 11580
rect 17773 11571 17831 11577
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18417 11571 18475 11577
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 3421 11543 3479 11549
rect 3421 11540 3433 11543
rect 2096 11512 3433 11540
rect 2096 11500 2102 11512
rect 3421 11509 3433 11512
rect 3467 11509 3479 11543
rect 3421 11503 3479 11509
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 5537 11543 5595 11549
rect 5537 11540 5549 11543
rect 5500 11512 5549 11540
rect 5500 11500 5506 11512
rect 5537 11509 5549 11512
rect 5583 11509 5595 11543
rect 5537 11503 5595 11509
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 9858 11540 9864 11552
rect 9819 11512 9864 11540
rect 6825 11503 6883 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 11330 11540 11336 11552
rect 11291 11512 11336 11540
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 14642 11540 14648 11552
rect 14603 11512 14648 11540
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 15841 11543 15899 11549
rect 15841 11540 15853 11543
rect 15620 11512 15853 11540
rect 15620 11500 15626 11512
rect 15841 11509 15853 11512
rect 15887 11540 15899 11543
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 15887 11512 16405 11540
rect 15887 11509 15899 11512
rect 15841 11503 15899 11509
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 17184 11512 17417 11540
rect 17184 11500 17190 11512
rect 17405 11509 17417 11512
rect 17451 11509 17463 11543
rect 21726 11540 21732 11552
rect 21687 11512 21732 11540
rect 17405 11503 17463 11509
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1854 11336 1860 11348
rect 1627 11308 1860 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2004 11308 2049 11336
rect 2004 11296 2010 11308
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2280 11308 2421 11336
rect 2280 11296 2286 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2869 11339 2927 11345
rect 2409 11299 2467 11305
rect 2700 11308 2820 11336
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2700 11200 2728 11308
rect 2792 11268 2820 11308
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3326 11336 3332 11348
rect 2915 11308 3332 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 3510 11336 3516 11348
rect 3471 11308 3516 11336
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 5534 11336 5540 11348
rect 5495 11308 5540 11336
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5994 11336 6000 11348
rect 5955 11308 6000 11336
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 8202 11336 8208 11348
rect 8163 11308 8208 11336
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11336 8634 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 8628 11308 8861 11336
rect 8628 11296 8634 11308
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 8849 11299 8907 11305
rect 9861 11339 9919 11345
rect 9861 11305 9873 11339
rect 9907 11336 9919 11339
rect 11790 11336 11796 11348
rect 9907 11308 11796 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 13354 11336 13360 11348
rect 13315 11308 13360 11336
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16264 11308 16681 11336
rect 16264 11296 16270 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 17957 11339 18015 11345
rect 17957 11305 17969 11339
rect 18003 11336 18015 11339
rect 19978 11336 19984 11348
rect 18003 11308 19984 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 3528 11268 3556 11296
rect 5258 11268 5264 11280
rect 2792 11240 3556 11268
rect 3620 11240 5264 11268
rect 1443 11172 2728 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 3620 11200 3648 11240
rect 5258 11228 5264 11240
rect 5316 11228 5322 11280
rect 6448 11271 6506 11277
rect 6448 11237 6460 11271
rect 6494 11268 6506 11271
rect 6822 11268 6828 11280
rect 6494 11240 6828 11268
rect 6494 11237 6506 11240
rect 6448 11231 6506 11237
rect 6822 11228 6828 11240
rect 6880 11228 6886 11280
rect 8386 11228 8392 11280
rect 8444 11268 8450 11280
rect 9217 11271 9275 11277
rect 9217 11268 9229 11271
rect 8444 11240 9229 11268
rect 8444 11228 8450 11240
rect 9217 11237 9229 11240
rect 9263 11237 9275 11271
rect 9217 11231 9275 11237
rect 11140 11271 11198 11277
rect 11140 11237 11152 11271
rect 11186 11268 11198 11271
rect 11238 11268 11244 11280
rect 11186 11240 11244 11268
rect 11186 11237 11198 11240
rect 11140 11231 11198 11237
rect 11238 11228 11244 11240
rect 11296 11228 11302 11280
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 13262 11268 13268 11280
rect 11388 11240 13268 11268
rect 11388 11228 11394 11240
rect 13262 11228 13268 11240
rect 13320 11268 13326 11280
rect 13725 11271 13783 11277
rect 13725 11268 13737 11271
rect 13320 11240 13737 11268
rect 13320 11228 13326 11240
rect 13725 11237 13737 11240
rect 13771 11237 13783 11271
rect 16684 11268 16712 11299
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 18325 11271 18383 11277
rect 18325 11268 18337 11271
rect 16684 11240 18337 11268
rect 13725 11231 13783 11237
rect 18325 11237 18337 11240
rect 18371 11268 18383 11271
rect 18598 11268 18604 11280
rect 18371 11240 18604 11268
rect 18371 11237 18383 11240
rect 18325 11231 18383 11237
rect 18598 11228 18604 11240
rect 18656 11228 18662 11280
rect 2832 11172 3648 11200
rect 2832 11160 2838 11172
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 6178 11200 6184 11212
rect 4580 11172 4625 11200
rect 6139 11172 6184 11200
rect 4580 11160 4586 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 14642 11200 14648 11212
rect 14507 11172 14648 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 14642 11160 14648 11172
rect 14700 11200 14706 11212
rect 15556 11203 15614 11209
rect 15556 11200 15568 11203
rect 14700 11172 15568 11200
rect 14700 11160 14706 11172
rect 15556 11169 15568 11172
rect 15602 11200 15614 11203
rect 15838 11200 15844 11212
rect 15602 11172 15844 11200
rect 15602 11169 15614 11172
rect 15556 11163 15614 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 17770 11200 17776 11212
rect 17731 11172 17776 11200
rect 17770 11160 17776 11172
rect 17828 11160 17834 11212
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 3053 11095 3111 11101
rect 2317 11067 2375 11073
rect 2317 11033 2329 11067
rect 2363 11064 2375 11067
rect 2590 11064 2596 11076
rect 2363 11036 2596 11064
rect 2363 11033 2375 11036
rect 2317 11027 2375 11033
rect 2590 11024 2596 11036
rect 2648 11024 2654 11076
rect 3068 10996 3096 11095
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10560 11104 10885 11132
rect 10560 11092 10566 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 13817 11135 13875 11141
rect 13817 11132 13829 11135
rect 13780 11104 13829 11132
rect 13780 11092 13786 11104
rect 13817 11101 13829 11104
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 15286 11132 15292 11144
rect 13964 11104 14009 11132
rect 15247 11104 15292 11132
rect 13964 11092 13970 11104
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 4062 11064 4068 11076
rect 4023 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5534 11064 5540 11076
rect 5307 11036 5540 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 10413 11067 10471 11073
rect 10413 11033 10425 11067
rect 10459 11064 10471 11067
rect 10778 11064 10784 11076
rect 10459 11036 10784 11064
rect 10459 11033 10471 11036
rect 10413 11027 10471 11033
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 12897 11067 12955 11073
rect 12897 11033 12909 11067
rect 12943 11064 12955 11067
rect 13265 11067 13323 11073
rect 13265 11064 13277 11067
rect 12943 11036 13277 11064
rect 12943 11033 12955 11036
rect 12897 11027 12955 11033
rect 13265 11033 13277 11036
rect 13311 11064 13323 11067
rect 13538 11064 13544 11076
rect 13311 11036 13544 11064
rect 13311 11033 13323 11036
rect 13265 11027 13323 11033
rect 13538 11024 13544 11036
rect 13596 11064 13602 11076
rect 13924 11064 13952 11092
rect 13596 11036 13952 11064
rect 13596 11024 13602 11036
rect 3142 10996 3148 11008
rect 3068 10968 3148 10996
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 7558 10996 7564 11008
rect 7519 10968 7564 10996
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 12253 10999 12311 11005
rect 12253 10965 12265 10999
rect 12299 10996 12311 10999
rect 12434 10996 12440 11008
rect 12299 10968 12440 10996
rect 12299 10965 12311 10968
rect 12253 10959 12311 10965
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 17126 10956 17132 11008
rect 17184 10996 17190 11008
rect 17221 10999 17279 11005
rect 17221 10996 17233 10999
rect 17184 10968 17233 10996
rect 17184 10956 17190 10968
rect 17221 10965 17233 10968
rect 17267 10965 17279 10999
rect 17221 10959 17279 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3384 10764 3525 10792
rect 3384 10752 3390 10764
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 3513 10755 3571 10761
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6822 10792 6828 10804
rect 6687 10764 6828 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 8628 10764 8677 10792
rect 8628 10752 8634 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 10502 10792 10508 10804
rect 8665 10755 8723 10761
rect 9784 10764 10508 10792
rect 6196 10724 6224 10752
rect 7101 10727 7159 10733
rect 7101 10724 7113 10727
rect 6196 10696 7113 10724
rect 7101 10693 7113 10696
rect 7147 10724 7159 10727
rect 7147 10696 7328 10724
rect 7147 10693 7159 10696
rect 7101 10687 7159 10693
rect 7300 10665 7328 10696
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 1581 10591 1639 10597
rect 1581 10557 1593 10591
rect 1627 10588 1639 10591
rect 2958 10588 2964 10600
rect 1627 10560 2964 10588
rect 1627 10557 1639 10560
rect 1581 10551 1639 10557
rect 2958 10548 2964 10560
rect 3016 10588 3022 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3016 10560 3985 10588
rect 3016 10548 3022 10560
rect 3973 10557 3985 10560
rect 4019 10588 4031 10591
rect 4062 10588 4068 10600
rect 4019 10560 4068 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4062 10548 4068 10560
rect 4120 10588 4126 10600
rect 5166 10588 5172 10600
rect 4120 10560 5172 10588
rect 4120 10548 4126 10560
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 7300 10588 7328 10619
rect 9784 10597 9812 10764
rect 10502 10752 10508 10764
rect 10560 10792 10566 10804
rect 11149 10795 11207 10801
rect 10560 10764 10732 10792
rect 10560 10752 10566 10764
rect 10704 10724 10732 10764
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 11238 10792 11244 10804
rect 11195 10764 11244 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 13906 10792 13912 10804
rect 13863 10764 13912 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 15746 10792 15752 10804
rect 15243 10764 15752 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 15896 10764 16221 10792
rect 15896 10752 15902 10764
rect 16209 10761 16221 10764
rect 16255 10761 16267 10795
rect 16942 10792 16948 10804
rect 16903 10764 16948 10792
rect 16209 10755 16267 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 19242 10792 19248 10804
rect 18555 10764 19248 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 11701 10727 11759 10733
rect 11701 10724 11713 10727
rect 10704 10696 11713 10724
rect 11701 10693 11713 10696
rect 11747 10724 11759 10727
rect 12161 10727 12219 10733
rect 12161 10724 12173 10727
rect 11747 10696 12173 10724
rect 11747 10693 11759 10696
rect 11701 10687 11759 10693
rect 12161 10693 12173 10696
rect 12207 10693 12219 10727
rect 12161 10687 12219 10693
rect 15105 10727 15163 10733
rect 15105 10693 15117 10727
rect 15151 10724 15163 10727
rect 15286 10724 15292 10736
rect 15151 10696 15292 10724
rect 15151 10693 15163 10696
rect 15105 10687 15163 10693
rect 12176 10656 12204 10687
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 12176 10628 12449 10656
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 15746 10656 15752 10668
rect 15707 10628 15752 10656
rect 12437 10619 12495 10625
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 7300 10560 9689 10588
rect 9677 10557 9689 10560
rect 9723 10588 9735 10591
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9723 10560 9781 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10025 10591 10083 10597
rect 10025 10588 10037 10591
rect 9916 10560 10037 10588
rect 9916 10548 9922 10560
rect 10025 10557 10037 10560
rect 10071 10557 10083 10591
rect 10025 10551 10083 10557
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 16577 10591 16635 10597
rect 16577 10588 16589 10591
rect 15712 10560 16589 10588
rect 15712 10548 15718 10560
rect 16577 10557 16589 10560
rect 16623 10557 16635 10591
rect 16758 10588 16764 10600
rect 16719 10560 16764 10588
rect 16577 10551 16635 10557
rect 16758 10548 16764 10560
rect 16816 10588 16822 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 16816 10560 17233 10588
rect 16816 10548 16822 10560
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 17221 10551 17279 10557
rect 18230 10548 18236 10600
rect 18288 10588 18294 10600
rect 18325 10591 18383 10597
rect 18325 10588 18337 10591
rect 18288 10560 18337 10588
rect 18288 10548 18294 10560
rect 18325 10557 18337 10560
rect 18371 10588 18383 10591
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 18371 10560 18889 10588
rect 18371 10557 18383 10560
rect 18325 10551 18383 10557
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 1848 10523 1906 10529
rect 1848 10489 1860 10523
rect 1894 10520 1906 10523
rect 2038 10520 2044 10532
rect 1894 10492 2044 10520
rect 1894 10489 1906 10492
rect 1848 10483 1906 10489
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 2590 10480 2596 10532
rect 2648 10520 2654 10532
rect 4332 10523 4390 10529
rect 4332 10520 4344 10523
rect 2648 10492 4344 10520
rect 2648 10480 2654 10492
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 2406 10452 2412 10464
rect 2280 10424 2412 10452
rect 2280 10412 2286 10424
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 2976 10461 3004 10492
rect 4332 10489 4344 10492
rect 4378 10520 4390 10523
rect 4890 10520 4896 10532
rect 4378 10492 4896 10520
rect 4378 10489 4390 10492
rect 4332 10483 4390 10489
rect 4890 10480 4896 10492
rect 4948 10480 4954 10532
rect 7558 10529 7564 10532
rect 7552 10520 7564 10529
rect 7471 10492 7564 10520
rect 7552 10483 7564 10492
rect 7616 10520 7622 10532
rect 8662 10520 8668 10532
rect 7616 10492 8668 10520
rect 7558 10480 7564 10483
rect 7616 10480 7622 10492
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 9309 10523 9367 10529
rect 9309 10489 9321 10523
rect 9355 10520 9367 10523
rect 9490 10520 9496 10532
rect 9355 10492 9496 10520
rect 9355 10489 9367 10492
rect 9309 10483 9367 10489
rect 9490 10480 9496 10492
rect 9548 10520 9554 10532
rect 9876 10520 9904 10548
rect 9548 10492 9904 10520
rect 9548 10480 9554 10492
rect 12434 10480 12440 10532
rect 12492 10520 12498 10532
rect 12682 10523 12740 10529
rect 12682 10520 12694 10523
rect 12492 10492 12694 10520
rect 12492 10480 12498 10492
rect 12682 10489 12694 10492
rect 12728 10489 12740 10523
rect 12682 10483 12740 10489
rect 14737 10523 14795 10529
rect 14737 10489 14749 10523
rect 14783 10520 14795 10523
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 14783 10492 15577 10520
rect 14783 10489 14795 10492
rect 14737 10483 14795 10489
rect 15565 10489 15577 10492
rect 15611 10520 15623 10523
rect 16482 10520 16488 10532
rect 15611 10492 16488 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 16482 10480 16488 10492
rect 16540 10480 16546 10532
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 4028 10424 5457 10452
rect 4028 10412 4034 10424
rect 5445 10421 5457 10424
rect 5491 10421 5503 10455
rect 15654 10452 15660 10464
rect 15615 10424 15660 10452
rect 5445 10415 5503 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 2774 10248 2780 10260
rect 2700 10220 2780 10248
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10180 2375 10183
rect 2700 10180 2728 10220
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 3878 10248 3884 10260
rect 3839 10220 3884 10248
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 4614 10248 4620 10260
rect 4575 10220 4620 10248
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 4890 10248 4896 10260
rect 4851 10220 4896 10248
rect 4890 10208 4896 10220
rect 4948 10208 4954 10260
rect 8662 10248 8668 10260
rect 8623 10220 8668 10248
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9490 10248 9496 10260
rect 9451 10220 9496 10248
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10870 10248 10876 10260
rect 9723 10220 10876 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 10965 10251 11023 10257
rect 10965 10217 10977 10251
rect 11011 10248 11023 10251
rect 11238 10248 11244 10260
rect 11011 10220 11244 10248
rect 11011 10217 11023 10220
rect 10965 10211 11023 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13446 10248 13452 10260
rect 13407 10220 13452 10248
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13872 10220 13921 10248
rect 13872 10208 13878 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 17126 10248 17132 10260
rect 17087 10220 17132 10248
rect 13909 10211 13967 10217
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 17368 10220 18429 10248
rect 17368 10208 17374 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 18417 10211 18475 10217
rect 3510 10180 3516 10192
rect 2363 10152 2728 10180
rect 3423 10152 3516 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 3510 10140 3516 10152
rect 3568 10180 3574 10192
rect 3970 10180 3976 10192
rect 3568 10152 3976 10180
rect 3568 10140 3574 10152
rect 3970 10140 3976 10152
rect 4028 10140 4034 10192
rect 4632 10180 4660 10208
rect 5350 10180 5356 10192
rect 4632 10152 5356 10180
rect 5350 10140 5356 10152
rect 5408 10189 5414 10192
rect 5408 10183 5472 10189
rect 5408 10149 5426 10183
rect 5460 10149 5472 10183
rect 9508 10180 9536 10208
rect 9508 10152 10272 10180
rect 5408 10143 5472 10149
rect 5408 10140 5414 10143
rect 2774 10072 2780 10124
rect 2832 10112 2838 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 2832 10084 4077 10112
rect 2832 10072 2838 10084
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 5166 10112 5172 10124
rect 5079 10084 5172 10112
rect 4065 10075 4123 10081
rect 5166 10072 5172 10084
rect 5224 10112 5230 10124
rect 5994 10112 6000 10124
rect 5224 10084 6000 10112
rect 5224 10072 5230 10084
rect 5994 10072 6000 10084
rect 6052 10112 6058 10124
rect 6178 10112 6184 10124
rect 6052 10084 6184 10112
rect 6052 10072 6058 10084
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 7466 10072 7472 10124
rect 7524 10112 7530 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 7524 10084 7573 10112
rect 7524 10072 7530 10084
rect 7561 10081 7573 10084
rect 7607 10112 7619 10115
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7607 10084 8033 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 8021 10081 8033 10084
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9456 10084 10057 10112
rect 9456 10072 9462 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3142 10044 3148 10056
rect 3099 10016 3148 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3142 10004 3148 10016
rect 3200 10044 3206 10056
rect 3510 10044 3516 10056
rect 3200 10016 3516 10044
rect 3200 10004 3206 10016
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 8110 10044 8116 10056
rect 7239 10016 7972 10044
rect 8071 10016 8116 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7650 9976 7656 9988
rect 7611 9948 7656 9976
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 7944 9976 7972 10016
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 8205 10007 8263 10013
rect 8018 9976 8024 9988
rect 7931 9948 8024 9976
rect 8018 9936 8024 9948
rect 8076 9976 8082 9988
rect 8220 9976 8248 10007
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10244 10053 10272 10152
rect 15746 10140 15752 10192
rect 15804 10180 15810 10192
rect 15994 10183 16052 10189
rect 15994 10180 16006 10183
rect 15804 10152 16006 10180
rect 15804 10140 15810 10152
rect 15994 10149 16006 10152
rect 16040 10149 16052 10183
rect 15994 10143 16052 10149
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 13814 10112 13820 10124
rect 11756 10084 11801 10112
rect 13775 10084 13820 10112
rect 11756 10072 11762 10084
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18196 10084 18245 10112
rect 18196 10072 18202 10084
rect 18233 10081 18245 10084
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 10137 10047 10195 10053
rect 9732 10016 9996 10044
rect 9732 10004 9738 10016
rect 9968 9988 9996 10016
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 10229 10007 10287 10013
rect 8076 9948 8248 9976
rect 8076 9936 8082 9948
rect 9950 9936 9956 9988
rect 10008 9936 10014 9988
rect 10152 9976 10180 10007
rect 11790 10004 11796 10016
rect 11848 10044 11854 10056
rect 12434 10044 12440 10056
rect 11848 10016 12440 10044
rect 11848 10004 11854 10016
rect 12434 10004 12440 10016
rect 12492 10044 12498 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12492 10016 12817 10044
rect 12492 10004 12498 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 14090 10044 14096 10056
rect 14051 10016 14096 10044
rect 12805 10007 12863 10013
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 15286 10004 15292 10056
rect 15344 10044 15350 10056
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15344 10016 15761 10044
rect 15344 10004 15350 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 10410 9976 10416 9988
rect 10152 9948 10416 9976
rect 10410 9936 10416 9948
rect 10468 9936 10474 9988
rect 11241 9979 11299 9985
rect 11241 9945 11253 9979
rect 11287 9976 11299 9979
rect 13722 9976 13728 9988
rect 11287 9948 13728 9976
rect 11287 9945 11299 9948
rect 11241 9939 11299 9945
rect 13722 9936 13728 9948
rect 13780 9976 13786 9988
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 13780 9948 14473 9976
rect 13780 9936 13786 9948
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 14461 9939 14519 9945
rect 6546 9908 6552 9920
rect 6507 9880 6552 9908
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9582 9908 9588 9920
rect 9171 9880 9588 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10686 9908 10692 9920
rect 9732 9880 10692 9908
rect 9732 9868 9738 9880
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12986 9908 12992 9920
rect 12575 9880 12992 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 15565 9911 15623 9917
rect 15565 9877 15577 9911
rect 15611 9908 15623 9911
rect 15746 9908 15752 9920
rect 15611 9880 15752 9908
rect 15611 9877 15623 9880
rect 15565 9871 15623 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 3510 9704 3516 9716
rect 2832 9676 2877 9704
rect 3471 9676 3516 9704
rect 2832 9664 2838 9676
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 5350 9704 5356 9716
rect 5311 9676 5356 9704
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 9582 9704 9588 9716
rect 8220 9676 9588 9704
rect 1397 9639 1455 9645
rect 1397 9605 1409 9639
rect 1443 9636 1455 9639
rect 2130 9636 2136 9648
rect 1443 9608 2136 9636
rect 1443 9605 1455 9608
rect 1397 9599 1455 9605
rect 2130 9596 2136 9608
rect 2188 9596 2194 9648
rect 2406 9636 2412 9648
rect 2367 9608 2412 9636
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 3145 9639 3203 9645
rect 3145 9636 3157 9639
rect 2556 9608 3157 9636
rect 2556 9596 2562 9608
rect 3145 9605 3157 9608
rect 3191 9605 3203 9639
rect 3145 9599 3203 9605
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 3528 9568 3556 9664
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 5368 9636 5396 9664
rect 6273 9639 6331 9645
rect 6273 9636 6285 9639
rect 5368 9608 6285 9636
rect 6273 9605 6285 9608
rect 6319 9605 6331 9639
rect 7558 9636 7564 9648
rect 7519 9608 7564 9636
rect 6273 9599 6331 9605
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 8021 9639 8079 9645
rect 8021 9605 8033 9639
rect 8067 9636 8079 9639
rect 8220 9636 8248 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 10410 9704 10416 9716
rect 9692 9676 10416 9704
rect 9033 9639 9091 9645
rect 9033 9636 9045 9639
rect 8067 9608 8248 9636
rect 8496 9608 9045 9636
rect 8067 9605 8079 9608
rect 8021 9599 8079 9605
rect 5000 9568 5028 9596
rect 5442 9568 5448 9580
rect 3528 9540 4108 9568
rect 5000 9540 5448 9568
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 1452 9472 1777 9500
rect 1452 9460 1458 9472
rect 1765 9469 1777 9472
rect 1811 9500 1823 9503
rect 1854 9500 1860 9512
rect 1811 9472 1860 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 3970 9500 3976 9512
rect 3927 9472 3976 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4080 9500 4108 9540
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 5592 9540 6837 9568
rect 5592 9528 5598 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 7576 9568 7604 9596
rect 8496 9577 8524 9608
rect 9033 9605 9045 9608
rect 9079 9636 9091 9639
rect 9692 9636 9720 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 11238 9704 11244 9716
rect 11151 9676 11244 9704
rect 11238 9664 11244 9676
rect 11296 9704 11302 9716
rect 11698 9704 11704 9716
rect 11296 9676 11704 9704
rect 11296 9664 11302 9676
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 12066 9664 12072 9716
rect 12124 9704 12130 9716
rect 12250 9704 12256 9716
rect 12124 9676 12256 9704
rect 12124 9664 12130 9676
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 13906 9704 13912 9716
rect 13867 9676 13912 9704
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 14277 9707 14335 9713
rect 14277 9673 14289 9707
rect 14323 9704 14335 9707
rect 15286 9704 15292 9716
rect 14323 9676 15292 9704
rect 14323 9673 14335 9676
rect 14277 9667 14335 9673
rect 15286 9664 15292 9676
rect 15344 9704 15350 9716
rect 16301 9707 16359 9713
rect 16301 9704 16313 9707
rect 15344 9676 16313 9704
rect 15344 9664 15350 9676
rect 16301 9673 16313 9676
rect 16347 9673 16359 9707
rect 18230 9704 18236 9716
rect 18191 9676 18236 9704
rect 16301 9667 16359 9673
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 9079 9608 9720 9636
rect 9079 9605 9091 9608
rect 9033 9599 9091 9605
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 12216 9608 14412 9636
rect 12216 9596 12222 9608
rect 8481 9571 8539 9577
rect 8481 9568 8493 9571
rect 7576 9540 8493 9568
rect 6825 9531 6883 9537
rect 8481 9537 8493 9540
rect 8527 9537 8539 9571
rect 8662 9568 8668 9580
rect 8623 9540 8668 9568
rect 8481 9531 8539 9537
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 9640 9540 10057 9568
rect 9640 9528 9646 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10686 9568 10692 9580
rect 10275 9540 10692 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 14384 9577 14412 9608
rect 18138 9596 18144 9648
rect 18196 9636 18202 9648
rect 18509 9639 18567 9645
rect 18509 9636 18521 9639
rect 18196 9608 18521 9636
rect 18196 9596 18202 9608
rect 18509 9605 18521 9608
rect 18555 9605 18567 9639
rect 18509 9599 18567 9605
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16632 9540 16865 9568
rect 16632 9528 16638 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 4246 9509 4252 9512
rect 4229 9503 4252 9509
rect 4229 9500 4241 9503
rect 4080 9472 4241 9500
rect 4229 9469 4241 9472
rect 4304 9500 4310 9512
rect 18046 9500 18052 9512
rect 4304 9472 4377 9500
rect 18007 9472 18052 9500
rect 4229 9463 4252 9469
rect 4246 9460 4252 9463
rect 4304 9460 4310 9472
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 18104 9472 18889 9500
rect 18104 9460 18110 9472
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 11379 9404 12173 9432
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 12161 9401 12173 9404
rect 12207 9432 12219 9435
rect 12805 9435 12863 9441
rect 12805 9432 12817 9435
rect 12207 9404 12817 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12805 9401 12817 9404
rect 12851 9401 12863 9435
rect 12805 9395 12863 9401
rect 14090 9392 14096 9444
rect 14148 9432 14154 9444
rect 14614 9435 14672 9441
rect 14614 9432 14626 9435
rect 14148 9404 14626 9432
rect 14148 9392 14154 9404
rect 14614 9401 14626 9404
rect 14660 9401 14672 9435
rect 14614 9395 14672 9401
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 1820 9336 1869 9364
rect 1820 9324 1826 9336
rect 1857 9333 1869 9336
rect 1903 9333 1915 9367
rect 5994 9364 6000 9376
rect 5907 9336 6000 9364
rect 1857 9327 1915 9333
rect 5994 9324 6000 9336
rect 6052 9364 6058 9376
rect 6638 9364 6644 9376
rect 6052 9336 6644 9364
rect 6052 9324 6058 9336
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7834 9364 7840 9376
rect 7795 9336 7840 9364
rect 7834 9324 7840 9336
rect 7892 9364 7898 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 7892 9336 8401 9364
rect 7892 9324 7898 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 9398 9364 9404 9376
rect 9359 9336 9404 9364
rect 8389 9327 8447 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9732 9336 9965 9364
rect 9732 9324 9738 9336
rect 9953 9333 9965 9336
rect 9999 9364 10011 9367
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 9999 9336 10609 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10597 9333 10609 9336
rect 10643 9333 10655 9367
rect 10597 9327 10655 9333
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11664 9336 11805 9364
rect 11664 9324 11670 9336
rect 11793 9333 11805 9336
rect 11839 9333 11851 9367
rect 11793 9327 11851 9333
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12894 9364 12900 9376
rect 12492 9336 12537 9364
rect 12855 9336 12900 9364
rect 12492 9324 12498 9336
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9364 13510 9376
rect 13722 9364 13728 9376
rect 13504 9336 13728 9364
rect 13504 9324 13510 9336
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 15746 9364 15752 9376
rect 15707 9336 15752 9364
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 1670 9160 1676 9172
rect 1627 9132 1676 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1912 9132 1961 9160
rect 1912 9120 1918 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 1949 9123 2007 9129
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2096 9132 2329 9160
rect 2096 9120 2102 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2317 9123 2375 9129
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 4062 9160 4068 9172
rect 3927 9132 4068 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4246 9160 4252 9172
rect 4207 9132 4252 9160
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 4580 9132 4629 9160
rect 4580 9120 4586 9132
rect 4617 9129 4629 9132
rect 4663 9129 4675 9163
rect 4617 9123 4675 9129
rect 5442 9120 5448 9172
rect 5500 9160 5506 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 5500 9132 5549 9160
rect 5500 9120 5506 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 8018 9160 8024 9172
rect 7979 9132 8024 9160
rect 5537 9123 5595 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 11790 9160 11796 9172
rect 11747 9132 11796 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 11885 9163 11943 9169
rect 11885 9129 11897 9163
rect 11931 9160 11943 9163
rect 12894 9160 12900 9172
rect 11931 9132 12900 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13044 9132 13553 9160
rect 13044 9120 13050 9132
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 14090 9160 14096 9172
rect 14051 9132 14096 9160
rect 13541 9123 13599 9129
rect 14090 9120 14096 9132
rect 14148 9160 14154 9172
rect 14461 9163 14519 9169
rect 14461 9160 14473 9163
rect 14148 9132 14473 9160
rect 14148 9120 14154 9132
rect 14461 9129 14473 9132
rect 14507 9129 14519 9163
rect 15746 9160 15752 9172
rect 15707 9132 15752 9160
rect 14461 9123 14519 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 16761 9163 16819 9169
rect 16761 9129 16773 9163
rect 16807 9160 16819 9163
rect 17770 9160 17776 9172
rect 16807 9132 17776 9160
rect 16807 9129 16819 9132
rect 16761 9123 16819 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 2682 9052 2688 9104
rect 2740 9092 2746 9104
rect 3329 9095 3387 9101
rect 3329 9092 3341 9095
rect 2740 9064 3341 9092
rect 2740 9052 2746 9064
rect 3329 9061 3341 9064
rect 3375 9061 3387 9095
rect 3329 9055 3387 9061
rect 6546 9052 6552 9104
rect 6604 9092 6610 9104
rect 6886 9095 6944 9101
rect 6886 9092 6898 9095
rect 6604 9064 6898 9092
rect 6604 9052 6610 9064
rect 6886 9061 6898 9064
rect 6932 9061 6944 9095
rect 8662 9092 8668 9104
rect 8575 9064 8668 9092
rect 6886 9055 6944 9061
rect 8662 9052 8668 9064
rect 8720 9092 8726 9104
rect 9858 9092 9864 9104
rect 8720 9064 9864 9092
rect 8720 9052 8726 9064
rect 9858 9052 9864 9064
rect 9916 9101 9922 9104
rect 9916 9095 9980 9101
rect 9916 9061 9934 9095
rect 9968 9061 9980 9095
rect 9916 9055 9980 9061
rect 15289 9095 15347 9101
rect 15289 9061 15301 9095
rect 15335 9092 15347 9095
rect 16390 9092 16396 9104
rect 15335 9064 16396 9092
rect 15335 9061 15347 9064
rect 15289 9055 15347 9061
rect 9916 9052 9922 9055
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 2590 9024 2596 9036
rect 2547 8996 2596 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 5350 8984 5356 9036
rect 5408 9024 5414 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 5408 8996 5457 9024
rect 5408 8984 5414 8996
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 6564 9024 6592 9052
rect 5445 8987 5503 8993
rect 5736 8996 6592 9024
rect 5736 8965 5764 8996
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 7374 9024 7380 9036
rect 6696 8996 7380 9024
rect 6696 8984 6702 8996
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 10226 9024 10232 9036
rect 9723 8996 10232 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 12417 9027 12475 9033
rect 12417 9024 12429 9027
rect 11940 8996 12429 9024
rect 11940 8984 11946 8996
rect 12417 8993 12429 8996
rect 12463 8993 12475 9027
rect 16574 9024 16580 9036
rect 16535 8996 16580 9024
rect 12417 8987 12475 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 8938 8956 8944 8968
rect 8899 8928 8944 8956
rect 5721 8919 5779 8925
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 12158 8956 12164 8968
rect 12119 8928 12164 8956
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 2682 8888 2688 8900
rect 2643 8860 2688 8888
rect 2682 8848 2688 8860
rect 2740 8848 2746 8900
rect 5074 8888 5080 8900
rect 5035 8860 5080 8888
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 10686 8820 10692 8832
rect 9539 8792 10692 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 10686 8780 10692 8792
rect 10744 8820 10750 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10744 8792 11069 8820
rect 10744 8780 10750 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11756 8792 11897 8820
rect 11756 8780 11762 8792
rect 11885 8789 11897 8792
rect 11931 8820 11943 8823
rect 11977 8823 12035 8829
rect 11977 8820 11989 8823
rect 11931 8792 11989 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 11977 8789 11989 8792
rect 12023 8789 12035 8823
rect 11977 8783 12035 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 2314 8616 2320 8628
rect 1995 8588 2320 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1964 8412 1992 8579
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 5442 8616 5448 8628
rect 5403 8588 5448 8616
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5905 8619 5963 8625
rect 5905 8585 5917 8619
rect 5951 8616 5963 8619
rect 6546 8616 6552 8628
rect 5951 8588 6552 8616
rect 5951 8585 5963 8588
rect 5905 8579 5963 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 10100 8588 10241 8616
rect 10100 8576 10106 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 11698 8616 11704 8628
rect 10827 8588 11704 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 5350 8548 5356 8560
rect 5215 8520 5356 8548
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 9858 8548 9864 8560
rect 9355 8520 9864 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10244 8548 10272 8579
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 11882 8616 11888 8628
rect 11843 8588 11888 8616
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12713 8619 12771 8625
rect 12713 8616 12725 8619
rect 12216 8588 12725 8616
rect 12216 8576 12222 8588
rect 12713 8585 12725 8588
rect 12759 8585 12771 8619
rect 12713 8579 12771 8585
rect 10244 8520 11284 8548
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7466 8480 7472 8492
rect 6963 8452 7472 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 10594 8480 10600 8492
rect 10555 8452 10600 8480
rect 10594 8440 10600 8452
rect 10652 8480 10658 8492
rect 11256 8489 11284 8520
rect 11241 8483 11299 8489
rect 10652 8452 11192 8480
rect 10652 8440 10658 8452
rect 2590 8412 2596 8424
rect 1443 8384 1992 8412
rect 2551 8384 2596 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7760 8384 7941 8412
rect 7760 8344 7788 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 8018 8372 8024 8424
rect 8076 8412 8082 8424
rect 11164 8421 11192 8452
rect 11241 8449 11253 8483
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 11425 8483 11483 8489
rect 11425 8449 11437 8483
rect 11471 8480 11483 8483
rect 11882 8480 11888 8492
rect 11471 8452 11888 8480
rect 11471 8449 11483 8452
rect 11425 8443 11483 8449
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 12728 8480 12756 8579
rect 14090 8576 14096 8628
rect 14148 8616 14154 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 14148 8588 14289 8616
rect 14148 8576 14154 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 16574 8616 16580 8628
rect 16535 8588 16580 8616
rect 14277 8579 14335 8585
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12728 8452 12909 8480
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 8185 8415 8243 8421
rect 8185 8412 8197 8415
rect 8076 8384 8197 8412
rect 8076 8372 8082 8384
rect 8185 8381 8197 8384
rect 8231 8381 8243 8415
rect 8185 8375 8243 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13153 8415 13211 8421
rect 13153 8412 13165 8415
rect 13044 8384 13165 8412
rect 13044 8372 13050 8384
rect 13153 8381 13165 8384
rect 13199 8381 13211 8415
rect 13153 8375 13211 8381
rect 9861 8347 9919 8353
rect 9861 8344 9873 8347
rect 7760 8316 9873 8344
rect 7466 8276 7472 8288
rect 7427 8248 7472 8276
rect 7466 8236 7472 8248
rect 7524 8276 7530 8288
rect 7760 8285 7788 8316
rect 9861 8313 9873 8316
rect 9907 8344 9919 8347
rect 10226 8344 10232 8356
rect 9907 8316 10232 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 10226 8304 10232 8316
rect 10284 8344 10290 8356
rect 12158 8344 12164 8356
rect 10284 8316 12164 8344
rect 10284 8304 10290 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 7524 8248 7757 8276
rect 7524 8236 7530 8248
rect 7745 8245 7757 8248
rect 7791 8245 7803 8279
rect 7745 8239 7803 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 8032 1400 8084
rect 1452 8032 1458 8084
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1544 8044 1593 8072
rect 1544 8032 1550 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 8018 8072 8024 8084
rect 7979 8044 8024 8072
rect 2225 8035 2283 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 9858 8072 9864 8084
rect 9819 8044 9864 8072
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 11882 8072 11888 8084
rect 11747 8044 11888 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 11882 8032 11888 8044
rect 11940 8072 11946 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 11940 8044 12265 8072
rect 11940 8032 11946 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12986 8072 12992 8084
rect 12947 8044 12992 8072
rect 12253 8035 12311 8041
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 1412 8004 1440 8032
rect 1857 8007 1915 8013
rect 1857 8004 1869 8007
rect 1412 7976 1869 8004
rect 1857 7973 1869 7976
rect 1903 7973 1915 8007
rect 1857 7967 1915 7973
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1670 7936 1676 7948
rect 1443 7908 1676 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1670 7896 1676 7908
rect 1728 7936 1734 7948
rect 2222 7936 2228 7948
rect 1728 7908 2228 7936
rect 1728 7896 1734 7908
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 10594 7945 10600 7948
rect 10321 7939 10379 7945
rect 10321 7936 10333 7939
rect 10192 7908 10333 7936
rect 10192 7896 10198 7908
rect 10321 7905 10333 7908
rect 10367 7905 10379 7939
rect 10588 7936 10600 7945
rect 10555 7908 10600 7936
rect 10321 7899 10379 7905
rect 10588 7899 10600 7908
rect 10594 7896 10600 7899
rect 10652 7896 10658 7948
rect 566 7760 572 7812
rect 624 7800 630 7812
rect 9398 7800 9404 7812
rect 624 7772 9404 7800
rect 624 7760 630 7772
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1670 7528 1676 7540
rect 1631 7500 1676 7528
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10192 7500 10333 7528
rect 10192 7488 10198 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 10594 7488 10600 7540
rect 10652 7528 10658 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 10652 7500 10701 7528
rect 10652 7488 10658 7500
rect 10689 7497 10701 7500
rect 10735 7497 10747 7531
rect 10689 7491 10747 7497
rect 9674 7392 9680 7404
rect 9635 7364 9680 7392
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 10778 5352 10784 5364
rect 10643 5324 10784 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 9214 5148 9220 5160
rect 9175 5120 9220 5148
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9490 5089 9496 5092
rect 9125 5083 9183 5089
rect 9125 5049 9137 5083
rect 9171 5080 9183 5083
rect 9484 5080 9496 5089
rect 9171 5052 9496 5080
rect 9171 5049 9183 5052
rect 9125 5043 9183 5049
rect 9484 5043 9496 5052
rect 9490 5040 9496 5043
rect 9548 5040 9554 5092
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 7466 4468 7472 4480
rect 4672 4440 7472 4468
rect 4672 4428 4678 4440
rect 7466 4428 7472 4440
rect 7524 4468 7530 4480
rect 9214 4468 9220 4480
rect 7524 4440 9220 4468
rect 7524 4428 7530 4440
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 2136 25372 2188 25424
rect 2780 25372 2832 25424
rect 3424 25372 3476 25424
rect 1768 25304 1820 25356
rect 2320 25304 2372 25356
rect 3056 25347 3108 25356
rect 3056 25313 3065 25347
rect 3065 25313 3099 25347
rect 3099 25313 3108 25347
rect 3056 25304 3108 25313
rect 4712 25279 4764 25288
rect 4712 25245 4721 25279
rect 4721 25245 4755 25279
rect 4755 25245 4764 25279
rect 4712 25236 4764 25245
rect 1400 25168 1452 25220
rect 2596 25168 2648 25220
rect 4620 25168 4672 25220
rect 5080 25236 5132 25288
rect 6920 25279 6972 25288
rect 6920 25245 6929 25279
rect 6929 25245 6963 25279
rect 6963 25245 6972 25279
rect 6920 25236 6972 25245
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 2412 25143 2464 25152
rect 2412 25109 2421 25143
rect 2421 25109 2455 25143
rect 2455 25109 2464 25143
rect 2412 25100 2464 25109
rect 2780 25100 2832 25152
rect 6092 25100 6144 25152
rect 7840 25143 7892 25152
rect 7840 25109 7849 25143
rect 7849 25109 7883 25143
rect 7883 25109 7892 25143
rect 7840 25100 7892 25109
rect 13084 25100 13136 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1768 24896 1820 24948
rect 5080 24939 5132 24948
rect 2320 24871 2372 24880
rect 2320 24837 2329 24871
rect 2329 24837 2363 24871
rect 2363 24837 2372 24871
rect 2320 24828 2372 24837
rect 5080 24905 5089 24939
rect 5089 24905 5123 24939
rect 5123 24905 5132 24939
rect 5080 24896 5132 24905
rect 5356 24896 5408 24948
rect 2412 24760 2464 24812
rect 6184 24803 6236 24812
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 2504 24692 2556 24744
rect 2872 24692 2924 24744
rect 3516 24735 3568 24744
rect 3516 24701 3525 24735
rect 3525 24701 3559 24735
rect 3559 24701 3568 24735
rect 3516 24692 3568 24701
rect 4988 24692 5040 24744
rect 6184 24769 6193 24803
rect 6193 24769 6227 24803
rect 6227 24769 6236 24803
rect 6184 24760 6236 24769
rect 7380 24760 7432 24812
rect 12256 24803 12308 24812
rect 12256 24769 12265 24803
rect 12265 24769 12299 24803
rect 12299 24769 12308 24803
rect 12256 24760 12308 24769
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 9772 24692 9824 24744
rect 1768 24624 1820 24676
rect 8208 24667 8260 24676
rect 8208 24633 8217 24667
rect 8217 24633 8251 24667
rect 8251 24633 8260 24667
rect 8208 24624 8260 24633
rect 10048 24624 10100 24676
rect 2320 24556 2372 24608
rect 2504 24556 2556 24608
rect 3056 24556 3108 24608
rect 3976 24599 4028 24608
rect 3976 24565 3985 24599
rect 3985 24565 4019 24599
rect 4019 24565 4028 24599
rect 3976 24556 4028 24565
rect 4436 24599 4488 24608
rect 4436 24565 4445 24599
rect 4445 24565 4479 24599
rect 4479 24565 4488 24599
rect 4436 24556 4488 24565
rect 5540 24556 5592 24608
rect 7380 24556 7432 24608
rect 7748 24599 7800 24608
rect 7748 24565 7757 24599
rect 7757 24565 7791 24599
rect 7791 24565 7800 24599
rect 7748 24556 7800 24565
rect 7840 24556 7892 24608
rect 11152 24556 11204 24608
rect 11796 24599 11848 24608
rect 11796 24565 11805 24599
rect 11805 24565 11839 24599
rect 11839 24565 11848 24599
rect 11796 24556 11848 24565
rect 12624 24556 12676 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 2504 24395 2556 24404
rect 2504 24361 2513 24395
rect 2513 24361 2547 24395
rect 2547 24361 2556 24395
rect 2504 24352 2556 24361
rect 3976 24352 4028 24404
rect 7748 24352 7800 24404
rect 9680 24352 9732 24404
rect 11060 24352 11112 24404
rect 15660 24395 15712 24404
rect 15660 24361 15669 24395
rect 15669 24361 15703 24395
rect 15703 24361 15712 24395
rect 15660 24352 15712 24361
rect 17316 24395 17368 24404
rect 17316 24361 17325 24395
rect 17325 24361 17359 24395
rect 17359 24361 17368 24395
rect 17316 24352 17368 24361
rect 21824 24395 21876 24404
rect 21824 24361 21833 24395
rect 21833 24361 21867 24395
rect 21867 24361 21876 24395
rect 21824 24352 21876 24361
rect 22928 24395 22980 24404
rect 22928 24361 22937 24395
rect 22937 24361 22971 24395
rect 22971 24361 22980 24395
rect 22928 24352 22980 24361
rect 24032 24395 24084 24404
rect 24032 24361 24041 24395
rect 24041 24361 24075 24395
rect 24075 24361 24084 24395
rect 24032 24352 24084 24361
rect 2872 24284 2924 24336
rect 3792 24284 3844 24336
rect 4712 24284 4764 24336
rect 3056 24216 3108 24268
rect 8116 24284 8168 24336
rect 9772 24284 9824 24336
rect 4988 24259 5040 24268
rect 4988 24225 5022 24259
rect 5022 24225 5040 24259
rect 4988 24216 5040 24225
rect 6552 24216 6604 24268
rect 9220 24216 9272 24268
rect 11336 24259 11388 24268
rect 11336 24225 11345 24259
rect 11345 24225 11379 24259
rect 11379 24225 11388 24259
rect 11336 24216 11388 24225
rect 11612 24259 11664 24268
rect 11612 24225 11646 24259
rect 11646 24225 11664 24259
rect 11612 24216 11664 24225
rect 15476 24259 15528 24268
rect 15476 24225 15485 24259
rect 15485 24225 15519 24259
rect 15519 24225 15528 24259
rect 15476 24216 15528 24225
rect 17316 24216 17368 24268
rect 21548 24216 21600 24268
rect 22744 24259 22796 24268
rect 22744 24225 22753 24259
rect 22753 24225 22787 24259
rect 22787 24225 22796 24259
rect 22744 24216 22796 24225
rect 23848 24259 23900 24268
rect 23848 24225 23857 24259
rect 23857 24225 23891 24259
rect 23891 24225 23900 24259
rect 23848 24216 23900 24225
rect 2872 24148 2924 24200
rect 4436 24148 4488 24200
rect 7380 24123 7432 24132
rect 7380 24089 7389 24123
rect 7389 24089 7423 24123
rect 7423 24089 7432 24123
rect 9956 24148 10008 24200
rect 7380 24080 7432 24089
rect 2228 24012 2280 24064
rect 4620 24012 4672 24064
rect 7472 24055 7524 24064
rect 7472 24021 7481 24055
rect 7481 24021 7515 24055
rect 7515 24021 7524 24055
rect 7472 24012 7524 24021
rect 10140 24012 10192 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2412 23808 2464 23860
rect 3884 23808 3936 23860
rect 4712 23808 4764 23860
rect 8116 23851 8168 23860
rect 8116 23817 8125 23851
rect 8125 23817 8159 23851
rect 8159 23817 8168 23851
rect 8116 23808 8168 23817
rect 9220 23851 9272 23860
rect 9220 23817 9229 23851
rect 9229 23817 9263 23851
rect 9263 23817 9272 23851
rect 9220 23808 9272 23817
rect 9680 23851 9732 23860
rect 9680 23817 9689 23851
rect 9689 23817 9723 23851
rect 9723 23817 9732 23851
rect 9680 23808 9732 23817
rect 10048 23808 10100 23860
rect 11336 23808 11388 23860
rect 11704 23851 11756 23860
rect 11704 23817 11713 23851
rect 11713 23817 11747 23851
rect 11747 23817 11756 23851
rect 11704 23808 11756 23817
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 18604 23851 18656 23860
rect 18604 23817 18613 23851
rect 18613 23817 18647 23851
rect 18647 23817 18656 23851
rect 18604 23808 18656 23817
rect 21364 23808 21416 23860
rect 21916 23851 21968 23860
rect 21916 23817 21925 23851
rect 21925 23817 21959 23851
rect 21959 23817 21968 23851
rect 21916 23808 21968 23817
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 21824 23740 21876 23792
rect 25320 23740 25372 23792
rect 5356 23715 5408 23724
rect 5356 23681 5365 23715
rect 5365 23681 5399 23715
rect 5399 23681 5408 23715
rect 5356 23672 5408 23681
rect 5448 23715 5500 23724
rect 5448 23681 5457 23715
rect 5457 23681 5491 23715
rect 5491 23681 5500 23715
rect 5448 23672 5500 23681
rect 7012 23672 7064 23724
rect 5264 23647 5316 23656
rect 5264 23613 5273 23647
rect 5273 23613 5307 23647
rect 5307 23613 5316 23647
rect 5264 23604 5316 23613
rect 6828 23604 6880 23656
rect 7472 23647 7524 23656
rect 7472 23613 7481 23647
rect 7481 23613 7515 23647
rect 7515 23613 7524 23647
rect 7472 23604 7524 23613
rect 7748 23604 7800 23656
rect 9496 23604 9548 23656
rect 9772 23647 9824 23656
rect 9772 23613 9781 23647
rect 9781 23613 9815 23647
rect 9815 23613 9824 23647
rect 9772 23604 9824 23613
rect 2412 23579 2464 23588
rect 2412 23545 2446 23579
rect 2446 23545 2464 23579
rect 2412 23536 2464 23545
rect 2964 23536 3016 23588
rect 2688 23468 2740 23520
rect 2872 23468 2924 23520
rect 4436 23468 4488 23520
rect 6644 23536 6696 23588
rect 9956 23536 10008 23588
rect 11060 23536 11112 23588
rect 11612 23536 11664 23588
rect 12348 23536 12400 23588
rect 18420 23647 18472 23656
rect 13820 23536 13872 23588
rect 6552 23511 6604 23520
rect 6552 23477 6561 23511
rect 6561 23477 6595 23511
rect 6595 23477 6604 23511
rect 6552 23468 6604 23477
rect 6736 23468 6788 23520
rect 9680 23468 9732 23520
rect 12716 23511 12768 23520
rect 12716 23477 12725 23511
rect 12725 23477 12759 23511
rect 12759 23477 12768 23511
rect 12716 23468 12768 23477
rect 13544 23511 13596 23520
rect 13544 23477 13553 23511
rect 13553 23477 13587 23511
rect 13587 23477 13596 23511
rect 13544 23468 13596 23477
rect 15108 23511 15160 23520
rect 15108 23477 15117 23511
rect 15117 23477 15151 23511
rect 15151 23477 15160 23511
rect 15108 23468 15160 23477
rect 15476 23468 15528 23520
rect 18420 23613 18429 23647
rect 18429 23613 18463 23647
rect 18463 23613 18472 23647
rect 18420 23604 18472 23613
rect 19340 23604 19392 23656
rect 19248 23536 19300 23588
rect 21180 23604 21232 23656
rect 23480 23604 23532 23656
rect 23848 23604 23900 23656
rect 24768 23647 24820 23656
rect 24768 23613 24777 23647
rect 24777 23613 24811 23647
rect 24811 23613 24820 23647
rect 24768 23604 24820 23613
rect 16948 23468 17000 23520
rect 17316 23468 17368 23520
rect 21548 23511 21600 23520
rect 21548 23477 21557 23511
rect 21557 23477 21591 23511
rect 21591 23477 21600 23511
rect 21548 23468 21600 23477
rect 22744 23511 22796 23520
rect 22744 23477 22753 23511
rect 22753 23477 22787 23511
rect 22787 23477 22796 23511
rect 22744 23468 22796 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2136 23196 2188 23248
rect 2504 23196 2556 23248
rect 2872 23264 2924 23316
rect 4988 23264 5040 23316
rect 6828 23264 6880 23316
rect 7012 23307 7064 23316
rect 7012 23273 7021 23307
rect 7021 23273 7055 23307
rect 7055 23273 7064 23307
rect 7012 23264 7064 23273
rect 9496 23307 9548 23316
rect 9496 23273 9505 23307
rect 9505 23273 9539 23307
rect 9539 23273 9548 23307
rect 9496 23264 9548 23273
rect 12440 23264 12492 23316
rect 16488 23264 16540 23316
rect 16764 23307 16816 23316
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 16764 23264 16816 23273
rect 19340 23264 19392 23316
rect 21548 23264 21600 23316
rect 22376 23307 22428 23316
rect 22376 23273 22385 23307
rect 22385 23273 22419 23307
rect 22419 23273 22428 23307
rect 22376 23264 22428 23273
rect 23848 23264 23900 23316
rect 9772 23196 9824 23248
rect 10140 23239 10192 23248
rect 10140 23205 10149 23239
rect 10149 23205 10183 23239
rect 10183 23205 10192 23239
rect 10140 23196 10192 23205
rect 12072 23239 12124 23248
rect 12072 23205 12106 23239
rect 12106 23205 12124 23239
rect 12072 23196 12124 23205
rect 3056 23128 3108 23180
rect 3424 23128 3476 23180
rect 4436 23128 4488 23180
rect 4712 23128 4764 23180
rect 6644 23128 6696 23180
rect 7104 23171 7156 23180
rect 7104 23137 7113 23171
rect 7113 23137 7147 23171
rect 7147 23137 7156 23171
rect 7104 23128 7156 23137
rect 7380 23171 7432 23180
rect 7380 23137 7414 23171
rect 7414 23137 7432 23171
rect 7380 23128 7432 23137
rect 9680 23128 9732 23180
rect 11704 23128 11756 23180
rect 15568 23128 15620 23180
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 17868 23171 17920 23180
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 18880 23171 18932 23180
rect 18880 23137 18889 23171
rect 18889 23137 18923 23171
rect 18923 23137 18932 23171
rect 18880 23128 18932 23137
rect 20720 23128 20772 23180
rect 22192 23171 22244 23180
rect 22192 23137 22201 23171
rect 22201 23137 22235 23171
rect 22235 23137 22244 23171
rect 22192 23128 22244 23137
rect 23296 23171 23348 23180
rect 23296 23137 23305 23171
rect 23305 23137 23339 23171
rect 23339 23137 23348 23171
rect 23296 23128 23348 23137
rect 10140 23060 10192 23112
rect 1676 22924 1728 22976
rect 2872 22992 2924 23044
rect 19248 22992 19300 23044
rect 2136 22924 2188 22976
rect 6276 22924 6328 22976
rect 10048 22924 10100 22976
rect 10784 22967 10836 22976
rect 10784 22933 10793 22967
rect 10793 22933 10827 22967
rect 10827 22933 10836 22967
rect 10784 22924 10836 22933
rect 13820 22967 13872 22976
rect 13820 22933 13829 22967
rect 13829 22933 13863 22967
rect 13863 22933 13872 22967
rect 13820 22924 13872 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2504 22720 2556 22772
rect 7104 22763 7156 22772
rect 1492 22380 1544 22432
rect 7104 22729 7113 22763
rect 7113 22729 7147 22763
rect 7147 22729 7156 22763
rect 7104 22720 7156 22729
rect 8024 22720 8076 22772
rect 9680 22763 9732 22772
rect 9680 22729 9689 22763
rect 9689 22729 9723 22763
rect 9723 22729 9732 22763
rect 9680 22720 9732 22729
rect 10140 22720 10192 22772
rect 11704 22720 11756 22772
rect 11980 22720 12032 22772
rect 12072 22720 12124 22772
rect 13820 22720 13872 22772
rect 16304 22763 16356 22772
rect 16304 22729 16313 22763
rect 16313 22729 16347 22763
rect 16347 22729 16356 22763
rect 16304 22720 16356 22729
rect 16580 22720 16632 22772
rect 16764 22720 16816 22772
rect 6276 22584 6328 22636
rect 7380 22584 7432 22636
rect 6552 22516 6604 22568
rect 8208 22516 8260 22568
rect 1676 22448 1728 22500
rect 2688 22448 2740 22500
rect 6000 22448 6052 22500
rect 7012 22448 7064 22500
rect 7564 22448 7616 22500
rect 10784 22584 10836 22636
rect 10692 22516 10744 22568
rect 11060 22584 11112 22636
rect 13544 22559 13596 22568
rect 13544 22525 13553 22559
rect 13553 22525 13587 22559
rect 13587 22525 13596 22559
rect 13544 22516 13596 22525
rect 15844 22516 15896 22568
rect 10876 22448 10928 22500
rect 12440 22491 12492 22500
rect 12440 22457 12449 22491
rect 12449 22457 12483 22491
rect 12483 22457 12492 22491
rect 12440 22448 12492 22457
rect 2596 22380 2648 22432
rect 2872 22380 2924 22432
rect 3976 22380 4028 22432
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 6276 22423 6328 22432
rect 6276 22389 6285 22423
rect 6285 22389 6319 22423
rect 6319 22389 6328 22423
rect 6276 22380 6328 22389
rect 9036 22423 9088 22432
rect 9036 22389 9045 22423
rect 9045 22389 9079 22423
rect 9079 22389 9088 22423
rect 9036 22380 9088 22389
rect 9772 22380 9824 22432
rect 11980 22380 12032 22432
rect 13084 22423 13136 22432
rect 13084 22389 13093 22423
rect 13093 22389 13127 22423
rect 13127 22389 13136 22423
rect 14556 22448 14608 22500
rect 15936 22448 15988 22500
rect 17868 22448 17920 22500
rect 15568 22423 15620 22432
rect 13084 22380 13136 22389
rect 15568 22389 15577 22423
rect 15577 22389 15611 22423
rect 15611 22389 15620 22423
rect 15568 22380 15620 22389
rect 18880 22423 18932 22432
rect 18880 22389 18889 22423
rect 18889 22389 18923 22423
rect 18923 22389 18932 22423
rect 18880 22380 18932 22389
rect 20720 22380 20772 22432
rect 22192 22423 22244 22432
rect 22192 22389 22201 22423
rect 22201 22389 22235 22423
rect 22235 22389 22244 22423
rect 22192 22380 22244 22389
rect 23296 22423 23348 22432
rect 23296 22389 23305 22423
rect 23305 22389 23339 22423
rect 23339 22389 23348 22423
rect 23296 22380 23348 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1676 22219 1728 22228
rect 1676 22185 1685 22219
rect 1685 22185 1719 22219
rect 1719 22185 1728 22219
rect 1676 22176 1728 22185
rect 2136 22219 2188 22228
rect 2136 22185 2145 22219
rect 2145 22185 2179 22219
rect 2179 22185 2188 22219
rect 4712 22219 4764 22228
rect 2136 22176 2188 22185
rect 4712 22185 4721 22219
rect 4721 22185 4755 22219
rect 4755 22185 4764 22219
rect 4712 22176 4764 22185
rect 5172 22176 5224 22228
rect 5356 22151 5408 22160
rect 5356 22117 5365 22151
rect 5365 22117 5399 22151
rect 5399 22117 5408 22151
rect 5356 22108 5408 22117
rect 2228 22015 2280 22024
rect 2228 21981 2237 22015
rect 2237 21981 2271 22015
rect 2271 21981 2280 22015
rect 2228 21972 2280 21981
rect 2688 21972 2740 22024
rect 3056 22040 3108 22092
rect 6828 22176 6880 22228
rect 7564 22219 7616 22228
rect 7564 22185 7573 22219
rect 7573 22185 7607 22219
rect 7607 22185 7616 22219
rect 7564 22176 7616 22185
rect 8668 22219 8720 22228
rect 8668 22185 8677 22219
rect 8677 22185 8711 22219
rect 8711 22185 8720 22219
rect 8668 22176 8720 22185
rect 9036 22176 9088 22228
rect 9772 22176 9824 22228
rect 10784 22176 10836 22228
rect 12716 22176 12768 22228
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 9588 22040 9640 22092
rect 10692 22040 10744 22092
rect 11060 22083 11112 22092
rect 11060 22049 11069 22083
rect 11069 22049 11103 22083
rect 11103 22049 11112 22083
rect 11060 22040 11112 22049
rect 6184 21972 6236 22024
rect 6736 21972 6788 22024
rect 7840 21972 7892 22024
rect 8668 21972 8720 22024
rect 10968 21972 11020 22024
rect 10784 21904 10836 21956
rect 12072 21972 12124 22024
rect 12624 21972 12676 22024
rect 12256 21904 12308 21956
rect 13728 21972 13780 22024
rect 2136 21836 2188 21888
rect 3240 21836 3292 21888
rect 3424 21836 3476 21888
rect 4988 21879 5040 21888
rect 4988 21845 4997 21879
rect 4997 21845 5031 21879
rect 5031 21845 5040 21879
rect 4988 21836 5040 21845
rect 6644 21836 6696 21888
rect 8392 21836 8444 21888
rect 13176 21836 13228 21888
rect 13544 21879 13596 21888
rect 13544 21845 13553 21879
rect 13553 21845 13587 21879
rect 13587 21845 13596 21879
rect 13544 21836 13596 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2044 21675 2096 21684
rect 2044 21641 2053 21675
rect 2053 21641 2087 21675
rect 2087 21641 2096 21675
rect 2044 21632 2096 21641
rect 2688 21632 2740 21684
rect 5356 21632 5408 21684
rect 6552 21675 6604 21684
rect 6552 21641 6561 21675
rect 6561 21641 6595 21675
rect 6595 21641 6604 21675
rect 6552 21632 6604 21641
rect 6828 21675 6880 21684
rect 6828 21641 6837 21675
rect 6837 21641 6871 21675
rect 6871 21641 6880 21675
rect 6828 21632 6880 21641
rect 7840 21675 7892 21684
rect 7840 21641 7849 21675
rect 7849 21641 7883 21675
rect 7883 21641 7892 21675
rect 7840 21632 7892 21641
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12716 21675 12768 21684
rect 12716 21641 12725 21675
rect 12725 21641 12759 21675
rect 12759 21641 12768 21675
rect 12716 21632 12768 21641
rect 14556 21675 14608 21684
rect 14556 21641 14565 21675
rect 14565 21641 14599 21675
rect 14599 21641 14608 21675
rect 14556 21632 14608 21641
rect 3700 21539 3752 21548
rect 3700 21505 3709 21539
rect 3709 21505 3743 21539
rect 3743 21505 3752 21539
rect 3700 21496 3752 21505
rect 5724 21539 5776 21548
rect 2044 21428 2096 21480
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 10968 21564 11020 21616
rect 12624 21564 12676 21616
rect 7472 21539 7524 21548
rect 7472 21505 7481 21539
rect 7481 21505 7515 21539
rect 7515 21505 7524 21539
rect 7472 21496 7524 21505
rect 11796 21496 11848 21548
rect 6000 21428 6052 21480
rect 6920 21428 6972 21480
rect 3424 21360 3476 21412
rect 8668 21428 8720 21480
rect 1860 21292 1912 21344
rect 2044 21292 2096 21344
rect 2872 21292 2924 21344
rect 3240 21335 3292 21344
rect 3240 21301 3249 21335
rect 3249 21301 3283 21335
rect 3283 21301 3292 21335
rect 3240 21292 3292 21301
rect 5264 21292 5316 21344
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 5540 21292 5592 21301
rect 8024 21292 8076 21344
rect 9496 21360 9548 21412
rect 9956 21335 10008 21344
rect 9956 21301 9965 21335
rect 9965 21301 9999 21335
rect 9999 21301 10008 21335
rect 9956 21292 10008 21301
rect 11336 21335 11388 21344
rect 11336 21301 11345 21335
rect 11345 21301 11379 21335
rect 11379 21301 11388 21335
rect 11336 21292 11388 21301
rect 12716 21292 12768 21344
rect 13544 21360 13596 21412
rect 14096 21360 14148 21412
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 2228 21088 2280 21140
rect 6736 21088 6788 21140
rect 9956 21088 10008 21140
rect 10784 21131 10836 21140
rect 10784 21097 10793 21131
rect 10793 21097 10827 21131
rect 10827 21097 10836 21131
rect 10784 21088 10836 21097
rect 11336 21088 11388 21140
rect 14096 21131 14148 21140
rect 14096 21097 14105 21131
rect 14105 21097 14139 21131
rect 14139 21097 14148 21131
rect 14096 21088 14148 21097
rect 1492 21020 1544 21072
rect 1952 21063 2004 21072
rect 1952 21029 1961 21063
rect 1961 21029 1995 21063
rect 1995 21029 2004 21063
rect 1952 21020 2004 21029
rect 6276 21020 6328 21072
rect 6920 21020 6972 21072
rect 13084 21020 13136 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 3976 20952 4028 21004
rect 9680 20995 9732 21004
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9680 20952 9732 20961
rect 2688 20859 2740 20868
rect 2688 20825 2697 20859
rect 2697 20825 2731 20859
rect 2731 20825 2740 20859
rect 2688 20816 2740 20825
rect 2228 20748 2280 20800
rect 3792 20791 3844 20800
rect 3792 20757 3801 20791
rect 3801 20757 3835 20791
rect 3835 20757 3844 20791
rect 3792 20748 3844 20757
rect 3976 20748 4028 20800
rect 5448 20884 5500 20936
rect 5724 20816 5776 20868
rect 5080 20748 5132 20800
rect 11060 20884 11112 20936
rect 11796 20927 11848 20936
rect 7656 20816 7708 20868
rect 8116 20816 8168 20868
rect 11796 20893 11805 20927
rect 11805 20893 11839 20927
rect 11839 20893 11848 20927
rect 11796 20884 11848 20893
rect 11980 20884 12032 20936
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 12348 20816 12400 20868
rect 6736 20748 6788 20800
rect 7840 20748 7892 20800
rect 8576 20791 8628 20800
rect 8576 20757 8585 20791
rect 8585 20757 8619 20791
rect 8619 20757 8628 20791
rect 8576 20748 8628 20757
rect 10140 20748 10192 20800
rect 11704 20748 11756 20800
rect 12532 20791 12584 20800
rect 12532 20757 12541 20791
rect 12541 20757 12575 20791
rect 12575 20757 12584 20791
rect 12532 20748 12584 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1400 20544 1452 20596
rect 2964 20544 3016 20596
rect 3976 20587 4028 20596
rect 3976 20553 3985 20587
rect 3985 20553 4019 20587
rect 4019 20553 4028 20587
rect 3976 20544 4028 20553
rect 5540 20587 5592 20596
rect 5540 20553 5549 20587
rect 5549 20553 5583 20587
rect 5583 20553 5592 20587
rect 5540 20544 5592 20553
rect 6092 20544 6144 20596
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 4896 20408 4948 20460
rect 2228 20383 2280 20392
rect 2228 20349 2262 20383
rect 2262 20349 2280 20383
rect 2228 20340 2280 20349
rect 4804 20383 4856 20392
rect 4804 20349 4813 20383
rect 4813 20349 4847 20383
rect 4847 20349 4856 20383
rect 4804 20340 4856 20349
rect 6920 20544 6972 20596
rect 11060 20544 11112 20596
rect 11336 20587 11388 20596
rect 11336 20553 11345 20587
rect 11345 20553 11379 20587
rect 11379 20553 11388 20587
rect 11336 20544 11388 20553
rect 11980 20544 12032 20596
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 13820 20587 13872 20596
rect 12440 20544 12492 20553
rect 13820 20553 13829 20587
rect 13829 20553 13863 20587
rect 13863 20553 13872 20587
rect 13820 20544 13872 20553
rect 9404 20476 9456 20528
rect 9956 20476 10008 20528
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 12808 20476 12860 20528
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 13084 20408 13136 20417
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 8116 20383 8168 20392
rect 8116 20349 8150 20383
rect 8150 20349 8168 20383
rect 1952 20272 2004 20324
rect 3976 20272 4028 20324
rect 4068 20272 4120 20324
rect 5448 20272 5500 20324
rect 8116 20340 8168 20349
rect 12532 20340 12584 20392
rect 13820 20340 13872 20392
rect 8024 20272 8076 20324
rect 10692 20315 10744 20324
rect 10692 20281 10701 20315
rect 10701 20281 10735 20315
rect 10735 20281 10744 20315
rect 10692 20272 10744 20281
rect 4436 20247 4488 20256
rect 4436 20213 4445 20247
rect 4445 20213 4479 20247
rect 4479 20213 4488 20247
rect 4436 20204 4488 20213
rect 6736 20204 6788 20256
rect 7012 20247 7064 20256
rect 7012 20213 7021 20247
rect 7021 20213 7055 20247
rect 7055 20213 7064 20247
rect 7012 20204 7064 20213
rect 9220 20247 9272 20256
rect 9220 20213 9229 20247
rect 9229 20213 9263 20247
rect 9263 20213 9272 20247
rect 9220 20204 9272 20213
rect 9772 20204 9824 20256
rect 14004 20247 14056 20256
rect 14004 20213 14013 20247
rect 14013 20213 14047 20247
rect 14047 20213 14056 20247
rect 14004 20204 14056 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2228 20000 2280 20052
rect 2596 20000 2648 20052
rect 3240 20000 3292 20052
rect 4804 20000 4856 20052
rect 5448 20043 5500 20052
rect 5448 20009 5457 20043
rect 5457 20009 5491 20043
rect 5491 20009 5500 20043
rect 5448 20000 5500 20009
rect 8116 20000 8168 20052
rect 8300 20000 8352 20052
rect 10692 20000 10744 20052
rect 11796 20043 11848 20052
rect 11796 20009 11805 20043
rect 11805 20009 11839 20043
rect 11839 20009 11848 20043
rect 11796 20000 11848 20009
rect 13084 20000 13136 20052
rect 1676 19932 1728 19984
rect 1952 19932 2004 19984
rect 6184 19932 6236 19984
rect 7840 19932 7892 19984
rect 2964 19864 3016 19916
rect 6736 19864 6788 19916
rect 9864 19864 9916 19916
rect 11060 19864 11112 19916
rect 11980 19864 12032 19916
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 12624 19907 12676 19916
rect 12624 19873 12658 19907
rect 12658 19873 12676 19907
rect 12624 19864 12676 19873
rect 11244 19839 11296 19848
rect 5080 19728 5132 19780
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 15292 19839 15344 19848
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 15292 19796 15344 19805
rect 9680 19728 9732 19780
rect 3148 19660 3200 19712
rect 4896 19703 4948 19712
rect 4896 19669 4905 19703
rect 4905 19669 4939 19703
rect 4939 19669 4948 19703
rect 4896 19660 4948 19669
rect 5172 19660 5224 19712
rect 9312 19660 9364 19712
rect 10140 19660 10192 19712
rect 10784 19703 10836 19712
rect 10784 19669 10793 19703
rect 10793 19669 10827 19703
rect 10827 19669 10836 19703
rect 10784 19660 10836 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2596 19499 2648 19508
rect 2596 19465 2605 19499
rect 2605 19465 2639 19499
rect 2639 19465 2648 19499
rect 2596 19456 2648 19465
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 3148 19499 3200 19508
rect 3148 19465 3157 19499
rect 3157 19465 3191 19499
rect 3191 19465 3200 19499
rect 3148 19456 3200 19465
rect 4804 19456 4856 19508
rect 9772 19456 9824 19508
rect 10048 19456 10100 19508
rect 11428 19499 11480 19508
rect 11428 19465 11437 19499
rect 11437 19465 11471 19499
rect 11471 19465 11480 19499
rect 11428 19456 11480 19465
rect 12624 19456 12676 19508
rect 3240 19320 3292 19372
rect 3148 19252 3200 19304
rect 3516 19295 3568 19304
rect 3516 19261 3525 19295
rect 3525 19261 3559 19295
rect 3559 19261 3568 19295
rect 4436 19320 4488 19372
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 5172 19295 5224 19304
rect 3516 19252 3568 19261
rect 2412 19184 2464 19236
rect 5172 19261 5181 19295
rect 5181 19261 5215 19295
rect 5215 19261 5224 19295
rect 5172 19252 5224 19261
rect 5264 19295 5316 19304
rect 5264 19261 5273 19295
rect 5273 19261 5307 19295
rect 5307 19261 5316 19295
rect 5264 19252 5316 19261
rect 5540 19252 5592 19304
rect 6184 19295 6236 19304
rect 6184 19261 6193 19295
rect 6193 19261 6227 19295
rect 6227 19261 6236 19295
rect 6184 19252 6236 19261
rect 7932 19295 7984 19304
rect 7932 19261 7941 19295
rect 7941 19261 7975 19295
rect 7975 19261 7984 19295
rect 7932 19252 7984 19261
rect 10048 19320 10100 19372
rect 10784 19320 10836 19372
rect 19432 19320 19484 19372
rect 19984 19320 20036 19372
rect 20720 19320 20772 19372
rect 20904 19320 20956 19372
rect 8944 19295 8996 19304
rect 8944 19261 8953 19295
rect 8953 19261 8987 19295
rect 8987 19261 8996 19295
rect 8944 19252 8996 19261
rect 12532 19252 12584 19304
rect 14096 19252 14148 19304
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 4344 19159 4396 19168
rect 4344 19125 4353 19159
rect 4353 19125 4387 19159
rect 4387 19125 4396 19159
rect 4344 19116 4396 19125
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 6828 19116 6880 19168
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 7564 19116 7616 19168
rect 9220 19184 9272 19236
rect 9864 19184 9916 19236
rect 10232 19184 10284 19236
rect 12716 19227 12768 19236
rect 12716 19193 12750 19227
rect 12750 19193 12768 19227
rect 12716 19184 12768 19193
rect 10784 19116 10836 19168
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 15108 19159 15160 19168
rect 15108 19125 15117 19159
rect 15117 19125 15151 19159
rect 15151 19125 15160 19159
rect 15108 19116 15160 19125
rect 15844 19116 15896 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1676 18955 1728 18964
rect 1676 18921 1685 18955
rect 1685 18921 1719 18955
rect 1719 18921 1728 18955
rect 1676 18912 1728 18921
rect 2964 18912 3016 18964
rect 3516 18955 3568 18964
rect 3516 18921 3525 18955
rect 3525 18921 3559 18955
rect 3559 18921 3568 18955
rect 3516 18912 3568 18921
rect 5264 18912 5316 18964
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 9220 18912 9272 18964
rect 11244 18912 11296 18964
rect 13360 18912 13412 18964
rect 5356 18844 5408 18896
rect 5540 18844 5592 18896
rect 7472 18844 7524 18896
rect 9772 18844 9824 18896
rect 1400 18776 1452 18828
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 7656 18776 7708 18828
rect 8116 18819 8168 18828
rect 8116 18785 8125 18819
rect 8125 18785 8159 18819
rect 8159 18785 8168 18819
rect 10784 18819 10836 18828
rect 8116 18776 8168 18785
rect 10784 18785 10818 18819
rect 10818 18785 10836 18819
rect 10784 18776 10836 18785
rect 13360 18819 13412 18828
rect 13360 18785 13369 18819
rect 13369 18785 13403 18819
rect 13403 18785 13412 18819
rect 13360 18776 13412 18785
rect 2228 18751 2280 18760
rect 2228 18717 2237 18751
rect 2237 18717 2271 18751
rect 2271 18717 2280 18751
rect 2228 18708 2280 18717
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 2964 18708 3016 18760
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 9220 18708 9272 18760
rect 15292 18751 15344 18760
rect 1952 18572 2004 18624
rect 2688 18572 2740 18624
rect 2872 18615 2924 18624
rect 2872 18581 2881 18615
rect 2881 18581 2915 18615
rect 2915 18581 2924 18615
rect 2872 18572 2924 18581
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 5172 18572 5224 18624
rect 6920 18572 6972 18624
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 12256 18640 12308 18692
rect 12716 18640 12768 18692
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 16304 18751 16356 18760
rect 16304 18717 16313 18751
rect 16313 18717 16347 18751
rect 16347 18717 16356 18751
rect 16304 18708 16356 18717
rect 10692 18572 10744 18624
rect 11796 18572 11848 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 13636 18572 13688 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1676 18368 1728 18420
rect 2964 18368 3016 18420
rect 4344 18368 4396 18420
rect 8208 18411 8260 18420
rect 8208 18377 8217 18411
rect 8217 18377 8251 18411
rect 8251 18377 8260 18411
rect 8208 18368 8260 18377
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 10784 18368 10836 18420
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 13360 18411 13412 18420
rect 13360 18377 13369 18411
rect 13369 18377 13403 18411
rect 13403 18377 13412 18411
rect 13360 18368 13412 18377
rect 24768 18368 24820 18420
rect 9220 18300 9272 18352
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 6092 18275 6144 18284
rect 5356 18232 5408 18241
rect 6092 18241 6101 18275
rect 6101 18241 6135 18275
rect 6135 18241 6144 18275
rect 6092 18232 6144 18241
rect 9772 18275 9824 18284
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 11888 18300 11940 18352
rect 13268 18300 13320 18352
rect 14924 18343 14976 18352
rect 14924 18309 14933 18343
rect 14933 18309 14967 18343
rect 14967 18309 14976 18343
rect 14924 18300 14976 18309
rect 11060 18232 11112 18284
rect 2872 18164 2924 18216
rect 5080 18207 5132 18216
rect 5080 18173 5089 18207
rect 5089 18173 5123 18207
rect 5123 18173 5132 18207
rect 5080 18164 5132 18173
rect 5540 18164 5592 18216
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 8944 18164 8996 18216
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 10968 18164 11020 18216
rect 13636 18164 13688 18216
rect 23664 18207 23716 18216
rect 4988 18096 5040 18148
rect 6920 18096 6972 18148
rect 13820 18139 13872 18148
rect 13820 18105 13854 18139
rect 13854 18105 13872 18139
rect 13820 18096 13872 18105
rect 1400 18028 1452 18080
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 10692 18028 10744 18080
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 23664 18173 23673 18207
rect 23673 18173 23707 18207
rect 23707 18173 23716 18207
rect 23664 18164 23716 18173
rect 17040 18028 17092 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2228 17867 2280 17876
rect 2228 17833 2237 17867
rect 2237 17833 2271 17867
rect 2271 17833 2280 17867
rect 2228 17824 2280 17833
rect 2780 17824 2832 17876
rect 3884 17824 3936 17876
rect 4068 17824 4120 17876
rect 2044 17756 2096 17808
rect 4436 17756 4488 17808
rect 2320 17688 2372 17740
rect 2228 17620 2280 17672
rect 4620 17688 4672 17740
rect 5540 17824 5592 17876
rect 6092 17867 6144 17876
rect 6092 17833 6101 17867
rect 6101 17833 6135 17867
rect 6135 17833 6144 17867
rect 6092 17824 6144 17833
rect 7656 17867 7708 17876
rect 7656 17833 7665 17867
rect 7665 17833 7699 17867
rect 7699 17833 7708 17867
rect 7656 17824 7708 17833
rect 9588 17824 9640 17876
rect 12256 17824 12308 17876
rect 13452 17867 13504 17876
rect 13452 17833 13461 17867
rect 13461 17833 13495 17867
rect 13495 17833 13504 17867
rect 13452 17824 13504 17833
rect 17040 17867 17092 17876
rect 17040 17833 17049 17867
rect 17049 17833 17083 17867
rect 17083 17833 17092 17867
rect 17040 17824 17092 17833
rect 5172 17756 5224 17808
rect 8116 17756 8168 17808
rect 8208 17756 8260 17808
rect 9496 17756 9548 17808
rect 10784 17756 10836 17808
rect 5356 17688 5408 17740
rect 8024 17731 8076 17740
rect 8024 17697 8033 17731
rect 8033 17697 8067 17731
rect 8067 17697 8076 17731
rect 8024 17688 8076 17697
rect 10692 17688 10744 17740
rect 11152 17688 11204 17740
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 17868 17731 17920 17740
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2964 17663 3016 17672
rect 2780 17620 2832 17629
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 8116 17663 8168 17672
rect 8116 17629 8125 17663
rect 8125 17629 8159 17663
rect 8159 17629 8168 17663
rect 8116 17620 8168 17629
rect 8300 17663 8352 17672
rect 8300 17629 8309 17663
rect 8309 17629 8343 17663
rect 8343 17629 8352 17663
rect 8300 17620 8352 17629
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 15384 17620 15436 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 2044 17552 2096 17604
rect 13084 17595 13136 17604
rect 13084 17561 13093 17595
rect 13093 17561 13127 17595
rect 13127 17561 13136 17595
rect 13084 17552 13136 17561
rect 17868 17697 17877 17731
rect 17877 17697 17911 17731
rect 17911 17697 17920 17731
rect 17868 17688 17920 17697
rect 17224 17552 17276 17604
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 9680 17484 9732 17536
rect 12992 17484 13044 17536
rect 17960 17484 18012 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 2044 17323 2096 17332
rect 2044 17289 2053 17323
rect 2053 17289 2087 17323
rect 2087 17289 2096 17323
rect 2044 17280 2096 17289
rect 2228 17323 2280 17332
rect 2228 17289 2237 17323
rect 2237 17289 2271 17323
rect 2271 17289 2280 17323
rect 2228 17280 2280 17289
rect 3516 17323 3568 17332
rect 3516 17289 3525 17323
rect 3525 17289 3559 17323
rect 3559 17289 3568 17323
rect 3516 17280 3568 17289
rect 4160 17280 4212 17332
rect 5540 17280 5592 17332
rect 7564 17323 7616 17332
rect 7564 17289 7573 17323
rect 7573 17289 7607 17323
rect 7607 17289 7616 17323
rect 7564 17280 7616 17289
rect 2504 17212 2556 17264
rect 2780 17212 2832 17264
rect 5448 17212 5500 17264
rect 3884 17144 3936 17196
rect 6920 17144 6972 17196
rect 10784 17280 10836 17332
rect 13728 17280 13780 17332
rect 15660 17280 15712 17332
rect 17224 17323 17276 17332
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 17868 17280 17920 17332
rect 8300 17212 8352 17264
rect 8944 17255 8996 17264
rect 8944 17221 8953 17255
rect 8953 17221 8987 17255
rect 8987 17221 8996 17255
rect 8944 17212 8996 17221
rect 19340 17212 19392 17264
rect 20260 17212 20312 17264
rect 18052 17187 18104 17196
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 3516 17076 3568 17128
rect 4712 17076 4764 17128
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 8208 17076 8260 17128
rect 9404 17119 9456 17128
rect 9404 17085 9438 17119
rect 9438 17085 9456 17119
rect 9404 17076 9456 17085
rect 4988 17008 5040 17060
rect 3056 16940 3108 16992
rect 4804 16940 4856 16992
rect 5356 16940 5408 16992
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 13084 17051 13136 17060
rect 13084 17017 13118 17051
rect 13118 17017 13136 17051
rect 13084 17008 13136 17017
rect 13636 16940 13688 16992
rect 15844 17076 15896 17128
rect 16212 16940 16264 16992
rect 16580 16940 16632 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1400 16779 1452 16788
rect 1400 16745 1409 16779
rect 1409 16745 1443 16779
rect 1443 16745 1452 16779
rect 1400 16736 1452 16745
rect 2688 16736 2740 16788
rect 4712 16736 4764 16788
rect 5448 16736 5500 16788
rect 7932 16736 7984 16788
rect 9404 16736 9456 16788
rect 9680 16736 9732 16788
rect 11428 16779 11480 16788
rect 11428 16745 11437 16779
rect 11437 16745 11471 16779
rect 11471 16745 11480 16779
rect 11428 16736 11480 16745
rect 13544 16736 13596 16788
rect 14280 16779 14332 16788
rect 14280 16745 14289 16779
rect 14289 16745 14323 16779
rect 14323 16745 14332 16779
rect 14280 16736 14332 16745
rect 15476 16779 15528 16788
rect 15476 16745 15485 16779
rect 15485 16745 15519 16779
rect 15519 16745 15528 16779
rect 15476 16736 15528 16745
rect 15844 16779 15896 16788
rect 15844 16745 15853 16779
rect 15853 16745 15887 16779
rect 15887 16745 15896 16779
rect 15844 16736 15896 16745
rect 19432 16736 19484 16788
rect 4804 16668 4856 16720
rect 4896 16668 4948 16720
rect 7012 16668 7064 16720
rect 7380 16668 7432 16720
rect 8116 16668 8168 16720
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 2780 16600 2832 16609
rect 2228 16396 2280 16448
rect 2412 16439 2464 16448
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 4988 16600 5040 16652
rect 5080 16643 5132 16652
rect 5080 16609 5089 16643
rect 5089 16609 5123 16643
rect 5123 16609 5132 16643
rect 6368 16643 6420 16652
rect 5080 16600 5132 16609
rect 6368 16609 6377 16643
rect 6377 16609 6411 16643
rect 6411 16609 6420 16643
rect 6368 16600 6420 16609
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 8024 16600 8076 16652
rect 8392 16643 8444 16652
rect 8392 16609 8401 16643
rect 8401 16609 8435 16643
rect 8435 16609 8444 16643
rect 8392 16600 8444 16609
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 6552 16464 6604 16516
rect 9404 16532 9456 16584
rect 9772 16600 9824 16652
rect 13452 16711 13504 16720
rect 13452 16677 13461 16711
rect 13461 16677 13495 16711
rect 13495 16677 13504 16711
rect 13452 16668 13504 16677
rect 13728 16668 13780 16720
rect 15384 16668 15436 16720
rect 16856 16668 16908 16720
rect 12256 16600 12308 16652
rect 10692 16532 10744 16584
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 13084 16600 13136 16652
rect 14188 16600 14240 16652
rect 14648 16600 14700 16652
rect 16120 16600 16172 16652
rect 19156 16643 19208 16652
rect 19156 16609 19165 16643
rect 19165 16609 19199 16643
rect 19199 16609 19208 16643
rect 19156 16600 19208 16609
rect 12440 16532 12492 16541
rect 12348 16464 12400 16516
rect 16212 16532 16264 16584
rect 22100 16600 22152 16652
rect 22468 16600 22520 16652
rect 19892 16532 19944 16584
rect 3884 16396 3936 16448
rect 5264 16396 5316 16448
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 9956 16396 10008 16448
rect 10968 16439 11020 16448
rect 10968 16405 10977 16439
rect 10977 16405 11011 16439
rect 11011 16405 11020 16439
rect 10968 16396 11020 16405
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 14740 16396 14792 16448
rect 15384 16396 15436 16448
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 3148 16192 3200 16244
rect 5080 16192 5132 16244
rect 5356 16192 5408 16244
rect 6276 16192 6328 16244
rect 5448 16124 5500 16176
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 2872 16056 2924 16108
rect 3884 16099 3936 16108
rect 3884 16065 3893 16099
rect 3893 16065 3927 16099
rect 3927 16065 3936 16099
rect 3884 16056 3936 16065
rect 5264 16056 5316 16108
rect 7380 16192 7432 16244
rect 9404 16192 9456 16244
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 13728 16192 13780 16244
rect 15844 16192 15896 16244
rect 19892 16235 19944 16244
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 20628 16235 20680 16244
rect 20628 16201 20637 16235
rect 20637 16201 20671 16235
rect 20671 16201 20680 16235
rect 20628 16192 20680 16201
rect 6828 16124 6880 16176
rect 8944 16124 8996 16176
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 7840 16056 7892 16108
rect 8392 16056 8444 16108
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 13176 16056 13228 16108
rect 13636 16056 13688 16108
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 3608 16031 3660 16040
rect 3608 15997 3617 16031
rect 3617 15997 3651 16031
rect 3651 15997 3660 16031
rect 3608 15988 3660 15997
rect 4620 15988 4672 16040
rect 6460 15988 6512 16040
rect 2136 15963 2188 15972
rect 2136 15929 2145 15963
rect 2145 15929 2179 15963
rect 2179 15929 2188 15963
rect 2136 15920 2188 15929
rect 2688 15920 2740 15972
rect 9220 15920 9272 15972
rect 11612 15920 11664 15972
rect 12440 15920 12492 15972
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 14924 16031 14976 16040
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2780 15895 2832 15904
rect 2780 15861 2789 15895
rect 2789 15861 2823 15895
rect 2823 15861 2832 15895
rect 2780 15852 2832 15861
rect 3332 15852 3384 15904
rect 3700 15895 3752 15904
rect 3700 15861 3709 15895
rect 3709 15861 3743 15895
rect 3743 15861 3752 15895
rect 3700 15852 3752 15861
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6000 15852 6052 15904
rect 7012 15852 7064 15904
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10692 15852 10744 15904
rect 10968 15895 11020 15904
rect 10968 15861 10977 15895
rect 10977 15861 11011 15895
rect 11011 15861 11020 15895
rect 10968 15852 11020 15861
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 12256 15852 12308 15904
rect 12624 15852 12676 15904
rect 14924 15997 14958 16031
rect 14958 15997 14976 16031
rect 14924 15988 14976 15997
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 19064 16031 19116 16040
rect 19064 15997 19073 16031
rect 19073 15997 19107 16031
rect 19107 15997 19116 16031
rect 19064 15988 19116 15997
rect 20444 16031 20496 16040
rect 20444 15997 20453 16031
rect 20453 15997 20487 16031
rect 20487 15997 20496 16031
rect 20444 15988 20496 15997
rect 14648 15852 14700 15904
rect 16212 15852 16264 15904
rect 16856 15852 16908 15904
rect 18236 15895 18288 15904
rect 18236 15861 18245 15895
rect 18245 15861 18279 15895
rect 18279 15861 18288 15895
rect 18236 15852 18288 15861
rect 19248 15895 19300 15904
rect 19248 15861 19257 15895
rect 19257 15861 19291 15895
rect 19291 15861 19300 15895
rect 19248 15852 19300 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 3608 15648 3660 15700
rect 4620 15691 4672 15700
rect 4620 15657 4629 15691
rect 4629 15657 4663 15691
rect 4663 15657 4672 15691
rect 4620 15648 4672 15657
rect 6920 15648 6972 15700
rect 4160 15580 4212 15632
rect 4528 15580 4580 15632
rect 7012 15623 7064 15632
rect 7012 15589 7021 15623
rect 7021 15589 7055 15623
rect 7055 15589 7064 15623
rect 7012 15580 7064 15589
rect 8392 15648 8444 15700
rect 8944 15691 8996 15700
rect 8944 15657 8953 15691
rect 8953 15657 8987 15691
rect 8987 15657 8996 15691
rect 8944 15648 8996 15657
rect 12348 15691 12400 15700
rect 12348 15657 12357 15691
rect 12357 15657 12391 15691
rect 12391 15657 12400 15691
rect 12348 15648 12400 15657
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 14924 15648 14976 15700
rect 15568 15648 15620 15700
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 16856 15648 16908 15700
rect 10048 15580 10100 15632
rect 10876 15580 10928 15632
rect 13360 15580 13412 15632
rect 1768 15555 1820 15564
rect 1768 15521 1802 15555
rect 1802 15521 1820 15555
rect 4712 15555 4764 15564
rect 1768 15512 1820 15521
rect 4712 15521 4721 15555
rect 4721 15521 4755 15555
rect 4755 15521 4764 15555
rect 4712 15512 4764 15521
rect 5264 15512 5316 15564
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 8300 15512 8352 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 17408 15512 17460 15564
rect 7288 15444 7340 15496
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 12440 15444 12492 15496
rect 12808 15419 12860 15428
rect 12808 15385 12817 15419
rect 12817 15385 12851 15419
rect 12851 15385 12860 15419
rect 12808 15376 12860 15385
rect 13176 15376 13228 15428
rect 16212 15444 16264 15496
rect 1676 15308 1728 15360
rect 3884 15351 3936 15360
rect 3884 15317 3893 15351
rect 3893 15317 3927 15351
rect 3927 15317 3936 15351
rect 3884 15308 3936 15317
rect 4620 15308 4672 15360
rect 9220 15308 9272 15360
rect 10048 15308 10100 15360
rect 11704 15351 11756 15360
rect 11704 15317 11713 15351
rect 11713 15317 11747 15351
rect 11747 15317 11756 15351
rect 11704 15308 11756 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1492 15104 1544 15156
rect 3148 15104 3200 15156
rect 4712 15104 4764 15156
rect 4988 15036 5040 15088
rect 6552 15104 6604 15156
rect 8300 15104 8352 15156
rect 9036 15104 9088 15156
rect 10876 15104 10928 15156
rect 12348 15104 12400 15156
rect 17408 15147 17460 15156
rect 17408 15113 17417 15147
rect 17417 15113 17451 15147
rect 17451 15113 17460 15147
rect 17408 15104 17460 15113
rect 20444 15104 20496 15156
rect 6368 14968 6420 15020
rect 2688 14900 2740 14952
rect 3148 14943 3200 14952
rect 3148 14909 3182 14943
rect 3182 14909 3200 14943
rect 1676 14832 1728 14884
rect 3148 14900 3200 14909
rect 3884 14900 3936 14952
rect 5448 14900 5500 14952
rect 6460 14943 6512 14952
rect 6460 14909 6469 14943
rect 6469 14909 6503 14943
rect 6503 14909 6512 14943
rect 6460 14900 6512 14909
rect 16856 14968 16908 15020
rect 4712 14832 4764 14884
rect 7840 14900 7892 14952
rect 8944 14832 8996 14884
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 10324 14900 10376 14952
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 19432 14943 19484 14952
rect 13912 14900 13964 14909
rect 10048 14875 10100 14884
rect 10048 14841 10082 14875
rect 10082 14841 10100 14875
rect 10048 14832 10100 14841
rect 10692 14832 10744 14884
rect 13176 14832 13228 14884
rect 14004 14832 14056 14884
rect 19432 14909 19441 14943
rect 19441 14909 19475 14943
rect 19475 14909 19484 14943
rect 19432 14900 19484 14909
rect 16764 14875 16816 14884
rect 16764 14841 16773 14875
rect 16773 14841 16807 14875
rect 16807 14841 16816 14875
rect 16764 14832 16816 14841
rect 11888 14764 11940 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 15476 14764 15528 14816
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 16488 14764 16540 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1768 14560 1820 14612
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 2136 14560 2188 14612
rect 2688 14560 2740 14612
rect 4436 14603 4488 14612
rect 3332 14492 3384 14544
rect 3792 14492 3844 14544
rect 4436 14569 4445 14603
rect 4445 14569 4479 14603
rect 4479 14569 4488 14603
rect 4436 14560 4488 14569
rect 4528 14603 4580 14612
rect 4528 14569 4537 14603
rect 4537 14569 4571 14603
rect 4571 14569 4580 14603
rect 4528 14560 4580 14569
rect 5264 14560 5316 14612
rect 10048 14603 10100 14612
rect 10048 14569 10057 14603
rect 10057 14569 10091 14603
rect 10091 14569 10100 14603
rect 10048 14560 10100 14569
rect 10876 14560 10928 14612
rect 14004 14603 14056 14612
rect 14004 14569 14013 14603
rect 14013 14569 14047 14603
rect 14047 14569 14056 14603
rect 14004 14560 14056 14569
rect 15384 14560 15436 14612
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 16764 14560 16816 14612
rect 4896 14492 4948 14544
rect 6552 14492 6604 14544
rect 12072 14535 12124 14544
rect 12072 14501 12106 14535
rect 12106 14501 12124 14535
rect 12072 14492 12124 14501
rect 15200 14492 15252 14544
rect 16304 14535 16356 14544
rect 16304 14501 16313 14535
rect 16313 14501 16347 14535
rect 16347 14501 16356 14535
rect 16304 14492 16356 14501
rect 3240 14424 3292 14476
rect 6092 14467 6144 14476
rect 6092 14433 6108 14467
rect 6108 14433 6142 14467
rect 6142 14433 6144 14467
rect 8392 14467 8444 14476
rect 6092 14424 6144 14433
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 10324 14424 10376 14476
rect 11888 14424 11940 14476
rect 16856 14424 16908 14476
rect 3148 14356 3200 14408
rect 4620 14399 4672 14408
rect 3240 14288 3292 14340
rect 2504 14220 2556 14272
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 9588 14288 9640 14340
rect 4988 14220 5040 14272
rect 5448 14263 5500 14272
rect 5448 14229 5457 14263
rect 5457 14229 5491 14263
rect 5491 14229 5500 14263
rect 5448 14220 5500 14229
rect 6368 14220 6420 14272
rect 7288 14220 7340 14272
rect 9680 14263 9732 14272
rect 9680 14229 9689 14263
rect 9689 14229 9723 14263
rect 9723 14229 9732 14263
rect 9680 14220 9732 14229
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 13176 14220 13228 14229
rect 14004 14220 14056 14272
rect 15568 14288 15620 14340
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 4344 14059 4396 14068
rect 4344 14025 4353 14059
rect 4353 14025 4387 14059
rect 4387 14025 4396 14059
rect 4344 14016 4396 14025
rect 4436 14016 4488 14068
rect 6184 14059 6236 14068
rect 4528 13948 4580 14000
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 6368 14016 6420 14068
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 6920 14016 6972 14068
rect 8944 14059 8996 14068
rect 2504 13880 2556 13932
rect 2964 13880 3016 13932
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 4988 13923 5040 13932
rect 4988 13889 4997 13923
rect 4997 13889 5031 13923
rect 5031 13889 5040 13923
rect 4988 13880 5040 13889
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 10048 14016 10100 14068
rect 11428 14059 11480 14068
rect 11428 14025 11437 14059
rect 11437 14025 11471 14059
rect 11471 14025 11480 14059
rect 11428 14016 11480 14025
rect 12072 14016 12124 14068
rect 14096 14016 14148 14068
rect 15568 14016 15620 14068
rect 15660 14016 15712 14068
rect 16488 14016 16540 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 8116 13880 8168 13932
rect 10324 13948 10376 14000
rect 12716 13948 12768 14000
rect 15016 13948 15068 14000
rect 7472 13812 7524 13864
rect 8300 13812 8352 13864
rect 4068 13744 4120 13796
rect 13360 13880 13412 13932
rect 16304 13880 16356 13932
rect 17040 13880 17092 13932
rect 13452 13812 13504 13864
rect 13912 13812 13964 13864
rect 9588 13744 9640 13796
rect 14648 13744 14700 13796
rect 2596 13676 2648 13728
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 4712 13676 4764 13685
rect 5540 13676 5592 13728
rect 7564 13719 7616 13728
rect 7564 13685 7573 13719
rect 7573 13685 7607 13719
rect 7607 13685 7616 13719
rect 7564 13676 7616 13685
rect 10692 13676 10744 13728
rect 11888 13719 11940 13728
rect 11888 13685 11897 13719
rect 11897 13685 11931 13719
rect 11931 13685 11940 13719
rect 11888 13676 11940 13685
rect 16120 13719 16172 13728
rect 16120 13685 16129 13719
rect 16129 13685 16163 13719
rect 16163 13685 16172 13719
rect 16120 13676 16172 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 848 13472 900 13524
rect 3148 13515 3200 13524
rect 2596 13404 2648 13456
rect 3148 13481 3157 13515
rect 3157 13481 3191 13515
rect 3191 13481 3200 13515
rect 3148 13472 3200 13481
rect 3884 13515 3936 13524
rect 3884 13481 3893 13515
rect 3893 13481 3927 13515
rect 3927 13481 3936 13515
rect 3884 13472 3936 13481
rect 4252 13472 4304 13524
rect 4712 13472 4764 13524
rect 6000 13472 6052 13524
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 8116 13515 8168 13524
rect 8116 13481 8125 13515
rect 8125 13481 8159 13515
rect 8159 13481 8168 13515
rect 8116 13472 8168 13481
rect 9956 13472 10008 13524
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 13820 13472 13872 13524
rect 15016 13515 15068 13524
rect 15016 13481 15025 13515
rect 15025 13481 15059 13515
rect 15059 13481 15068 13515
rect 15016 13472 15068 13481
rect 17040 13472 17092 13524
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 21180 13472 21232 13524
rect 4620 13404 4672 13456
rect 7104 13404 7156 13456
rect 7288 13404 7340 13456
rect 1952 13336 2004 13388
rect 7840 13336 7892 13388
rect 8760 13336 8812 13388
rect 9680 13336 9732 13388
rect 11520 13336 11572 13388
rect 13176 13336 13228 13388
rect 16212 13336 16264 13388
rect 18144 13336 18196 13388
rect 20812 13336 20864 13388
rect 3976 13200 4028 13252
rect 6184 13268 6236 13320
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 10692 13268 10744 13320
rect 11888 13268 11940 13320
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 17960 13268 18012 13320
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 2228 13132 2280 13184
rect 3884 13132 3936 13184
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 7288 13175 7340 13184
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 9588 13132 9640 13184
rect 13360 13175 13412 13184
rect 13360 13141 13369 13175
rect 13369 13141 13403 13175
rect 13403 13141 13412 13175
rect 13360 13132 13412 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 3516 12928 3568 12980
rect 3976 12971 4028 12980
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 4528 12928 4580 12980
rect 4620 12903 4672 12912
rect 4620 12869 4629 12903
rect 4629 12869 4663 12903
rect 4663 12869 4672 12903
rect 4620 12860 4672 12869
rect 5080 12860 5132 12912
rect 6276 12928 6328 12980
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 9220 12971 9272 12980
rect 9220 12937 9229 12971
rect 9229 12937 9263 12971
rect 9263 12937 9272 12971
rect 9220 12928 9272 12937
rect 10140 12928 10192 12980
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 14004 12971 14056 12980
rect 12440 12928 12492 12937
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 15936 12928 15988 12980
rect 22008 12928 22060 12980
rect 23388 12928 23440 12980
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 6828 12860 6880 12912
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 7012 12792 7064 12844
rect 9312 12792 9364 12844
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 12532 12792 12584 12844
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 14648 12835 14700 12844
rect 14648 12801 14657 12835
rect 14657 12801 14691 12835
rect 14691 12801 14700 12835
rect 14648 12792 14700 12801
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 1584 12724 1636 12776
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 3332 12724 3384 12776
rect 4528 12724 4580 12776
rect 5724 12724 5776 12776
rect 6368 12724 6420 12776
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 12164 12724 12216 12776
rect 13820 12724 13872 12776
rect 18144 12724 18196 12776
rect 20812 12724 20864 12776
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 7288 12699 7340 12708
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2596 12588 2648 12640
rect 2964 12588 3016 12640
rect 7288 12665 7297 12699
rect 7297 12665 7331 12699
rect 7331 12665 7340 12699
rect 7288 12656 7340 12665
rect 14372 12699 14424 12708
rect 14372 12665 14381 12699
rect 14381 12665 14415 12699
rect 14415 12665 14424 12699
rect 14372 12656 14424 12665
rect 16212 12656 16264 12708
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7196 12631 7248 12640
rect 7196 12597 7205 12631
rect 7205 12597 7239 12631
rect 7239 12597 7248 12631
rect 7196 12588 7248 12597
rect 7840 12631 7892 12640
rect 7840 12597 7849 12631
rect 7849 12597 7883 12631
rect 7883 12597 7892 12631
rect 7840 12588 7892 12597
rect 15568 12588 15620 12640
rect 15936 12588 15988 12640
rect 16488 12588 16540 12640
rect 17960 12588 18012 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3240 12427 3292 12436
rect 3240 12393 3249 12427
rect 3249 12393 3283 12427
rect 3283 12393 3292 12427
rect 3240 12384 3292 12393
rect 2780 12316 2832 12368
rect 3976 12384 4028 12436
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 4344 12384 4396 12436
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 9312 12427 9364 12436
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 11704 12384 11756 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 13084 12384 13136 12436
rect 13452 12384 13504 12436
rect 16396 12427 16448 12436
rect 5540 12316 5592 12368
rect 5816 12316 5868 12368
rect 8576 12316 8628 12368
rect 10140 12359 10192 12368
rect 10140 12325 10149 12359
rect 10149 12325 10183 12359
rect 10183 12325 10192 12359
rect 10140 12316 10192 12325
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 22744 12384 22796 12436
rect 16672 12316 16724 12368
rect 17132 12316 17184 12368
rect 2136 12291 2188 12300
rect 2136 12257 2145 12291
rect 2145 12257 2179 12291
rect 2179 12257 2188 12291
rect 2136 12248 2188 12257
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 2688 12248 2740 12300
rect 4160 12248 4212 12300
rect 5264 12291 5316 12300
rect 5264 12257 5273 12291
rect 5273 12257 5307 12291
rect 5307 12257 5316 12291
rect 5264 12248 5316 12257
rect 6460 12248 6512 12300
rect 8208 12248 8260 12300
rect 9956 12248 10008 12300
rect 11520 12248 11572 12300
rect 13084 12248 13136 12300
rect 15476 12248 15528 12300
rect 21732 12291 21784 12300
rect 21732 12257 21741 12291
rect 21741 12257 21775 12291
rect 21775 12257 21784 12291
rect 21732 12248 21784 12257
rect 2596 12180 2648 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 2044 12112 2096 12164
rect 7748 12155 7800 12164
rect 7748 12121 7757 12155
rect 7757 12121 7791 12155
rect 7791 12121 7800 12155
rect 7748 12112 7800 12121
rect 9680 12112 9732 12164
rect 10784 12180 10836 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12716 12180 12768 12232
rect 13820 12180 13872 12232
rect 14648 12180 14700 12232
rect 15292 12180 15344 12232
rect 15936 12180 15988 12232
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 17960 12112 18012 12164
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 7564 12044 7616 12096
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 15476 12087 15528 12096
rect 15476 12053 15485 12087
rect 15485 12053 15519 12087
rect 15519 12053 15528 12087
rect 15476 12044 15528 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11840 1636 11892
rect 4160 11840 4212 11892
rect 5172 11883 5224 11892
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 5172 11840 5224 11849
rect 6184 11840 6236 11892
rect 6460 11840 6512 11892
rect 7104 11772 7156 11824
rect 5540 11704 5592 11756
rect 7564 11704 7616 11756
rect 10140 11840 10192 11892
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 11796 11840 11848 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 16488 11840 16540 11892
rect 16672 11840 16724 11892
rect 17868 11840 17920 11892
rect 18052 11883 18104 11892
rect 18052 11849 18061 11883
rect 18061 11849 18095 11883
rect 18095 11849 18104 11883
rect 18052 11840 18104 11849
rect 16304 11704 16356 11756
rect 17132 11704 17184 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 2780 11636 2832 11688
rect 8576 11636 8628 11688
rect 13360 11636 13412 11688
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 2964 11568 3016 11620
rect 3700 11568 3752 11620
rect 6552 11611 6604 11620
rect 6552 11577 6561 11611
rect 6561 11577 6595 11611
rect 6595 11577 6604 11611
rect 6552 11568 6604 11577
rect 9680 11568 9732 11620
rect 9956 11568 10008 11620
rect 11060 11568 11112 11620
rect 11520 11568 11572 11620
rect 13544 11611 13596 11620
rect 13544 11577 13578 11611
rect 13578 11577 13596 11611
rect 13544 11568 13596 11577
rect 16580 11568 16632 11620
rect 2044 11500 2096 11552
rect 5448 11500 5500 11552
rect 6736 11500 6788 11552
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 11336 11543 11388 11552
rect 11336 11509 11345 11543
rect 11345 11509 11379 11543
rect 11379 11509 11388 11543
rect 11336 11500 11388 11509
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 14648 11543 14700 11552
rect 14648 11509 14657 11543
rect 14657 11509 14691 11543
rect 14691 11509 14700 11543
rect 14648 11500 14700 11509
rect 15568 11500 15620 11552
rect 17132 11500 17184 11552
rect 21732 11543 21784 11552
rect 21732 11509 21741 11543
rect 21741 11509 21775 11543
rect 21775 11509 21784 11543
rect 21732 11500 21784 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1860 11296 1912 11348
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 2228 11296 2280 11348
rect 3332 11296 3384 11348
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 8208 11339 8260 11348
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 11796 11296 11848 11348
rect 13360 11339 13412 11348
rect 13360 11305 13369 11339
rect 13369 11305 13403 11339
rect 13403 11305 13412 11339
rect 13360 11296 13412 11305
rect 16212 11296 16264 11348
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 5264 11228 5316 11280
rect 6828 11228 6880 11280
rect 8392 11228 8444 11280
rect 11244 11228 11296 11280
rect 11336 11228 11388 11280
rect 13268 11228 13320 11280
rect 19984 11296 20036 11348
rect 18604 11228 18656 11280
rect 2780 11160 2832 11169
rect 4160 11160 4212 11212
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 6184 11203 6236 11212
rect 4528 11160 4580 11169
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 14648 11160 14700 11212
rect 15844 11160 15896 11212
rect 17776 11203 17828 11212
rect 17776 11169 17785 11203
rect 17785 11169 17819 11203
rect 17819 11169 17828 11203
rect 17776 11160 17828 11169
rect 4620 11135 4672 11144
rect 2596 11024 2648 11076
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 10508 11092 10560 11144
rect 13728 11092 13780 11144
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 15292 11135 15344 11144
rect 13912 11092 13964 11101
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 4068 11067 4120 11076
rect 4068 11033 4077 11067
rect 4077 11033 4111 11067
rect 4111 11033 4120 11067
rect 4068 11024 4120 11033
rect 5540 11024 5592 11076
rect 10784 11024 10836 11076
rect 13544 11024 13596 11076
rect 3148 10956 3200 11008
rect 7564 10999 7616 11008
rect 7564 10965 7573 10999
rect 7573 10965 7607 10999
rect 7607 10965 7616 10999
rect 7564 10956 7616 10965
rect 12440 10956 12492 11008
rect 17132 10956 17184 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3332 10752 3384 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 6828 10752 6880 10804
rect 8576 10752 8628 10804
rect 2964 10548 3016 10600
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 5172 10548 5224 10600
rect 10508 10752 10560 10804
rect 11244 10752 11296 10804
rect 13912 10752 13964 10804
rect 15752 10752 15804 10804
rect 15844 10752 15896 10804
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 19248 10752 19300 10804
rect 15292 10684 15344 10736
rect 15752 10659 15804 10668
rect 15752 10625 15761 10659
rect 15761 10625 15795 10659
rect 15795 10625 15804 10659
rect 15752 10616 15804 10625
rect 9864 10548 9916 10600
rect 15660 10548 15712 10600
rect 16764 10591 16816 10600
rect 16764 10557 16773 10591
rect 16773 10557 16807 10591
rect 16807 10557 16816 10591
rect 16764 10548 16816 10557
rect 18236 10548 18288 10600
rect 2044 10480 2096 10532
rect 2596 10480 2648 10532
rect 2228 10412 2280 10464
rect 2412 10412 2464 10464
rect 4896 10480 4948 10532
rect 7564 10523 7616 10532
rect 7564 10489 7598 10523
rect 7598 10489 7616 10523
rect 7564 10480 7616 10489
rect 8668 10480 8720 10532
rect 9496 10480 9548 10532
rect 12440 10480 12492 10532
rect 16488 10480 16540 10532
rect 3976 10412 4028 10464
rect 15660 10455 15712 10464
rect 15660 10421 15669 10455
rect 15669 10421 15703 10455
rect 15703 10421 15712 10455
rect 15660 10412 15712 10421
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 2780 10208 2832 10260
rect 3884 10251 3936 10260
rect 3884 10217 3893 10251
rect 3893 10217 3927 10251
rect 3927 10217 3936 10251
rect 3884 10208 3936 10217
rect 4620 10251 4672 10260
rect 4620 10217 4629 10251
rect 4629 10217 4663 10251
rect 4663 10217 4672 10251
rect 4620 10208 4672 10217
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 8668 10251 8720 10260
rect 8668 10217 8677 10251
rect 8677 10217 8711 10251
rect 8711 10217 8720 10251
rect 8668 10208 8720 10217
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 10876 10208 10928 10260
rect 11244 10208 11296 10260
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 13820 10208 13872 10260
rect 17132 10251 17184 10260
rect 17132 10217 17141 10251
rect 17141 10217 17175 10251
rect 17175 10217 17184 10251
rect 17132 10208 17184 10217
rect 17316 10208 17368 10260
rect 3516 10183 3568 10192
rect 3516 10149 3525 10183
rect 3525 10149 3559 10183
rect 3559 10149 3568 10183
rect 3516 10140 3568 10149
rect 3976 10140 4028 10192
rect 5356 10140 5408 10192
rect 2780 10115 2832 10124
rect 2780 10081 2789 10115
rect 2789 10081 2823 10115
rect 2823 10081 2832 10115
rect 2780 10072 2832 10081
rect 5172 10115 5224 10124
rect 5172 10081 5181 10115
rect 5181 10081 5215 10115
rect 5215 10081 5224 10115
rect 5172 10072 5224 10081
rect 6000 10072 6052 10124
rect 6184 10072 6236 10124
rect 7472 10072 7524 10124
rect 9404 10072 9456 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3148 10004 3200 10056
rect 3516 10004 3568 10056
rect 8116 10047 8168 10056
rect 7656 9979 7708 9988
rect 7656 9945 7665 9979
rect 7665 9945 7699 9979
rect 7699 9945 7708 9979
rect 7656 9936 7708 9945
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8024 9936 8076 9988
rect 9680 10004 9732 10056
rect 15752 10140 15804 10192
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 13820 10115 13872 10124
rect 11704 10072 11756 10081
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 18144 10072 18196 10124
rect 11796 10047 11848 10056
rect 9956 9936 10008 9988
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 12440 10004 12492 10056
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 15292 10004 15344 10056
rect 10416 9936 10468 9988
rect 13728 9936 13780 9988
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 9588 9868 9640 9920
rect 9680 9868 9732 9920
rect 10692 9868 10744 9920
rect 12992 9868 13044 9920
rect 15752 9868 15804 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2780 9707 2832 9716
rect 2780 9673 2789 9707
rect 2789 9673 2823 9707
rect 2823 9673 2832 9707
rect 3516 9707 3568 9716
rect 2780 9664 2832 9673
rect 3516 9673 3525 9707
rect 3525 9673 3559 9707
rect 3559 9673 3568 9707
rect 3516 9664 3568 9673
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 2136 9596 2188 9648
rect 2412 9639 2464 9648
rect 2412 9605 2421 9639
rect 2421 9605 2455 9639
rect 2455 9605 2464 9639
rect 2412 9596 2464 9605
rect 2504 9596 2556 9648
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 4988 9596 5040 9648
rect 7564 9639 7616 9648
rect 7564 9605 7573 9639
rect 7573 9605 7607 9639
rect 7607 9605 7616 9639
rect 7564 9596 7616 9605
rect 9588 9664 9640 9716
rect 1400 9460 1452 9512
rect 1860 9460 1912 9512
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 5448 9528 5500 9580
rect 5540 9528 5592 9580
rect 10416 9664 10468 9716
rect 11244 9707 11296 9716
rect 11244 9673 11253 9707
rect 11253 9673 11287 9707
rect 11287 9673 11296 9707
rect 11244 9664 11296 9673
rect 11704 9664 11756 9716
rect 12072 9664 12124 9716
rect 12256 9664 12308 9716
rect 13912 9707 13964 9716
rect 13912 9673 13921 9707
rect 13921 9673 13955 9707
rect 13955 9673 13964 9707
rect 13912 9664 13964 9673
rect 15292 9664 15344 9716
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 12164 9596 12216 9648
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9588 9528 9640 9580
rect 10692 9528 10744 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 18144 9596 18196 9648
rect 16580 9528 16632 9580
rect 4252 9503 4304 9512
rect 4252 9469 4275 9503
rect 4275 9469 4304 9503
rect 18052 9503 18104 9512
rect 4252 9460 4304 9469
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 14096 9392 14148 9444
rect 1768 9324 1820 9376
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 6644 9324 6696 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 9680 9324 9732 9376
rect 11612 9324 11664 9376
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12900 9367 12952 9376
rect 12440 9324 12492 9333
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 13728 9324 13780 9376
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1676 9120 1728 9172
rect 1860 9120 1912 9172
rect 2044 9120 2096 9172
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 4068 9120 4120 9172
rect 4252 9163 4304 9172
rect 4252 9129 4261 9163
rect 4261 9129 4295 9163
rect 4295 9129 4304 9163
rect 4252 9120 4304 9129
rect 4528 9120 4580 9172
rect 5448 9120 5500 9172
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 11796 9120 11848 9172
rect 12900 9120 12952 9172
rect 12992 9120 13044 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 15752 9163 15804 9172
rect 15752 9129 15761 9163
rect 15761 9129 15795 9163
rect 15795 9129 15804 9163
rect 15752 9120 15804 9129
rect 17776 9120 17828 9172
rect 2688 9052 2740 9104
rect 6552 9052 6604 9104
rect 8668 9095 8720 9104
rect 8668 9061 8677 9095
rect 8677 9061 8711 9095
rect 8711 9061 8720 9095
rect 8668 9052 8720 9061
rect 9864 9052 9916 9104
rect 16396 9052 16448 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 2596 8984 2648 9036
rect 5356 8984 5408 9036
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 7380 8984 7432 9036
rect 10232 8984 10284 9036
rect 11888 8984 11940 9036
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 12164 8959 12216 8968
rect 12164 8925 12173 8959
rect 12173 8925 12207 8959
rect 12207 8925 12216 8959
rect 12164 8916 12216 8925
rect 2688 8891 2740 8900
rect 2688 8857 2697 8891
rect 2697 8857 2731 8891
rect 2731 8857 2740 8891
rect 2688 8848 2740 8857
rect 5080 8891 5132 8900
rect 5080 8857 5089 8891
rect 5089 8857 5123 8891
rect 5123 8857 5132 8891
rect 5080 8848 5132 8857
rect 10692 8780 10744 8832
rect 11704 8780 11756 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2320 8576 2372 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 10048 8576 10100 8628
rect 5356 8508 5408 8560
rect 9864 8508 9916 8560
rect 11704 8576 11756 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 12164 8576 12216 8628
rect 7472 8440 7524 8492
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 2596 8415 2648 8424
rect 2596 8381 2605 8415
rect 2605 8381 2639 8415
rect 2639 8381 2648 8415
rect 2596 8372 2648 8381
rect 8024 8372 8076 8424
rect 11888 8440 11940 8492
rect 14096 8576 14148 8628
rect 16580 8619 16632 8628
rect 16580 8585 16589 8619
rect 16589 8585 16623 8619
rect 16623 8585 16632 8619
rect 16580 8576 16632 8585
rect 12992 8372 13044 8424
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 10232 8304 10284 8356
rect 12164 8347 12216 8356
rect 12164 8313 12173 8347
rect 12173 8313 12207 8347
rect 12207 8313 12216 8347
rect 12164 8304 12216 8313
rect 7472 8236 7524 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 8032 1452 8084
rect 1492 8032 1544 8084
rect 2136 8032 2188 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 11888 8032 11940 8084
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 1676 7896 1728 7948
rect 2228 7896 2280 7948
rect 10140 7896 10192 7948
rect 10600 7939 10652 7948
rect 10600 7905 10634 7939
rect 10634 7905 10652 7939
rect 10600 7896 10652 7905
rect 572 7760 624 7812
rect 9404 7760 9456 7812
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1676 7531 1728 7540
rect 1676 7497 1685 7531
rect 1685 7497 1719 7531
rect 1719 7497 1728 7531
rect 1676 7488 1728 7497
rect 10140 7488 10192 7540
rect 10600 7488 10652 7540
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 10784 5312 10836 5364
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 9496 5083 9548 5092
rect 9496 5049 9530 5083
rect 9530 5049 9548 5083
rect 9496 5040 9548 5049
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 4620 4428 4672 4480
rect 7472 4428 7524 4480
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 2778 27704 2834 27713
rect 2778 27639 2834 27648
rect 308 27418 336 27520
rect 216 27390 336 27418
rect 216 14929 244 27390
rect 202 14920 258 14929
rect 202 14855 258 14864
rect 860 13530 888 27520
rect 1412 25514 1440 27520
rect 1412 25486 1900 25514
rect 1768 25356 1820 25362
rect 1768 25298 1820 25304
rect 1400 25220 1452 25226
rect 1400 25162 1452 25168
rect 1412 24750 1440 25162
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1490 23624 1546 23633
rect 1490 23559 1546 23568
rect 1504 22794 1532 23559
rect 1596 23225 1624 25094
rect 1780 24954 1808 25298
rect 1768 24948 1820 24954
rect 1768 24890 1820 24896
rect 1768 24676 1820 24682
rect 1768 24618 1820 24624
rect 1582 23216 1638 23225
rect 1582 23151 1638 23160
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1412 22766 1532 22794
rect 1412 21010 1440 22766
rect 1582 22536 1638 22545
rect 1688 22506 1716 22918
rect 1582 22471 1638 22480
rect 1676 22500 1728 22506
rect 1492 22432 1544 22438
rect 1492 22374 1544 22380
rect 1504 21078 1532 22374
rect 1596 21690 1624 22471
rect 1676 22442 1728 22448
rect 1688 22234 1716 22442
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1582 21448 1638 21457
rect 1582 21383 1638 21392
rect 1596 21146 1624 21383
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1492 21072 1544 21078
rect 1492 21014 1544 21020
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 20602 1440 20946
rect 1400 20596 1452 20602
rect 1400 20538 1452 20544
rect 1676 19984 1728 19990
rect 1676 19926 1728 19932
rect 1582 19680 1638 19689
rect 1582 19615 1638 19624
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 18086 1440 18770
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 16794 1440 18022
rect 1490 17912 1546 17921
rect 1490 17847 1546 17856
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1504 15162 1532 17847
rect 1596 17338 1624 19615
rect 1688 18970 1716 19926
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1688 18426 1716 18906
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1674 17504 1730 17513
rect 1674 17439 1730 17448
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1688 15994 1716 17439
rect 1780 16561 1808 24618
rect 1872 21350 1900 25486
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 1964 21162 1992 27520
rect 2136 25424 2188 25430
rect 2136 25366 2188 25372
rect 2042 24712 2098 24721
rect 2042 24647 2098 24656
rect 2056 21690 2084 24647
rect 2148 23254 2176 25366
rect 2320 25356 2372 25362
rect 2320 25298 2372 25304
rect 2332 24886 2360 25298
rect 2412 25152 2464 25158
rect 2412 25094 2464 25100
rect 2320 24880 2372 24886
rect 2318 24848 2320 24857
rect 2372 24848 2374 24857
rect 2424 24818 2452 25094
rect 2318 24783 2374 24792
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2320 24608 2372 24614
rect 2320 24550 2372 24556
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 2136 23248 2188 23254
rect 2136 23190 2188 23196
rect 2136 22976 2188 22982
rect 2136 22918 2188 22924
rect 2148 22234 2176 22918
rect 2136 22228 2188 22234
rect 2136 22170 2188 22176
rect 2240 22030 2268 24006
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 2044 21684 2096 21690
rect 2044 21626 2096 21632
rect 2056 21486 2084 21626
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 2044 21344 2096 21350
rect 2044 21286 2096 21292
rect 1872 21134 1992 21162
rect 1766 16552 1822 16561
rect 1766 16487 1822 16496
rect 1596 15966 1716 15994
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13705 1440 14350
rect 1596 14074 1624 15966
rect 1676 15904 1728 15910
rect 1674 15872 1676 15881
rect 1728 15872 1730 15881
rect 1674 15807 1730 15816
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 14890 1716 15302
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1674 14648 1730 14657
rect 1780 14618 1808 15506
rect 1872 15337 1900 21134
rect 1952 21072 2004 21078
rect 1952 21014 2004 21020
rect 1964 20466 1992 21014
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 1964 20330 1992 20402
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1964 19990 1992 20266
rect 1952 19984 2004 19990
rect 1952 19926 2004 19932
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1964 18630 1992 19110
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 2056 17814 2084 21286
rect 2044 17808 2096 17814
rect 2044 17750 2096 17756
rect 2044 17604 2096 17610
rect 2044 17546 2096 17552
rect 2056 17338 2084 17546
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2148 17218 2176 21830
rect 2240 21146 2268 21966
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2240 20398 2268 20742
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2240 20058 2268 20334
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2332 19394 2360 24550
rect 2424 23866 2452 24754
rect 2516 24750 2544 27520
rect 2792 25430 2820 27639
rect 3146 27520 3202 28000
rect 3698 27520 3754 28000
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 2870 26616 2926 26625
rect 2870 26551 2926 26560
rect 2780 25424 2832 25430
rect 2780 25366 2832 25372
rect 2596 25220 2648 25226
rect 2596 25162 2648 25168
rect 2504 24744 2556 24750
rect 2504 24686 2556 24692
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2516 24410 2544 24550
rect 2504 24404 2556 24410
rect 2504 24346 2556 24352
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2424 23594 2452 23802
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 2608 23338 2636 25162
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2424 23310 2636 23338
rect 2424 22250 2452 23310
rect 2504 23248 2556 23254
rect 2504 23190 2556 23196
rect 2516 22778 2544 23190
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2516 22420 2544 22714
rect 2700 22506 2728 23462
rect 2688 22500 2740 22506
rect 2688 22442 2740 22448
rect 2596 22432 2648 22438
rect 2516 22392 2596 22420
rect 2596 22374 2648 22380
rect 2424 22222 2636 22250
rect 2608 20618 2636 22222
rect 2688 22024 2740 22030
rect 2792 22001 2820 25094
rect 2884 24750 2912 26551
rect 3054 25392 3110 25401
rect 3054 25327 3056 25336
rect 3108 25327 3110 25336
rect 3056 25298 3108 25304
rect 2872 24744 2924 24750
rect 2872 24686 2924 24692
rect 2884 24342 2912 24686
rect 3068 24614 3096 25298
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 2872 24336 2924 24342
rect 2872 24278 2924 24284
rect 3068 24274 3096 24550
rect 3056 24268 3108 24274
rect 3056 24210 3108 24216
rect 2872 24200 2924 24206
rect 2872 24142 2924 24148
rect 2884 23526 2912 24142
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 2872 23520 2924 23526
rect 2872 23462 2924 23468
rect 2884 23322 2912 23462
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2884 23050 2912 23258
rect 2872 23044 2924 23050
rect 2872 22986 2924 22992
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2688 21966 2740 21972
rect 2778 21992 2834 22001
rect 2700 21706 2728 21966
rect 2778 21927 2834 21936
rect 2884 21706 2912 22374
rect 2700 21690 2912 21706
rect 2688 21684 2912 21690
rect 2740 21678 2912 21684
rect 2688 21626 2740 21632
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2686 20904 2742 20913
rect 2686 20839 2688 20848
rect 2740 20839 2742 20848
rect 2688 20810 2740 20816
rect 2608 20590 2728 20618
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2608 19514 2636 19994
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2332 19366 2636 19394
rect 2412 19236 2464 19242
rect 2412 19178 2464 19184
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2240 17882 2268 18702
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2332 17746 2360 18702
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2240 17338 2268 17614
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2148 17190 2360 17218
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2042 16144 2098 16153
rect 2240 16114 2268 16390
rect 2042 16079 2098 16088
rect 2228 16108 2280 16114
rect 2056 16046 2084 16079
rect 2228 16050 2280 16056
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2134 16008 2190 16017
rect 2134 15943 2136 15952
rect 2188 15943 2190 15952
rect 2136 15914 2188 15920
rect 1858 15328 1914 15337
rect 1858 15263 1914 15272
rect 2148 14618 2176 15914
rect 1674 14583 1730 14592
rect 1768 14612 1820 14618
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 848 13524 900 13530
rect 848 13466 900 13472
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12782 1624 13126
rect 1584 12776 1636 12782
rect 1504 12724 1584 12730
rect 1504 12718 1636 12724
rect 1504 12702 1624 12718
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9518 1440 9998
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1398 9344 1454 9353
rect 1398 9279 1454 9288
rect 1412 9042 1440 9279
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 8090 1440 8978
rect 1504 8090 1532 12702
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1596 8634 1624 11834
rect 1688 9178 1716 14583
rect 1768 14554 1820 14560
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2240 14498 2268 16050
rect 2148 14470 2268 14498
rect 1858 13560 1914 13569
rect 1858 13495 1914 13504
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 10713 1808 12038
rect 1872 11354 1900 13495
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1964 13190 1992 13330
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12186 1992 13126
rect 2148 12782 2176 14470
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2240 12306 2268 13126
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 1964 12170 2084 12186
rect 1964 12164 2096 12170
rect 1964 12158 2044 12164
rect 2044 12106 2096 12112
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11354 1992 11630
rect 2056 11558 2084 12106
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1766 10704 1822 10713
rect 1766 10639 1822 10648
rect 1858 10568 1914 10577
rect 2056 10538 2084 11494
rect 1858 10503 1914 10512
rect 2044 10532 2096 10538
rect 1872 10266 1900 10503
rect 2044 10474 2096 10480
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1872 9874 1900 10202
rect 1780 9846 1900 9874
rect 1780 9382 1808 9846
rect 2056 9586 2084 10474
rect 2148 9654 2176 12242
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2240 11257 2268 11290
rect 2226 11248 2282 11257
rect 2226 11183 2282 11192
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1872 9178 1900 9454
rect 2056 9178 2084 9522
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2148 8090 2176 9590
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2240 7954 2268 10406
rect 2332 8634 2360 17190
rect 2424 16538 2452 19178
rect 2502 19136 2558 19145
rect 2502 19071 2558 19080
rect 2516 17270 2544 19071
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2424 16510 2544 16538
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2424 14521 2452 16390
rect 2410 14512 2466 14521
rect 2410 14447 2466 14456
rect 2516 14362 2544 16510
rect 2424 14334 2544 14362
rect 2424 10470 2452 14334
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 13938 2544 14214
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2410 10296 2466 10305
rect 2410 10231 2412 10240
rect 2464 10231 2466 10240
rect 2412 10202 2464 10208
rect 2410 10024 2466 10033
rect 2410 9959 2466 9968
rect 2424 9654 2452 9959
rect 2516 9654 2544 13874
rect 2608 13818 2636 19366
rect 2700 19145 2728 20590
rect 2686 19136 2742 19145
rect 2686 19071 2742 19080
rect 2884 18630 2912 21286
rect 2976 20602 3004 23530
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 3068 22098 3096 23122
rect 3056 22092 3108 22098
rect 3056 22034 3108 22040
rect 3160 21298 3188 27520
rect 3424 25424 3476 25430
rect 3424 25366 3476 25372
rect 3238 23760 3294 23769
rect 3238 23695 3294 23704
rect 3252 21894 3280 23695
rect 3330 23352 3386 23361
rect 3330 23287 3386 23296
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3068 21270 3188 21298
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2976 19514 3004 19858
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 2976 18970 3004 19450
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 2976 18766 3004 18906
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2688 18624 2740 18630
rect 2872 18624 2924 18630
rect 2740 18584 2820 18612
rect 2688 18566 2740 18572
rect 2792 17882 2820 18584
rect 2872 18566 2924 18572
rect 2884 18329 2912 18566
rect 2976 18426 3004 18702
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 2870 18320 2926 18329
rect 2870 18255 2926 18264
rect 2884 18222 2912 18255
rect 2872 18216 2924 18222
rect 2924 18164 3004 18170
rect 2872 18158 3004 18164
rect 2884 18142 3004 18158
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2976 17678 3004 18142
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2792 17270 2820 17614
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 3068 17082 3096 21270
rect 3146 21176 3202 21185
rect 3146 21111 3202 21120
rect 3160 21010 3188 21111
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3252 20058 3280 21286
rect 3344 20369 3372 23287
rect 3436 23186 3464 25366
rect 3712 24834 3740 27520
rect 3882 27160 3938 27169
rect 3882 27095 3938 27104
rect 3620 24806 3740 24834
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3528 24313 3556 24686
rect 3514 24304 3570 24313
rect 3514 24239 3570 24248
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3436 21418 3464 21830
rect 3424 21412 3476 21418
rect 3424 21354 3476 21360
rect 3330 20360 3386 20369
rect 3330 20295 3386 20304
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19514 3188 19654
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3160 19310 3188 19450
rect 3252 19378 3280 19994
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 18970 3556 19246
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3514 17640 3570 17649
rect 3514 17575 3570 17584
rect 3528 17338 3556 17575
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3528 17134 3556 17274
rect 2976 17054 3096 17082
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 2686 16960 2742 16969
rect 2686 16895 2742 16904
rect 2700 16794 2728 16895
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2686 16552 2742 16561
rect 2686 16487 2742 16496
rect 2700 15978 2728 16487
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2792 15910 2820 16594
rect 2976 16561 3004 17054
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2962 16552 3018 16561
rect 2962 16487 3018 16496
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2792 15042 2820 15846
rect 2884 15706 2912 16050
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2792 15014 2912 15042
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2700 14618 2728 14894
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2608 13790 2820 13818
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13462 2636 13670
rect 2792 13546 2820 13790
rect 2700 13518 2820 13546
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2608 13297 2636 13398
rect 2594 13288 2650 13297
rect 2594 13223 2650 13232
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2608 12646 2636 12786
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2700 12481 2728 13518
rect 2686 12472 2742 12481
rect 2686 12407 2742 12416
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11082 2636 12174
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2608 10538 2636 11018
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2700 9110 2728 12242
rect 2792 11694 2820 12310
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10266 2820 11154
rect 2884 11121 2912 15014
rect 2976 13938 3004 16487
rect 3068 16266 3096 16934
rect 3068 16250 3188 16266
rect 3068 16244 3200 16250
rect 3068 16238 3148 16244
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 11626 3004 12582
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2870 11112 2926 11121
rect 2870 11047 2926 11056
rect 2976 10606 3004 11562
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2792 9722 2820 10066
rect 2872 10056 2924 10062
rect 2870 10024 2872 10033
rect 2924 10024 2926 10033
rect 2870 9959 2926 9968
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2962 9616 3018 9625
rect 2962 9551 3018 9560
rect 2976 9518 3004 9551
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2976 9178 3004 9454
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2608 8430 2636 8978
rect 2686 8936 2742 8945
rect 2686 8871 2688 8880
rect 2740 8871 2742 8880
rect 2688 8842 2740 8848
rect 2596 8424 2648 8430
rect 2594 8392 2596 8401
rect 2648 8392 2650 8401
rect 2594 8327 2650 8336
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 572 7812 624 7818
rect 572 7754 624 7760
rect 584 4321 612 7754
rect 1688 7546 1716 7890
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 570 4312 626 4321
rect 570 4247 626 4256
rect 2686 3224 2742 3233
rect 2742 3182 2820 3210
rect 2686 3159 2742 3168
rect 2792 2961 2820 3182
rect 2778 2952 2834 2961
rect 2778 2887 2834 2896
rect 938 2544 994 2553
rect 938 2479 994 2488
rect 952 1737 980 2479
rect 938 1728 994 1737
rect 938 1663 994 1672
rect 3068 377 3096 16238
rect 3148 16186 3200 16192
rect 3620 16046 3648 24806
rect 3698 24440 3754 24449
rect 3698 24375 3754 24384
rect 3712 21554 3740 24375
rect 3792 24336 3844 24342
rect 3792 24278 3844 24284
rect 3804 23497 3832 24278
rect 3896 23866 3924 27095
rect 4066 26072 4122 26081
rect 4122 26030 4200 26058
rect 4066 26007 4122 26016
rect 4172 24698 4200 26030
rect 4264 24834 4292 27520
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4264 24806 4568 24834
rect 4172 24670 4292 24698
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 4066 24576 4122 24585
rect 3988 24410 4016 24550
rect 4066 24511 4122 24520
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 3790 23488 3846 23497
rect 3790 23423 3846 23432
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3988 21010 4016 22374
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3804 16153 3832 20742
rect 3988 20602 4016 20742
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3988 20330 4016 20538
rect 4080 20330 4108 24511
rect 4264 22001 4292 24670
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4448 24313 4476 24550
rect 4434 24304 4490 24313
rect 4434 24239 4490 24248
rect 4436 24200 4488 24206
rect 4436 24142 4488 24148
rect 4448 23526 4476 24142
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4448 23186 4476 23462
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4250 21992 4306 22001
rect 4250 21927 4306 21936
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4448 19378 4476 20198
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4066 19272 4122 19281
rect 4066 19207 4122 19216
rect 4080 18834 4108 19207
rect 4344 19168 4396 19174
rect 4158 19136 4214 19145
rect 4344 19110 4396 19116
rect 4158 19071 4214 19080
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 3882 17912 3938 17921
rect 4080 17882 4108 18770
rect 3882 17847 3884 17856
rect 3936 17847 3938 17856
rect 4068 17876 4120 17882
rect 3884 17818 3936 17824
rect 4068 17818 4120 17824
rect 3896 17202 3924 17818
rect 4172 17338 4200 19071
rect 4252 18624 4304 18630
rect 4250 18592 4252 18601
rect 4304 18592 4306 18601
rect 4250 18527 4306 18536
rect 4356 18426 4384 19110
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4436 17808 4488 17814
rect 4436 17750 4488 17756
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3790 16144 3846 16153
rect 3896 16114 3924 16390
rect 4342 16144 4398 16153
rect 3790 16079 3846 16088
rect 3884 16108 3936 16114
rect 4342 16079 4398 16088
rect 3884 16050 3936 16056
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3160 14958 3188 15098
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3344 14550 3372 15846
rect 3620 15706 3648 15982
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3620 14657 3648 15642
rect 3606 14648 3662 14657
rect 3606 14583 3662 14592
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3160 13530 3188 14350
rect 3252 14346 3280 14418
rect 3712 14385 3740 15846
rect 3896 15366 3924 16050
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4250 15600 4306 15609
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3896 14958 3924 15302
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3698 14376 3754 14385
rect 3240 14340 3292 14346
rect 3698 14311 3754 14320
rect 3240 14282 3292 14288
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3252 12442 3280 14282
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 13938 3464 14214
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3436 12968 3464 13874
rect 3516 12980 3568 12986
rect 3436 12940 3516 12968
rect 3516 12922 3568 12928
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3606 12744 3662 12753
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3344 11354 3372 12718
rect 3606 12679 3662 12688
rect 3422 11656 3478 11665
rect 3422 11591 3478 11600
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10062 3188 10950
rect 3344 10810 3372 11290
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3436 4865 3464 11591
rect 3514 11384 3570 11393
rect 3514 11319 3516 11328
rect 3568 11319 3570 11328
rect 3516 11290 3568 11296
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3528 10062 3556 10134
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3528 9722 3556 9998
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3620 6089 3648 12679
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3606 6080 3662 6089
rect 3606 6015 3662 6024
rect 3712 5409 3740 11562
rect 3804 11354 3832 14486
rect 3896 13530 3924 14894
rect 4172 13818 4200 15574
rect 4250 15535 4306 15544
rect 4264 15337 4292 15535
rect 4250 15328 4306 15337
rect 4250 15263 4306 15272
rect 4080 13802 4200 13818
rect 4068 13796 4200 13802
rect 4120 13790 4200 13796
rect 4068 13738 4120 13744
rect 4264 13530 4292 15263
rect 4356 14074 4384 16079
rect 4448 14618 4476 17750
rect 4540 15638 4568 24806
rect 4632 24070 4660 25162
rect 4724 24342 4752 25230
rect 4816 24449 4844 27520
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 5092 24954 5120 25230
rect 5368 24954 5396 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 5356 24948 5408 24954
rect 5356 24890 5408 24896
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 5000 24449 5028 24686
rect 5540 24608 5592 24614
rect 6012 24585 6040 27520
rect 6092 25152 6144 25158
rect 6092 25094 6144 25100
rect 5540 24550 5592 24556
rect 5998 24576 6054 24585
rect 4802 24440 4858 24449
rect 4802 24375 4858 24384
rect 4986 24440 5042 24449
rect 4986 24375 5042 24384
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4632 23746 4660 24006
rect 4724 23866 4752 24278
rect 4988 24268 5040 24274
rect 4988 24210 5040 24216
rect 5000 24177 5028 24210
rect 4986 24168 5042 24177
rect 4986 24103 5042 24112
rect 5446 24168 5502 24177
rect 5446 24103 5502 24112
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4632 23718 4752 23746
rect 4724 23186 4752 23718
rect 5000 23322 5028 24103
rect 5354 23760 5410 23769
rect 5460 23730 5488 24103
rect 5354 23695 5356 23704
rect 5408 23695 5410 23704
rect 5448 23724 5500 23730
rect 5356 23666 5408 23672
rect 5448 23666 5500 23672
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4724 22234 4752 23122
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22234 5212 22374
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 4802 21992 4858 22001
rect 4802 21927 4858 21936
rect 4816 20398 4844 21927
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 20913 5028 21830
rect 5276 21434 5304 23598
rect 5552 23361 5580 24550
rect 5998 24511 6054 24520
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5538 23352 5594 23361
rect 5538 23287 5594 23296
rect 5998 23080 6054 23089
rect 5998 23015 6054 23024
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5354 22536 5410 22545
rect 6012 22506 6040 23015
rect 5354 22471 5410 22480
rect 6000 22500 6052 22506
rect 5368 22166 5396 22471
rect 6000 22442 6052 22448
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5368 21690 5396 22102
rect 5998 21856 6054 21865
rect 5622 21788 5918 21808
rect 5998 21791 6054 21800
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5276 21406 5396 21434
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 4986 20904 5042 20913
rect 4986 20839 5042 20848
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4816 20058 4844 20334
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4816 19514 4844 19994
rect 4908 19718 4936 20402
rect 5092 19786 5120 20742
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4632 16130 4660 17682
rect 4724 17134 4752 18022
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16794 4752 17070
rect 4816 16998 4844 19110
rect 4908 18329 4936 19654
rect 5092 18612 5120 19722
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19310 5212 19654
rect 5276 19310 5304 21286
rect 5368 19496 5396 21406
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5552 21049 5580 21286
rect 5538 21040 5594 21049
rect 5538 20975 5594 20984
rect 5448 20936 5500 20942
rect 5500 20884 5580 20890
rect 5448 20878 5580 20884
rect 5460 20862 5580 20878
rect 5736 20874 5764 21490
rect 6012 21486 6040 21791
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 5552 20602 5580 20862
rect 5724 20868 5776 20874
rect 5724 20810 5776 20816
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6104 20602 6132 25094
rect 6182 24848 6238 24857
rect 6182 24783 6184 24792
rect 6236 24783 6238 24792
rect 6184 24754 6236 24760
rect 6564 24721 6592 27520
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6550 24712 6606 24721
rect 6550 24647 6606 24656
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6564 23526 6592 24210
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 6644 23588 6696 23594
rect 6644 23530 6696 23536
rect 6552 23520 6604 23526
rect 6550 23488 6552 23497
rect 6604 23488 6606 23497
rect 6550 23423 6606 23432
rect 6656 23186 6684 23530
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6288 22642 6316 22918
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6288 22438 6316 22578
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 5446 20360 5502 20369
rect 5446 20295 5448 20304
rect 5500 20295 5502 20304
rect 5448 20266 5500 20272
rect 5460 20058 5488 20266
rect 5448 20052 5500 20058
rect 5500 20012 5580 20040
rect 5448 19994 5500 20000
rect 5368 19468 5488 19496
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5276 18970 5304 19246
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5368 18902 5396 19314
rect 5356 18896 5408 18902
rect 5356 18838 5408 18844
rect 5172 18624 5224 18630
rect 5092 18584 5172 18612
rect 5172 18566 5224 18572
rect 4894 18320 4950 18329
rect 4894 18255 4950 18264
rect 5080 18216 5132 18222
rect 5078 18184 5080 18193
rect 5132 18184 5134 18193
rect 4988 18148 5040 18154
rect 5078 18119 5134 18128
rect 4988 18090 5040 18096
rect 5000 17066 5028 18090
rect 5184 17814 5212 18566
rect 5368 18290 5396 18838
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4816 16726 4844 16934
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4632 16102 4752 16130
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4632 15706 4660 15982
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4724 15570 4752 16102
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4526 14920 4582 14929
rect 4526 14855 4582 14864
rect 4540 14618 4568 14855
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4448 14074 4476 14554
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4540 14006 4568 14554
rect 4632 14414 4660 15302
rect 4724 15162 4752 15506
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4724 14890 4752 15098
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4908 14550 4936 16662
rect 5000 16658 5028 17002
rect 5368 16998 5396 17682
rect 5460 17270 5488 19468
rect 5552 19310 5580 20012
rect 6196 19990 6224 21966
rect 6288 21078 6316 22374
rect 6564 21690 6592 22510
rect 6748 22030 6776 23462
rect 6840 23322 6868 23598
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6458 20768 6514 20777
rect 6458 20703 6514 20712
rect 6184 19984 6236 19990
rect 6184 19926 6236 19932
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6196 19310 6224 19926
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5552 18222 5580 18838
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5552 17882 5580 18158
rect 6104 17882 6132 18226
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 5552 17338 5580 17818
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5078 16824 5134 16833
rect 5078 16759 5134 16768
rect 5092 16658 5120 16759
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5092 16250 5120 16594
rect 5368 16590 5396 16934
rect 5460 16794 5488 17206
rect 6472 16969 6500 20703
rect 6552 16992 6604 16998
rect 6182 16960 6238 16969
rect 6182 16895 6238 16904
rect 6458 16960 6514 16969
rect 6552 16934 6604 16940
rect 6458 16895 6514 16904
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 5276 16114 5304 16390
rect 5368 16250 5396 16526
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5460 16182 5488 16730
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5172 15904 5224 15910
rect 5170 15872 5172 15881
rect 5224 15872 5226 15881
rect 5170 15807 5226 15816
rect 5276 15570 5304 16050
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4896 14544 4948 14550
rect 4802 14512 4858 14521
rect 4896 14486 4948 14492
rect 4802 14447 4858 14456
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4264 13410 4292 13466
rect 4264 13382 4384 13410
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3896 10266 3924 13126
rect 3988 12986 4016 13194
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3988 12442 4016 12922
rect 4250 12880 4306 12889
rect 4250 12815 4306 12824
rect 4066 12608 4122 12617
rect 4066 12543 4122 12552
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4080 12322 4108 12543
rect 4264 12442 4292 12815
rect 4356 12442 4384 13382
rect 4540 12986 4568 13942
rect 4816 13870 4844 14447
rect 5000 14278 5028 15030
rect 5276 14822 5304 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5276 14618 5304 14758
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5460 14278 5488 14894
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5000 13938 5028 14214
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4804 13864 4856 13870
rect 4802 13832 4804 13841
rect 4856 13832 4858 13841
rect 4802 13767 4858 13776
rect 4712 13728 4764 13734
rect 4710 13696 4712 13705
rect 4764 13696 4766 13705
rect 4710 13631 4766 13640
rect 4724 13530 4752 13631
rect 5460 13569 5488 14214
rect 5552 13977 5580 14758
rect 6012 14521 6040 15846
rect 6196 14634 6224 16895
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6274 16552 6330 16561
rect 6274 16487 6330 16496
rect 6288 16250 6316 16487
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6380 15026 6408 16594
rect 6564 16522 6592 16934
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 16046 6500 16390
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6564 15162 6592 16458
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6196 14606 6316 14634
rect 5998 14512 6054 14521
rect 5998 14447 6054 14456
rect 6092 14476 6144 14482
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5538 13968 5594 13977
rect 5538 13903 5594 13912
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5446 13560 5502 13569
rect 4712 13524 4764 13530
rect 5446 13495 5502 13504
rect 4712 13466 4764 13472
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4540 12782 4568 12922
rect 4632 12918 4660 13398
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 5092 12356 5120 12854
rect 5552 12374 5580 13670
rect 6012 13530 6040 14447
rect 6144 14436 6224 14464
rect 6092 14418 6144 14424
rect 6196 14074 6224 14436
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6288 13818 6316 14606
rect 6380 14278 6408 14962
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6368 14068 6420 14074
rect 6472 14056 6500 14894
rect 6564 14550 6592 15098
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6564 14074 6592 14486
rect 6420 14028 6500 14056
rect 6368 14010 6420 14016
rect 6288 13790 6408 13818
rect 6274 13696 6330 13705
rect 6274 13631 6330 13640
rect 6288 13530 6316 13631
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6184 13320 6236 13326
rect 5998 13288 6054 13297
rect 6184 13262 6236 13268
rect 5998 13223 6054 13232
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5814 12880 5870 12889
rect 5814 12815 5816 12824
rect 5868 12815 5870 12824
rect 5816 12786 5868 12792
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 3988 12294 4108 12322
rect 5000 12328 5120 12356
rect 5540 12368 5592 12374
rect 5262 12336 5318 12345
rect 4160 12300 4212 12306
rect 3988 11801 4016 12294
rect 4160 12242 4212 12248
rect 4172 11898 4200 12242
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 4526 11248 4582 11257
rect 4160 11212 4212 11218
rect 4526 11183 4528 11192
rect 4160 11154 4212 11160
rect 4580 11183 4582 11192
rect 4528 11154 4580 11160
rect 4066 11112 4122 11121
rect 4066 11047 4068 11056
rect 4120 11047 4122 11056
rect 4068 11018 4120 11024
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3988 10198 4016 10406
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4080 10044 4108 10542
rect 4172 10305 4200 11154
rect 4158 10296 4214 10305
rect 4158 10231 4214 10240
rect 3988 10016 4108 10044
rect 3988 9518 4016 10016
rect 4172 9738 4200 10231
rect 4080 9710 4200 9738
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4080 9178 4108 9710
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4264 9178 4292 9454
rect 4540 9178 4568 11154
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4632 10266 4660 11086
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4908 10266 4936 10474
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 5000 9654 5028 12328
rect 5736 12345 5764 12718
rect 5828 12374 5856 12786
rect 5816 12368 5868 12374
rect 5540 12310 5592 12316
rect 5722 12336 5778 12345
rect 5262 12271 5264 12280
rect 5316 12271 5318 12280
rect 5264 12242 5316 12248
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 5184 11898 5212 12135
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5276 11286 5304 12242
rect 5552 11762 5580 12310
rect 5816 12310 5868 12316
rect 5722 12271 5778 12280
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 5460 11064 5488 11494
rect 5552 11354 5580 11698
rect 6012 11354 6040 13223
rect 6196 12646 6224 13262
rect 6288 12986 6316 13466
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6380 12782 6408 13790
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6184 12640 6236 12646
rect 6182 12608 6184 12617
rect 6236 12608 6238 12617
rect 6182 12543 6238 12552
rect 6380 12345 6408 12718
rect 6366 12336 6422 12345
rect 6472 12306 6500 14028
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6564 13326 6592 14010
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6550 13016 6606 13025
rect 6550 12951 6606 12960
rect 6564 12753 6592 12951
rect 6550 12744 6606 12753
rect 6550 12679 6606 12688
rect 6366 12271 6422 12280
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6472 11898 6500 12242
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6196 11218 6224 11834
rect 6550 11656 6606 11665
rect 6550 11591 6552 11600
rect 6604 11591 6606 11600
rect 6552 11562 6604 11568
rect 6656 11393 6684 21830
rect 6748 21146 6776 21966
rect 6840 21690 6868 22170
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6932 21486 6960 25230
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 7024 23322 7052 23666
rect 7116 23633 7144 27520
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7392 24614 7420 24754
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7392 24138 7420 24550
rect 7380 24132 7432 24138
rect 7380 24074 7432 24080
rect 7102 23624 7158 23633
rect 7102 23559 7158 23568
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 7024 22506 7052 23258
rect 7392 23186 7420 24074
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 23662 7512 24006
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7116 22778 7144 23122
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7392 22642 7420 23122
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7576 22234 7604 22442
rect 7564 22228 7616 22234
rect 7484 22188 7564 22216
rect 7484 21554 7512 22188
rect 7564 22170 7616 22176
rect 7562 22128 7618 22137
rect 7562 22063 7618 22072
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6748 20262 6776 20742
rect 6932 20602 6960 21014
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6748 19922 6776 20198
rect 6736 19916 6788 19922
rect 6788 19876 6868 19904
rect 6736 19858 6788 19864
rect 6840 19174 6868 19876
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18222 6868 19110
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6932 18154 6960 18566
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6932 17542 6960 18090
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17202 6960 17478
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7024 16726 7052 20198
rect 7576 19174 7604 22063
rect 7668 21185 7696 27520
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 7852 24614 7880 25094
rect 8220 24857 8248 27520
rect 8206 24848 8262 24857
rect 8206 24783 8262 24792
rect 8206 24712 8262 24721
rect 8206 24647 8208 24656
rect 8260 24647 8262 24656
rect 8208 24618 8260 24624
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7760 24410 7788 24550
rect 7852 24426 7880 24550
rect 7930 24440 7986 24449
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7852 24398 7930 24426
rect 7760 23662 7788 24346
rect 7748 23656 7800 23662
rect 7748 23598 7800 23604
rect 7852 22137 7880 24398
rect 7930 24375 7986 24384
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 8128 24041 8156 24278
rect 8114 24032 8170 24041
rect 8114 23967 8170 23976
rect 8128 23866 8156 23967
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8864 23361 8892 27520
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9232 23866 9260 24210
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 7930 23352 7986 23361
rect 7930 23287 7986 23296
rect 8850 23352 8906 23361
rect 8850 23287 8906 23296
rect 7838 22128 7894 22137
rect 7838 22063 7894 22072
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7852 21690 7880 21966
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7654 21176 7710 21185
rect 7654 21111 7710 21120
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7484 18902 7512 19110
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7576 18766 7604 19110
rect 7668 18970 7696 20810
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7852 19990 7880 20742
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7944 19310 7972 23287
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 8036 21350 8064 22714
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 8036 20330 8064 21286
rect 8128 20874 8156 22034
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 8114 20632 8170 20641
rect 8114 20567 8170 20576
rect 8128 20398 8156 20567
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8024 20324 8076 20330
rect 8024 20266 8076 20272
rect 8128 20058 8156 20334
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 8114 18864 8170 18873
rect 7656 18828 7708 18834
rect 8114 18799 8116 18808
rect 7656 18770 7708 18776
rect 8168 18799 8170 18808
rect 8116 18770 8168 18776
rect 7564 18760 7616 18766
rect 7562 18728 7564 18737
rect 7616 18728 7618 18737
rect 7562 18663 7618 18672
rect 7562 18592 7618 18601
rect 7562 18527 7618 18536
rect 7576 17338 7604 18527
rect 7668 17882 7696 18770
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 8128 17814 8156 18770
rect 8220 18426 8248 22510
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 9048 22234 9076 22374
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 8680 22030 8708 22170
rect 8668 22024 8720 22030
rect 8668 21966 8720 21972
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8116 17808 8168 17814
rect 8022 17776 8078 17785
rect 8116 17750 8168 17756
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8022 17711 8024 17720
rect 8076 17711 8078 17720
rect 8024 17682 8076 17688
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7930 17232 7986 17241
rect 7930 17167 7986 17176
rect 7944 17134 7972 17167
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16833 7420 16934
rect 7378 16824 7434 16833
rect 7944 16794 7972 17070
rect 7378 16759 7434 16768
rect 7932 16788 7984 16794
rect 7392 16726 7420 16759
rect 7932 16730 7984 16736
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6840 16182 6868 16594
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6932 15706 6960 16526
rect 7010 16416 7066 16425
rect 7010 16351 7066 16360
rect 7024 15910 7052 16351
rect 7392 16250 7420 16662
rect 8036 16658 8064 17682
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8128 16726 8156 17614
rect 8220 17134 8248 17750
rect 8312 17678 8340 19994
rect 8300 17672 8352 17678
rect 8404 17649 8432 21830
rect 8680 21486 8708 21966
rect 8668 21480 8720 21486
rect 9416 21457 9444 27520
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9692 23866 9720 24346
rect 9784 24342 9812 24686
rect 9772 24336 9824 24342
rect 9968 24290 9996 27520
rect 10520 25786 10548 27520
rect 10520 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10048 24676 10100 24682
rect 10048 24618 10100 24624
rect 9772 24278 9824 24284
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9784 23662 9812 24278
rect 9876 24262 9996 24290
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9508 23322 9536 23598
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 8668 21422 8720 21428
rect 9402 21448 9458 21457
rect 9508 21418 9536 23258
rect 9692 23186 9720 23462
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9692 22778 9720 23122
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9784 22522 9812 23190
rect 9876 23089 9904 24262
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9968 23594 9996 24142
rect 10060 23866 10088 24618
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9862 23080 9918 23089
rect 10060 23066 10088 23802
rect 10152 23254 10180 24006
rect 10704 23769 10732 25758
rect 10966 24848 11022 24857
rect 10966 24783 11022 24792
rect 10690 23760 10746 23769
rect 10690 23695 10746 23704
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 10140 23112 10192 23118
rect 10060 23060 10140 23066
rect 10060 23054 10192 23060
rect 10060 23038 10180 23054
rect 9862 23015 9918 23024
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 9692 22494 9812 22522
rect 9692 22216 9720 22494
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 22234 9812 22374
rect 9600 22188 9720 22216
rect 9772 22228 9824 22234
rect 9600 22098 9628 22188
rect 9772 22170 9824 22176
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9402 21383 9458 21392
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 21146 9996 21286
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8588 20641 8616 20742
rect 8574 20632 8630 20641
rect 8574 20567 8630 20576
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 8956 18222 8984 19246
rect 9232 19242 9260 20198
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9232 18970 9260 19178
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9232 18766 9260 18906
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9232 18358 9260 18702
rect 9324 18426 9352 19654
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8300 17614 8352 17620
rect 8390 17640 8446 17649
rect 8312 17270 8340 17614
rect 8390 17575 8446 17584
rect 8956 17270 8984 18158
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 9416 17134 9444 20470
rect 9692 19786 9720 20946
rect 9968 20534 9996 21082
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 9784 19666 9812 20198
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9692 19638 9812 19666
rect 9692 19496 9720 19638
rect 9508 19468 9720 19496
rect 9772 19508 9824 19514
rect 9508 17814 9536 19468
rect 9772 19450 9824 19456
rect 9678 19408 9734 19417
rect 9678 19343 9734 19352
rect 9692 18222 9720 19343
rect 9784 19009 9812 19450
rect 9876 19394 9904 19858
rect 10060 19514 10088 22918
rect 10152 22778 10180 23038
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10796 22642 10824 22918
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22098 10732 22510
rect 10796 22234 10824 22578
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10784 21956 10836 21962
rect 10784 21898 10836 21904
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10796 21146 10824 21898
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10690 21040 10746 21049
rect 10690 20975 10746 20984
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 10152 20040 10180 20742
rect 10704 20330 10732 20975
rect 10782 20496 10838 20505
rect 10782 20431 10784 20440
rect 10836 20431 10838 20440
rect 10784 20402 10836 20408
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20266
rect 10692 20052 10744 20058
rect 10152 20012 10272 20040
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9876 19366 9996 19394
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9770 19000 9826 19009
rect 9770 18935 9826 18944
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9784 18290 9812 18838
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 18034 9720 18158
rect 9600 18006 9720 18034
rect 9600 17882 9628 18006
rect 9876 17921 9904 19178
rect 9968 18630 9996 19366
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 9956 18624 10008 18630
rect 9954 18592 9956 18601
rect 10008 18592 10010 18601
rect 9954 18527 10010 18536
rect 9862 17912 9918 17921
rect 9588 17876 9640 17882
rect 9862 17847 9918 17856
rect 9588 17818 9640 17824
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17241 9720 17478
rect 9678 17232 9734 17241
rect 9678 17167 9734 17176
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9416 16794 9444 17070
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 7562 16280 7618 16289
rect 7380 16244 7432 16250
rect 7562 16215 7618 16224
rect 7380 16186 7432 16192
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7024 15638 7052 15846
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7300 14278 7328 15438
rect 7392 15337 7420 16050
rect 7576 15745 7604 16215
rect 8404 16114 8432 16594
rect 9416 16590 9444 16730
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9416 16250 9444 16526
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 7562 15736 7618 15745
rect 7562 15671 7618 15680
rect 7562 15600 7618 15609
rect 7562 15535 7564 15544
rect 7616 15535 7618 15544
rect 7564 15506 7616 15512
rect 7852 15502 7880 16050
rect 8404 15706 8432 16050
rect 8956 15706 8984 16118
rect 9494 16008 9550 16017
rect 9220 15972 9272 15978
rect 9494 15943 9550 15952
rect 9220 15914 9272 15920
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7378 15328 7434 15337
rect 7378 15263 7434 15272
rect 7852 15201 7880 15438
rect 7838 15192 7894 15201
rect 8312 15162 8340 15506
rect 9232 15366 9260 15914
rect 9508 15910 9536 15943
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 7838 15127 7894 15136
rect 8300 15156 8352 15162
rect 7852 14958 7880 15127
rect 8300 15098 8352 15104
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8390 14512 8446 14521
rect 8390 14447 8392 14456
rect 8444 14447 8446 14456
rect 8392 14418 8444 14424
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6932 13954 6960 14010
rect 6840 13926 6960 13954
rect 6840 12918 6868 13926
rect 7300 13462 7328 14214
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 7024 12850 7052 13126
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6826 12744 6882 12753
rect 6826 12679 6882 12688
rect 6840 12646 6868 12679
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6828 12436 6880 12442
rect 7024 12424 7052 12786
rect 6880 12396 7052 12424
rect 6828 12378 6880 12384
rect 6736 11552 6788 11558
rect 6734 11520 6736 11529
rect 6788 11520 6790 11529
rect 6734 11455 6790 11464
rect 6642 11384 6698 11393
rect 6642 11319 6698 11328
rect 6840 11286 6868 12378
rect 7116 11830 7144 13398
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12714 7328 13126
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7208 12209 7236 12582
rect 7194 12200 7250 12209
rect 7194 12135 7250 12144
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 5540 11076 5592 11082
rect 5460 11036 5540 11064
rect 5540 11018 5592 11024
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10130 5212 10542
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5368 9722 5396 10134
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5552 9586 5580 11018
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6196 10810 6224 11154
rect 6840 10810 6868 11222
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6196 10130 6224 10746
rect 7484 10418 7512 13806
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7576 13569 7604 13670
rect 7562 13560 7618 13569
rect 8128 13530 8156 13874
rect 8300 13864 8352 13870
rect 8298 13832 8300 13841
rect 8352 13832 8354 13841
rect 8298 13767 8354 13776
rect 8588 13705 8616 14350
rect 8956 14074 8984 14826
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8574 13696 8630 13705
rect 8574 13631 8630 13640
rect 7562 13495 7618 13504
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7668 13433 7696 13466
rect 7654 13424 7710 13433
rect 7654 13359 7710 13368
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 7852 12646 7880 13330
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12481 7880 12582
rect 7838 12472 7894 12481
rect 7838 12407 7894 12416
rect 8588 12374 8616 13262
rect 8772 12986 8800 13330
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7746 12200 7802 12209
rect 7746 12135 7748 12144
rect 7800 12135 7802 12144
rect 7748 12106 7800 12112
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7576 11762 7604 12038
rect 7944 11801 7972 12038
rect 7930 11792 7986 11801
rect 7564 11756 7616 11762
rect 7930 11727 7986 11736
rect 7564 11698 7616 11704
rect 7576 11014 7604 11698
rect 8220 11354 8248 12242
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8404 11529 8432 12174
rect 8588 11694 8616 12174
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8390 11520 8446 11529
rect 8390 11455 8446 11464
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8404 11286 8432 11455
rect 8588 11354 8616 11630
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10538 7604 10950
rect 8588 10810 8616 11290
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 7484 10390 7604 10418
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5354 9480 5410 9489
rect 5354 9415 5410 9424
rect 4894 9208 4950 9217
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4528 9172 4580 9178
rect 4894 9143 4950 9152
rect 4528 9114 4580 9120
rect 4908 8945 4936 9143
rect 5368 9042 5396 9415
rect 5460 9178 5488 9522
rect 6012 9382 6040 10066
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 4894 8936 4950 8945
rect 4894 8871 4950 8880
rect 5078 8936 5134 8945
rect 5078 8871 5080 8880
rect 5132 8871 5134 8880
rect 5080 8842 5132 8848
rect 5368 8566 5396 8978
rect 5460 8634 5488 9114
rect 6564 9110 6592 9862
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6564 8634 6592 9046
rect 6656 9042 6684 9318
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 7392 8378 7420 8978
rect 7484 8498 7512 10066
rect 7576 9654 7604 10390
rect 8680 10266 8708 10474
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8116 10056 8168 10062
rect 7654 10024 7710 10033
rect 8116 9998 8168 10004
rect 7654 9959 7656 9968
rect 7708 9959 7710 9968
rect 8024 9988 8076 9994
rect 7656 9930 7708 9936
rect 8024 9930 8076 9936
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 9081 7880 9318
rect 8036 9178 8064 9930
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7838 9072 7894 9081
rect 7838 9007 7894 9016
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 8036 8430 8064 9114
rect 8128 8945 8156 9998
rect 9048 9761 9076 15098
rect 9232 12986 9260 15302
rect 9692 15065 9720 16730
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9784 15881 9812 16594
rect 10060 16561 10088 19314
rect 10046 16552 10102 16561
rect 10046 16487 10102 16496
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 15910 9996 16390
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9956 15904 10008 15910
rect 9770 15872 9826 15881
rect 9956 15846 10008 15852
rect 9770 15807 9826 15816
rect 9678 15056 9734 15065
rect 9678 14991 9734 15000
rect 9770 14512 9826 14521
rect 9770 14447 9826 14456
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13802 9628 14282
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 13190 9628 13738
rect 9692 13394 9720 14214
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9324 12442 9352 12786
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9600 12322 9628 13126
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12442 9720 12718
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9600 12294 9720 12322
rect 9692 12170 9720 12294
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9508 10266 9536 10474
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9034 9752 9090 9761
rect 9034 9687 9090 9696
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8680 9110 8708 9522
rect 9416 9382 9444 10066
rect 9692 10062 9720 11562
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9600 9722 9628 9862
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9600 9586 9628 9658
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9586 9480 9642 9489
rect 9692 9466 9720 9862
rect 9784 9625 9812 14447
rect 9968 13530 9996 15846
rect 10060 15638 10088 16050
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 14890 10088 15302
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10046 14648 10102 14657
rect 10046 14583 10048 14592
rect 10100 14583 10102 14592
rect 10048 14554 10100 14560
rect 10060 14074 10088 14554
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10152 13954 10180 19654
rect 10244 19242 10272 20012
rect 10692 19994 10744 20000
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10796 19378 10824 19654
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10796 18834 10824 19110
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10704 18086 10732 18566
rect 10796 18426 10824 18770
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17746 10732 18022
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10796 17338 10824 17750
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10704 15910 10732 16526
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15609 10732 15846
rect 10888 15722 10916 22442
rect 10980 22030 11008 24783
rect 11072 24410 11100 27520
rect 11716 24857 11744 27520
rect 11702 24848 11758 24857
rect 12268 24818 12296 27520
rect 11702 24783 11758 24792
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 11164 24177 11192 24550
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11150 24168 11206 24177
rect 11150 24103 11206 24112
rect 11348 23866 11376 24210
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11624 23594 11652 24210
rect 11808 24041 11836 24550
rect 12162 24168 12218 24177
rect 12162 24103 12218 24112
rect 11794 24032 11850 24041
rect 11794 23967 11850 23976
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 11612 23588 11664 23594
rect 11612 23530 11664 23536
rect 11072 22642 11100 23530
rect 11716 23186 11744 23802
rect 12070 23488 12126 23497
rect 12070 23423 12126 23432
rect 12084 23254 12112 23423
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11716 22778 11744 23122
rect 12084 22778 12112 23190
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 11992 22438 12020 22714
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 10968 22024 11020 22030
rect 11072 22001 11100 22034
rect 10968 21966 11020 21972
rect 11058 21992 11114 22001
rect 10980 21622 11008 21966
rect 11058 21927 11114 21936
rect 11072 21690 11100 21927
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11348 21146 11376 21286
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20602 11100 20878
rect 11348 20602 11376 21082
rect 11808 20942 11836 21490
rect 11992 20942 12020 22374
rect 12084 22030 12112 22714
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11072 19174 11100 19858
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18290 11100 19110
rect 11256 18970 11284 19790
rect 11440 19514 11468 19790
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10980 16810 11008 18158
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17105 11100 18022
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11058 17096 11114 17105
rect 11058 17031 11114 17040
rect 11164 16998 11192 17682
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11426 16824 11482 16833
rect 10980 16782 11192 16810
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16153 11008 16390
rect 10966 16144 11022 16153
rect 10966 16079 11022 16088
rect 10968 15904 11020 15910
rect 10966 15872 10968 15881
rect 11020 15872 11022 15881
rect 10966 15807 11022 15816
rect 10796 15694 10916 15722
rect 10690 15600 10746 15609
rect 10690 15535 10746 15544
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 14958 10364 15438
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14385 10364 14418
rect 10322 14376 10378 14385
rect 10322 14311 10378 14320
rect 10336 14006 10364 14311
rect 10060 13926 10180 13954
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9968 11626 9996 12242
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 10606 9904 11494
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 10060 10441 10088 13926
rect 10704 13734 10732 14826
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10138 13560 10194 13569
rect 10289 13552 10585 13572
rect 10138 13495 10140 13504
rect 10192 13495 10194 13504
rect 10140 13466 10192 13472
rect 10152 12986 10180 13466
rect 10704 13326 10732 13670
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10244 12850 10272 13262
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12368 10192 12374
rect 10138 12336 10140 12345
rect 10192 12336 10194 12345
rect 10796 12322 10824 15694
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10888 15162 10916 15574
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10888 14618 10916 15098
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10138 12271 10194 12280
rect 10704 12294 10824 12322
rect 10152 11898 10180 12271
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10520 10810 10548 11086
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10046 10432 10102 10441
rect 10046 10367 10102 10376
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9862 10160 9918 10169
rect 10322 10160 10378 10169
rect 9918 10104 10180 10112
rect 9862 10095 10180 10104
rect 10322 10095 10378 10104
rect 9876 10084 10180 10095
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9862 9888 9918 9897
rect 9862 9823 9918 9832
rect 9770 9616 9826 9625
rect 9770 9551 9826 9560
rect 9692 9438 9812 9466
rect 9586 9415 9642 9424
rect 9600 9382 9628 9415
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8944 8968 8996 8974
rect 8114 8936 8170 8945
rect 8114 8871 8170 8880
rect 8942 8936 8944 8945
rect 8996 8936 8998 8945
rect 8942 8871 8998 8880
rect 8024 8424 8076 8430
rect 7392 8350 7512 8378
rect 8024 8366 8076 8372
rect 7484 8294 7512 8350
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 3974 7848 4030 7857
rect 3974 7783 4030 7792
rect 3698 5400 3754 5409
rect 3698 5335 3754 5344
rect 3422 4856 3478 4865
rect 3422 4791 3478 4800
rect 3988 3777 4016 7783
rect 4080 7177 4108 7919
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 7484 4486 7512 8230
rect 8036 8090 8064 8366
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 9416 7818 9444 9318
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9692 7410 9720 9318
rect 9784 8401 9812 9438
rect 9876 9217 9904 9823
rect 9862 9208 9918 9217
rect 9862 9143 9918 9152
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9876 8566 9904 9046
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9770 8392 9826 8401
rect 9770 8327 9826 8336
rect 9876 8090 9904 8502
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9232 4486 9260 5102
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 3974 3768 4030 3777
rect 3974 3703 4030 3712
rect 4632 480 4660 4422
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 9508 4049 9536 5034
rect 9494 4040 9550 4049
rect 9494 3975 9550 3984
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 9968 1329 9996 9930
rect 10152 9738 10180 10084
rect 10230 9752 10286 9761
rect 10060 9710 10230 9738
rect 10060 8634 10088 9710
rect 10230 9687 10286 9696
rect 10336 9364 10364 10095
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10428 9722 10456 9930
rect 10704 9926 10732 12294
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11082 10824 12174
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 11506 11100 11562
rect 10980 11478 11100 11506
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10152 9353 10364 9364
rect 10138 9344 10364 9353
rect 10194 9336 10364 9344
rect 10138 9279 10194 9288
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10244 8378 10272 8978
rect 10704 8838 10732 9522
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10598 8528 10654 8537
rect 10598 8463 10600 8472
rect 10652 8463 10654 8472
rect 10600 8434 10652 8440
rect 10152 8362 10272 8378
rect 10152 8356 10284 8362
rect 10152 8350 10232 8356
rect 10152 7954 10180 8350
rect 10232 8298 10284 8304
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7970 10732 8774
rect 10612 7954 10732 7970
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10600 7948 10732 7954
rect 10652 7942 10732 7948
rect 10600 7890 10652 7896
rect 10152 7546 10180 7890
rect 10612 7546 10640 7890
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10796 5370 10824 11018
rect 10876 10260 10928 10266
rect 10980 10248 11008 11478
rect 10928 10220 11008 10248
rect 10876 10202 10928 10208
rect 11164 9897 11192 16782
rect 11426 16759 11428 16768
rect 11480 16759 11482 16768
rect 11428 16730 11480 16736
rect 11716 16697 11744 20742
rect 11808 20058 11836 20878
rect 11992 20602 12020 20878
rect 12176 20777 12204 24103
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12360 23304 12388 23530
rect 12440 23316 12492 23322
rect 12360 23276 12440 23304
rect 12440 23258 12492 23264
rect 12438 22536 12494 22545
rect 12438 22471 12440 22480
rect 12492 22471 12494 22480
rect 12440 22442 12492 22448
rect 12636 22030 12664 24550
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12728 22234 12756 23462
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12268 21690 12296 21898
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12636 21622 12664 21966
rect 12728 21690 12756 22170
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 20942 12756 21286
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 12162 20768 12218 20777
rect 12162 20703 12218 20712
rect 12360 20618 12388 20810
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12360 20602 12480 20618
rect 11980 20596 12032 20602
rect 12360 20596 12492 20602
rect 12360 20590 12440 20596
rect 11980 20538 12032 20544
rect 12440 20538 12492 20544
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11992 19922 12020 20538
rect 12544 20398 12572 20742
rect 12820 20534 12848 27520
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13096 24818 13124 25094
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13096 22438 13124 24754
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13084 21072 13136 21078
rect 13084 21014 13136 21020
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 13096 20466 13124 21014
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 12532 20392 12584 20398
rect 12530 20360 12532 20369
rect 12584 20360 12586 20369
rect 12530 20295 12586 20304
rect 13096 20058 13124 20402
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12360 19292 12388 19858
rect 12636 19514 12664 19858
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12532 19304 12584 19310
rect 12360 19264 12532 19292
rect 12532 19246 12584 19252
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11808 18306 11836 18566
rect 12268 18426 12296 18634
rect 12544 18630 12572 19246
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 18698 12756 19178
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 11888 18352 11940 18358
rect 11808 18300 11888 18306
rect 11808 18294 11940 18300
rect 11808 18278 11928 18294
rect 11702 16688 11758 16697
rect 11702 16623 11758 16632
rect 11610 16416 11666 16425
rect 11610 16351 11666 16360
rect 11624 16250 11652 16351
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11624 15978 11652 16186
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15473 11284 15846
rect 11242 15464 11298 15473
rect 11242 15399 11298 15408
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11716 15201 11744 15302
rect 11702 15192 11758 15201
rect 11702 15127 11758 15136
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11440 13841 11468 14010
rect 11426 13832 11482 13841
rect 11426 13767 11482 13776
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11532 12986 11560 13330
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11256 12345 11284 12378
rect 11242 12336 11298 12345
rect 11242 12271 11298 12280
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11256 11286 11284 11834
rect 11532 11626 11560 12242
rect 11716 11778 11744 12378
rect 11808 12322 11836 18278
rect 12268 17882 12296 18362
rect 13188 17921 13216 21830
rect 13372 18986 13400 27520
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13556 22574 13584 23462
rect 13832 22982 13860 23530
rect 13820 22976 13872 22982
rect 13820 22918 13872 22924
rect 13832 22778 13860 22918
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 13728 22024 13780 22030
rect 13832 22012 13860 22714
rect 13780 21984 13860 22012
rect 13728 21966 13780 21972
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13556 21418 13584 21830
rect 13818 21448 13874 21457
rect 13544 21412 13596 21418
rect 13818 21383 13874 21392
rect 13544 21354 13596 21360
rect 13832 20602 13860 21383
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13832 20398 13860 20538
rect 13924 20505 13952 27520
rect 14568 24857 14596 27520
rect 15120 25242 15148 27520
rect 14752 25214 15148 25242
rect 14554 24848 14610 24857
rect 14554 24783 14610 24792
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14568 21690 14596 22442
rect 14752 21865 14780 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15672 24664 15700 27520
rect 15396 24636 15700 24664
rect 15396 24313 15424 24636
rect 15658 24576 15714 24585
rect 15658 24511 15714 24520
rect 15672 24410 15700 24511
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15382 24304 15438 24313
rect 15382 24239 15438 24248
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15488 23526 15516 24210
rect 15108 23520 15160 23526
rect 15106 23488 15108 23497
rect 15476 23520 15528 23526
rect 15160 23488 15162 23497
rect 15476 23462 15528 23468
rect 15106 23423 15162 23432
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14738 21856 14794 21865
rect 14738 21791 14794 21800
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14108 21146 14136 21354
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14094 20904 14150 20913
rect 14094 20839 14150 20848
rect 14278 20904 14334 20913
rect 14278 20839 14334 20848
rect 13910 20496 13966 20505
rect 13910 20431 13966 20440
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 13280 18970 13400 18986
rect 13280 18964 13412 18970
rect 13280 18958 13360 18964
rect 13280 18358 13308 18958
rect 13360 18906 13412 18912
rect 14016 18873 14044 20198
rect 14108 19310 14136 20839
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14002 18864 14058 18873
rect 13360 18828 13412 18834
rect 14002 18799 14058 18808
rect 13360 18770 13412 18776
rect 13372 18737 13400 18770
rect 13358 18728 13414 18737
rect 13358 18663 13414 18672
rect 13372 18426 13400 18663
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13648 18222 13676 18566
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13450 18048 13506 18057
rect 13450 17983 13506 17992
rect 13174 17912 13230 17921
rect 12256 17876 12308 17882
rect 13464 17882 13492 17983
rect 13174 17847 13230 17856
rect 13452 17876 13504 17882
rect 12256 17818 12308 17824
rect 13452 17818 13504 17824
rect 13082 17640 13138 17649
rect 13082 17575 13084 17584
rect 13136 17575 13138 17584
rect 13084 17546 13136 17552
rect 12992 17536 13044 17542
rect 13044 17484 13124 17490
rect 12992 17478 13124 17484
rect 13004 17462 13124 17478
rect 13096 17066 13124 17462
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13096 16969 13124 17002
rect 13082 16960 13138 16969
rect 13082 16895 13138 16904
rect 13096 16658 13124 16895
rect 13464 16726 13492 17818
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13556 16794 13584 17614
rect 13648 16998 13676 18158
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13832 17898 13860 18090
rect 13740 17870 13860 17898
rect 13740 17678 13768 17870
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13740 17338 13768 17614
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 14292 16794 14320 20839
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14554 20632 14610 20641
rect 14956 20624 15252 20644
rect 14554 20567 14610 20576
rect 14568 20466 14596 20567
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19417 15332 19790
rect 15290 19408 15346 19417
rect 15290 19343 15346 19352
rect 15106 19272 15162 19281
rect 15106 19207 15162 19216
rect 15120 19174 15148 19207
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14924 18352 14976 18358
rect 14922 18320 14924 18329
rect 14976 18320 14978 18329
rect 14922 18255 14978 18264
rect 15304 18057 15332 18702
rect 15290 18048 15346 18057
rect 15290 17983 15346 17992
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 15396 16726 15424 17614
rect 15488 16794 15516 23462
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15580 22438 15608 23122
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12268 15910 12296 16594
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 12070 14784 12126 14793
rect 11900 14482 11928 14758
rect 12070 14719 12126 14728
rect 12084 14550 12112 14719
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11900 13734 11928 14418
rect 12084 14074 12112 14486
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13326 11928 13670
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 12986 11928 13262
rect 12162 13016 12218 13025
rect 11888 12980 11940 12986
rect 12162 12951 12164 12960
rect 11888 12922 11940 12928
rect 12216 12951 12218 12960
rect 12164 12922 12216 12928
rect 12176 12782 12204 12922
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11808 12294 12020 12322
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11898 11836 12174
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11716 11750 11836 11778
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11808 11558 11836 11750
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11348 11286 11376 11494
rect 11808 11354 11836 11494
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11256 10810 11284 11222
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11256 10266 11284 10746
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11150 9888 11206 9897
rect 11150 9823 11206 9832
rect 11242 9752 11298 9761
rect 11242 9687 11244 9696
rect 11296 9687 11298 9696
rect 11244 9658 11296 9664
rect 11624 9382 11652 10066
rect 11716 9722 11744 10066
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 7857 11652 9318
rect 11808 9178 11836 9998
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11716 8634 11744 8774
rect 11900 8634 11928 8978
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11900 8498 11928 8570
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11900 8090 11928 8434
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11610 7848 11666 7857
rect 11610 7783 11666 7792
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 11992 3505 12020 12294
rect 12268 9722 12296 15846
rect 12360 15706 12388 16458
rect 12452 15978 12480 16526
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 16114 13216 16390
rect 13740 16250 13768 16662
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14002 16552 14058 16561
rect 14002 16487 14058 16496
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12452 15586 12480 15914
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12452 15558 12572 15586
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12348 15156 12400 15162
rect 12452 15144 12480 15438
rect 12400 15116 12480 15144
rect 12348 15098 12400 15104
rect 12452 12986 12480 15116
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12544 12850 12572 15558
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12544 12442 12572 12786
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10538 12480 10950
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 12452 10062 12480 10474
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 11978 3496 12034 3505
rect 11978 3431 12034 3440
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 12084 1601 12112 9658
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12176 8974 12204 9590
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12452 9382 12480 9415
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8634 12204 8910
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12176 8362 12204 8570
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12636 2553 12664 15846
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 12806 15464 12862 15473
rect 12806 15399 12808 15408
rect 12860 15399 12862 15408
rect 13176 15428 13228 15434
rect 12808 15370 12860 15376
rect 13176 15370 13228 15376
rect 13188 14890 13216 15370
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 13082 14784 13138 14793
rect 12912 14657 12940 14758
rect 13082 14719 13138 14728
rect 12898 14648 12954 14657
rect 12898 14583 12954 14592
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12728 12238 12756 13942
rect 13096 12850 13124 14719
rect 13188 14278 13216 14826
rect 13372 14822 13400 15574
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 13394 13216 14214
rect 13372 13938 13400 14758
rect 13648 13954 13676 16050
rect 14016 15881 14044 16487
rect 14200 15881 14228 16594
rect 14660 16289 14688 16594
rect 14740 16448 14792 16454
rect 14738 16416 14740 16425
rect 15384 16448 15436 16454
rect 14792 16416 14794 16425
rect 15382 16416 15384 16425
rect 15436 16416 15438 16425
rect 14738 16351 14794 16360
rect 14956 16348 15252 16368
rect 15382 16351 15438 16360
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14646 16280 14702 16289
rect 14956 16272 15252 16292
rect 14646 16215 14702 16224
rect 14922 16144 14978 16153
rect 14922 16079 14978 16088
rect 14936 16046 14964 16079
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14660 15910 14688 15982
rect 14648 15904 14700 15910
rect 14002 15872 14058 15881
rect 14002 15807 14058 15816
rect 14186 15872 14242 15881
rect 14648 15846 14700 15852
rect 14186 15807 14242 15816
rect 14200 15706 14228 15807
rect 14936 15706 14964 15982
rect 15290 15736 15346 15745
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14924 15700 14976 15706
rect 15580 15706 15608 22374
rect 15856 22012 15884 22510
rect 15936 22500 15988 22506
rect 15936 22442 15988 22448
rect 15764 21984 15884 22012
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15672 17513 15700 17682
rect 15658 17504 15714 17513
rect 15658 17439 15714 17448
rect 15672 17338 15700 17439
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15290 15671 15346 15680
rect 15568 15700 15620 15706
rect 14924 15642 14976 15648
rect 15304 15570 15332 15671
rect 15568 15642 15620 15648
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15198 15056 15254 15065
rect 15198 14991 15254 15000
rect 15382 15056 15438 15065
rect 15382 14991 15438 15000
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13648 13926 13860 13954
rect 13452 13864 13504 13870
rect 13648 13841 13676 13926
rect 13452 13806 13504 13812
rect 13634 13832 13690 13841
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12889 13400 13126
rect 13358 12880 13414 12889
rect 13084 12844 13136 12850
rect 13358 12815 13414 12824
rect 13084 12786 13136 12792
rect 13096 12442 13124 12786
rect 13464 12442 13492 13806
rect 13634 13767 13690 13776
rect 13832 13530 13860 13926
rect 13924 13870 13952 14894
rect 14004 14884 14056 14890
rect 14004 14826 14056 14832
rect 14016 14618 14044 14826
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14016 14362 14044 14554
rect 15212 14550 15240 14991
rect 15292 14816 15344 14822
rect 15290 14784 15292 14793
rect 15344 14784 15346 14793
rect 15290 14719 15346 14728
rect 15396 14618 15424 14991
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 14016 14334 14136 14362
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13832 12782 13860 13466
rect 14016 12986 14044 14214
rect 14108 14074 14136 14334
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 15488 13954 15516 14758
rect 15658 14648 15714 14657
rect 15658 14583 15660 14592
rect 15712 14583 15714 14592
rect 15660 14554 15712 14560
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 14074 15608 14282
rect 15672 14074 15700 14554
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 14646 13832 14702 13841
rect 14646 13767 14648 13776
rect 14700 13767 14702 13776
rect 14648 13738 14700 13744
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14660 12850 14688 13738
rect 15028 13530 15056 13942
rect 15488 13926 15608 13954
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15580 13326 15608 13926
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12728 11898 12756 12174
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 13096 11558 13124 12242
rect 13464 11778 13492 12378
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11801 13676 12038
rect 13372 11750 13492 11778
rect 13634 11792 13690 11801
rect 13372 11694 13400 11750
rect 13634 11727 13690 11736
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9586 13032 9862
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9178 12940 9318
rect 13004 9178 13032 9522
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 13004 8430 13032 9114
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13004 8090 13032 8366
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13096 2961 13124 11494
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13268 11280 13320 11286
rect 13372 11257 13400 11290
rect 13268 11222 13320 11228
rect 13358 11248 13414 11257
rect 13280 10266 13308 11222
rect 13358 11183 13414 11192
rect 13556 11082 13584 11562
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13450 10432 13506 10441
rect 13450 10367 13506 10376
rect 13464 10266 13492 10367
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13740 9994 13768 11086
rect 13832 10282 13860 12174
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10810 13952 11086
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13832 10266 13952 10282
rect 13820 10260 13952 10266
rect 13872 10254 13952 10260
rect 13820 10202 13872 10208
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13832 9466 13860 10066
rect 13924 9722 13952 10254
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13740 9438 13860 9466
rect 14108 9450 14136 9998
rect 14096 9444 14148 9450
rect 13740 9382 13768 9438
rect 14096 9386 14148 9392
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13464 7449 13492 9318
rect 14108 9178 14136 9386
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14108 8634 14136 9114
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13450 7440 13506 7449
rect 13450 7375 13506 7384
rect 14384 6905 14412 12650
rect 15580 12646 15608 13262
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 14660 11558 14688 12174
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11218 14688 11494
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 15304 11150 15332 12174
rect 15488 12102 15516 12242
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15292 11144 15344 11150
rect 15488 11121 15516 12038
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15292 11086 15344 11092
rect 15474 11112 15530 11121
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10742 15332 11086
rect 15474 11047 15530 11056
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15304 10062 15332 10678
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 9998
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15580 7993 15608 11494
rect 15764 10810 15792 21984
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 17785 15884 19110
rect 15842 17776 15898 17785
rect 15842 17711 15898 17720
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 17134 15884 17614
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15856 16794 15884 17070
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15856 16250 15884 16730
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15948 12986 15976 22442
rect 16224 20913 16252 27520
rect 16776 24154 16804 27520
rect 17420 24585 17448 27520
rect 17406 24576 17462 24585
rect 17406 24511 17462 24520
rect 17314 24440 17370 24449
rect 17314 24375 17316 24384
rect 17368 24375 17370 24384
rect 17316 24346 17368 24352
rect 17316 24268 17368 24274
rect 17316 24210 17368 24216
rect 16500 24126 16804 24154
rect 16394 23896 16450 23905
rect 16394 23831 16396 23840
rect 16448 23831 16450 23840
rect 16396 23802 16448 23808
rect 16302 23624 16358 23633
rect 16302 23559 16358 23568
rect 16316 22778 16344 23559
rect 16500 23322 16528 24126
rect 17328 23526 17356 24210
rect 17972 23905 18000 27520
rect 17958 23896 18014 23905
rect 17958 23831 18014 23840
rect 18420 23656 18472 23662
rect 18418 23624 18420 23633
rect 18472 23624 18474 23633
rect 18418 23559 18474 23568
rect 16948 23520 17000 23526
rect 16762 23488 16818 23497
rect 16948 23462 17000 23468
rect 17316 23520 17368 23526
rect 18524 23497 18552 27520
rect 19076 24449 19104 27520
rect 19628 25922 19656 27520
rect 19444 25894 19656 25922
rect 19062 24440 19118 24449
rect 19062 24375 19118 24384
rect 18602 23896 18658 23905
rect 18602 23831 18604 23840
rect 18656 23831 18658 23840
rect 18604 23802 18656 23808
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19248 23588 19300 23594
rect 19248 23530 19300 23536
rect 17316 23462 17368 23468
rect 18510 23488 18566 23497
rect 16762 23423 16818 23432
rect 16776 23322 16804 23423
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16592 22778 16620 23122
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16210 20904 16266 20913
rect 16210 20839 16266 20848
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16316 18193 16344 18702
rect 16302 18184 16358 18193
rect 16302 18119 16358 18128
rect 16486 18184 16542 18193
rect 16486 18119 16542 18128
rect 16500 18086 16528 18119
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16212 16992 16264 16998
rect 16580 16992 16632 16998
rect 16212 16934 16264 16940
rect 16578 16960 16580 16969
rect 16632 16960 16634 16969
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16132 15706 16160 16594
rect 16224 16590 16252 16934
rect 16578 16895 16634 16904
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16224 15910 16252 16526
rect 16776 16504 16804 22714
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16684 16476 16804 16504
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16224 15502 16252 15846
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 14822 16252 15438
rect 16394 14920 16450 14929
rect 16394 14855 16450 14864
rect 16408 14822 16436 14855
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 16316 13938 16344 14486
rect 16500 14074 16528 14758
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15948 12238 15976 12582
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15856 10810 15884 11154
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10470 15700 10542
rect 15660 10464 15712 10470
rect 15658 10432 15660 10441
rect 15712 10432 15714 10441
rect 15658 10367 15714 10376
rect 15764 10198 15792 10610
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15764 9926 15792 10134
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15764 9382 15792 9862
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 9178 15792 9318
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15566 7984 15622 7993
rect 15566 7919 15622 7928
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14370 6896 14426 6905
rect 14370 6831 14426 6840
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 13910 4040 13966 4049
rect 13910 3975 13966 3984
rect 13082 2952 13138 2961
rect 13082 2887 13138 2896
rect 12622 2544 12678 2553
rect 12622 2479 12678 2488
rect 12070 1592 12126 1601
rect 12070 1527 12126 1536
rect 9954 1320 10010 1329
rect 9954 1255 10010 1264
rect 13924 480 13952 3975
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 16132 1737 16160 13670
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16224 12714 16252 13330
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16224 11354 16252 12650
rect 16316 11762 16344 13874
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16394 12472 16450 12481
rect 16394 12407 16396 12416
rect 16448 12407 16450 12416
rect 16396 12378 16448 12384
rect 16500 11898 16528 12582
rect 16684 12374 16712 16476
rect 16868 15910 16896 16662
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15706 16896 15846
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16868 15026 16896 15642
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16776 14618 16804 14826
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16868 14482 16896 14962
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16684 11898 16712 12174
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16592 11506 16620 11562
rect 16408 11478 16620 11506
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16408 9110 16436 11478
rect 16960 10810 16988 23462
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 17052 17882 17080 18022
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17236 17338 17264 17546
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 13530 17080 13874
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 12481 17080 12786
rect 17038 12472 17094 12481
rect 17038 12407 17094 12416
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17144 11762 17172 12310
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17144 11558 17172 11698
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11014 17172 11494
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16762 10704 16818 10713
rect 16762 10639 16818 10648
rect 16776 10606 16804 10639
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16500 10418 16528 10474
rect 16500 10390 16620 10418
rect 16592 9586 16620 10390
rect 17144 10266 17172 10950
rect 17328 10266 17356 23462
rect 18510 23423 18566 23432
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 17880 22506 17908 23122
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 18892 22438 18920 23122
rect 19260 23050 19288 23530
rect 19352 23322 19380 23598
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 17866 17912 17922 17921
rect 17866 17847 17922 17856
rect 17880 17746 17908 17847
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 17338 17908 17682
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 18050 17504 18106 17513
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17972 16833 18000 17478
rect 18050 17439 18106 17448
rect 18064 17202 18092 17439
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17958 16824 18014 16833
rect 17958 16759 18014 16768
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 16153 18092 16390
rect 18050 16144 18106 16153
rect 18050 16079 18106 16088
rect 18052 16040 18104 16046
rect 18050 16008 18052 16017
rect 18104 16008 18106 16017
rect 18050 15943 18106 15952
rect 18236 15904 18288 15910
rect 18234 15872 18236 15881
rect 18288 15872 18290 15881
rect 18234 15807 18290 15816
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17420 15162 17448 15506
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17420 14074 17448 15098
rect 18892 15065 18920 22374
rect 19444 19378 19472 25894
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19154 16688 19210 16697
rect 19154 16623 19156 16632
rect 19208 16623 19210 16632
rect 19156 16594 19208 16600
rect 19062 16416 19118 16425
rect 19062 16351 19118 16360
rect 19076 16046 19104 16351
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19260 15609 19288 15846
rect 19246 15600 19302 15609
rect 19246 15535 19302 15544
rect 18878 15056 18934 15065
rect 18878 14991 18934 15000
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17972 12646 18000 13262
rect 18050 12880 18106 12889
rect 18050 12815 18106 12824
rect 17960 12640 18012 12646
rect 17880 12588 17960 12594
rect 17880 12582 18012 12588
rect 17880 12566 18000 12582
rect 17880 11898 17908 12566
rect 17958 12472 18014 12481
rect 17958 12407 18014 12416
rect 17972 12170 18000 12407
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 18064 11898 18092 12815
rect 18156 12782 18184 13330
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18156 12481 18184 12718
rect 18142 12472 18198 12481
rect 18142 12407 18198 12416
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 18510 11792 18566 11801
rect 18510 11727 18566 11736
rect 18604 11756 18656 11762
rect 18524 11694 18552 11727
rect 18604 11698 18656 11704
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18616 11286 18644 11698
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17788 10470 17816 11154
rect 19352 10826 19380 17206
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19444 16561 19472 16730
rect 19892 16584 19944 16590
rect 19430 16552 19486 16561
rect 19892 16526 19944 16532
rect 19430 16487 19486 16496
rect 19904 16250 19932 16526
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19430 15464 19486 15473
rect 19430 15399 19486 15408
rect 19444 14958 19472 15399
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19430 13832 19486 13841
rect 19430 13767 19486 13776
rect 19444 13530 19472 13767
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 19314
rect 20272 17270 20300 27520
rect 20824 23905 20852 27520
rect 20810 23896 20866 23905
rect 21376 23866 21404 27520
rect 21822 24440 21878 24449
rect 21822 24375 21824 24384
rect 21876 24375 21878 24384
rect 21824 24346 21876 24352
rect 21928 24290 21956 27520
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21836 24262 21956 24290
rect 20810 23831 20866 23840
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20732 22438 20760 23122
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 19378 20760 22374
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 20626 16280 20682 16289
rect 20626 16215 20628 16224
rect 20680 16215 20682 16224
rect 20628 16186 20680 16192
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20456 15162 20484 15982
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20824 12782 20852 13330
rect 20812 12776 20864 12782
rect 20810 12744 20812 12753
rect 20864 12744 20866 12753
rect 20810 12679 20866 12688
rect 20916 12209 20944 19314
rect 21192 13530 21220 23598
rect 21560 23526 21588 24210
rect 21836 23798 21864 24262
rect 21914 23896 21970 23905
rect 21914 23831 21916 23840
rect 21968 23831 21970 23840
rect 21916 23802 21968 23808
rect 21824 23792 21876 23798
rect 21824 23734 21876 23740
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21560 23322 21588 23462
rect 22374 23352 22430 23361
rect 21548 23316 21600 23322
rect 22374 23287 22376 23296
rect 21548 23258 21600 23264
rect 22428 23287 22430 23296
rect 22376 23258 22428 23264
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22204 22438 22232 23122
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22112 16289 22140 16594
rect 22098 16280 22154 16289
rect 22098 16215 22154 16224
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 22204 13002 22232 22374
rect 22480 16658 22508 27520
rect 22926 24576 22982 24585
rect 22926 24511 22982 24520
rect 22940 24410 22968 24511
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 22744 24268 22796 24274
rect 22744 24210 22796 24216
rect 22756 23526 22784 24210
rect 23124 23905 23152 27520
rect 23676 24449 23704 27520
rect 23662 24440 23718 24449
rect 23662 24375 23718 24384
rect 24030 24440 24086 24449
rect 24030 24375 24032 24384
rect 24084 24375 24086 24384
rect 24032 24346 24084 24352
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23110 23896 23166 23905
rect 23110 23831 23166 23840
rect 23860 23662 23888 24210
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22020 12986 22232 13002
rect 22008 12980 22232 12986
rect 22060 12974 22232 12980
rect 22008 12922 22060 12928
rect 22282 12880 22338 12889
rect 22282 12815 22338 12824
rect 22296 12782 22324 12815
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 21100 12345 21128 12718
rect 22756 12442 22784 23462
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23308 22438 23336 23122
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23308 14929 23336 22374
rect 23294 14920 23350 14929
rect 23294 14855 23350 14864
rect 23492 13002 23520 23598
rect 23860 23322 23888 23598
rect 24228 23361 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24780 24585 24808 27520
rect 24766 24576 24822 24585
rect 24766 24511 24822 24520
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24950 23896 25006 23905
rect 24950 23831 24952 23840
rect 25004 23831 25006 23840
rect 24952 23802 25004 23808
rect 25332 23798 25360 27520
rect 25976 24449 26004 27520
rect 25962 24440 26018 24449
rect 25962 24375 26018 24384
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 24768 23656 24820 23662
rect 24768 23598 24820 23604
rect 24214 23352 24270 23361
rect 23848 23316 23900 23322
rect 24214 23287 24270 23296
rect 23848 23258 23900 23264
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24780 18426 24808 23598
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 23664 18216 23716 18222
rect 26528 18193 26556 27520
rect 27080 23905 27108 27520
rect 27632 24721 27660 27520
rect 27618 24712 27674 24721
rect 27618 24647 27674 24656
rect 27066 23896 27122 23905
rect 27066 23831 27122 23840
rect 23664 18158 23716 18164
rect 26514 18184 26570 18193
rect 23676 17649 23704 18158
rect 26514 18119 26570 18128
rect 23662 17640 23718 17649
rect 23662 17575 23718 17584
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 23400 12986 23520 13002
rect 23388 12980 23520 12986
rect 23440 12974 23520 12980
rect 23388 12922 23440 12928
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 21086 12336 21142 12345
rect 21086 12271 21142 12280
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 20902 12200 20958 12209
rect 20902 12135 20958 12144
rect 21744 11558 21772 12242
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 21744 11257 21772 11494
rect 21730 11248 21786 11257
rect 21730 11183 21786 11192
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19260 10810 19380 10826
rect 19248 10804 19380 10810
rect 19300 10798 19380 10804
rect 19248 10746 19300 10752
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16578 9344 16634 9353
rect 16578 9279 16634 9288
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16592 9042 16620 9279
rect 17788 9178 17816 10406
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18156 10033 18184 10066
rect 18142 10024 18198 10033
rect 18142 9959 18198 9968
rect 18156 9654 18184 9959
rect 18248 9722 18276 10542
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 9512 18104 9518
rect 18050 9480 18052 9489
rect 18104 9480 18106 9489
rect 18050 9415 18106 9424
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 8634 16620 8978
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 23202 3496 23258 3505
rect 23202 3431 23258 3440
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 16118 1728 16174 1737
rect 16118 1663 16174 1672
rect 23216 480 23244 3431
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 3054 368 3110 377
rect 3054 303 3110 312
rect 4618 0 4674 480
rect 13910 0 13966 480
rect 23202 0 23258 480
<< via2 >>
rect 2778 27648 2834 27704
rect 202 14864 258 14920
rect 1490 23568 1546 23624
rect 1582 23160 1638 23216
rect 1582 22480 1638 22536
rect 1582 21392 1638 21448
rect 1582 19624 1638 19680
rect 1490 17856 1546 17912
rect 1674 17448 1730 17504
rect 2042 24656 2098 24712
rect 2318 24828 2320 24848
rect 2320 24828 2372 24848
rect 2372 24828 2374 24848
rect 2318 24792 2374 24828
rect 1766 16496 1822 16552
rect 1674 15852 1676 15872
rect 1676 15852 1728 15872
rect 1728 15852 1730 15872
rect 1674 15816 1730 15852
rect 1674 14592 1730 14648
rect 2870 26560 2926 26616
rect 3054 25356 3110 25392
rect 3054 25336 3056 25356
rect 3056 25336 3108 25356
rect 3108 25336 3110 25356
rect 2778 21936 2834 21992
rect 2686 20868 2742 20904
rect 2686 20848 2688 20868
rect 2688 20848 2740 20868
rect 2740 20848 2742 20868
rect 2042 16088 2098 16144
rect 2134 15972 2190 16008
rect 2134 15952 2136 15972
rect 2136 15952 2188 15972
rect 2188 15952 2190 15972
rect 1858 15272 1914 15328
rect 1398 13640 1454 13696
rect 1398 9288 1454 9344
rect 1582 12280 1638 12336
rect 1858 13504 1914 13560
rect 1766 10648 1822 10704
rect 1858 10512 1914 10568
rect 2226 11192 2282 11248
rect 2502 19080 2558 19136
rect 2410 14456 2466 14512
rect 2410 10260 2466 10296
rect 2410 10240 2412 10260
rect 2412 10240 2464 10260
rect 2464 10240 2466 10260
rect 2410 9968 2466 10024
rect 2686 19080 2742 19136
rect 3238 23704 3294 23760
rect 3330 23296 3386 23352
rect 2870 18264 2926 18320
rect 3146 21120 3202 21176
rect 3882 27104 3938 27160
rect 3514 24248 3570 24304
rect 3330 20304 3386 20360
rect 3514 17584 3570 17640
rect 2686 16904 2742 16960
rect 2686 16496 2742 16552
rect 2962 16496 3018 16552
rect 2594 13232 2650 13288
rect 2686 12416 2742 12472
rect 2870 11056 2926 11112
rect 2870 10004 2872 10024
rect 2872 10004 2924 10024
rect 2924 10004 2926 10024
rect 2870 9968 2926 10004
rect 2962 9560 3018 9616
rect 2686 8900 2742 8936
rect 2686 8880 2688 8900
rect 2688 8880 2740 8900
rect 2740 8880 2742 8900
rect 2594 8372 2596 8392
rect 2596 8372 2648 8392
rect 2648 8372 2650 8392
rect 2594 8336 2650 8372
rect 570 4256 626 4312
rect 2686 3168 2742 3224
rect 2778 2896 2834 2952
rect 938 2488 994 2544
rect 938 1672 994 1728
rect 3698 24384 3754 24440
rect 4066 26016 4122 26072
rect 4066 24520 4122 24576
rect 3790 23432 3846 23488
rect 4434 24248 4490 24304
rect 4250 21936 4306 21992
rect 4066 19216 4122 19272
rect 4158 19080 4214 19136
rect 3882 17876 3938 17912
rect 3882 17856 3884 17876
rect 3884 17856 3936 17876
rect 3936 17856 3938 17876
rect 4250 18572 4252 18592
rect 4252 18572 4304 18592
rect 4304 18572 4306 18592
rect 4250 18536 4306 18572
rect 3790 16088 3846 16144
rect 4342 16088 4398 16144
rect 3606 14592 3662 14648
rect 3698 14320 3754 14376
rect 3606 12688 3662 12744
rect 3422 11600 3478 11656
rect 3514 11348 3570 11384
rect 3514 11328 3516 11348
rect 3516 11328 3568 11348
rect 3568 11328 3570 11348
rect 3606 6024 3662 6080
rect 4250 15544 4306 15600
rect 4250 15272 4306 15328
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4802 24384 4858 24440
rect 4986 24384 5042 24440
rect 4986 24112 5042 24168
rect 5446 24112 5502 24168
rect 5354 23724 5410 23760
rect 5354 23704 5356 23724
rect 5356 23704 5408 23724
rect 5408 23704 5410 23724
rect 4802 21936 4858 21992
rect 5998 24520 6054 24576
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5538 23296 5594 23352
rect 5998 23024 6054 23080
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5354 22480 5410 22536
rect 5998 21800 6054 21856
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 4986 20848 5042 20904
rect 5538 20984 5594 21040
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 6182 24812 6238 24848
rect 6182 24792 6184 24812
rect 6184 24792 6236 24812
rect 6236 24792 6238 24812
rect 6550 24656 6606 24712
rect 6550 23468 6552 23488
rect 6552 23468 6604 23488
rect 6604 23468 6606 23488
rect 6550 23432 6606 23468
rect 5446 20324 5502 20360
rect 5446 20304 5448 20324
rect 5448 20304 5500 20324
rect 5500 20304 5502 20324
rect 4894 18264 4950 18320
rect 5078 18164 5080 18184
rect 5080 18164 5132 18184
rect 5132 18164 5134 18184
rect 5078 18128 5134 18164
rect 4526 14864 4582 14920
rect 6458 20712 6514 20768
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5078 16768 5134 16824
rect 6182 16904 6238 16960
rect 6458 16904 6514 16960
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5170 15852 5172 15872
rect 5172 15852 5224 15872
rect 5224 15852 5226 15872
rect 5170 15816 5226 15852
rect 4802 14456 4858 14512
rect 4250 12824 4306 12880
rect 4066 12552 4122 12608
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4802 13812 4804 13832
rect 4804 13812 4856 13832
rect 4856 13812 4858 13832
rect 4802 13776 4858 13812
rect 4710 13676 4712 13696
rect 4712 13676 4764 13696
rect 4764 13676 4766 13696
rect 4710 13640 4766 13676
rect 6274 16496 6330 16552
rect 5998 14456 6054 14512
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5538 13912 5594 13968
rect 5446 13504 5502 13560
rect 6274 13640 6330 13696
rect 5998 13232 6054 13288
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5814 12844 5870 12880
rect 5814 12824 5816 12844
rect 5816 12824 5868 12844
rect 5868 12824 5870 12844
rect 3974 11736 4030 11792
rect 4526 11212 4582 11248
rect 4526 11192 4528 11212
rect 4528 11192 4580 11212
rect 4580 11192 4582 11212
rect 4066 11076 4122 11112
rect 4066 11056 4068 11076
rect 4068 11056 4120 11076
rect 4120 11056 4122 11076
rect 4158 10240 4214 10296
rect 5262 12300 5318 12336
rect 5262 12280 5264 12300
rect 5264 12280 5316 12300
rect 5316 12280 5318 12300
rect 5170 12144 5226 12200
rect 5722 12280 5778 12336
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6182 12588 6184 12608
rect 6184 12588 6236 12608
rect 6236 12588 6238 12608
rect 6182 12552 6238 12588
rect 6366 12280 6422 12336
rect 6550 12960 6606 13016
rect 6550 12688 6606 12744
rect 6550 11620 6606 11656
rect 6550 11600 6552 11620
rect 6552 11600 6604 11620
rect 6604 11600 6606 11620
rect 7102 23568 7158 23624
rect 7562 22072 7618 22128
rect 8206 24792 8262 24848
rect 8206 24676 8262 24712
rect 8206 24656 8208 24676
rect 8208 24656 8260 24676
rect 8260 24656 8262 24676
rect 7930 24384 7986 24440
rect 8114 23976 8170 24032
rect 7930 23296 7986 23352
rect 8850 23296 8906 23352
rect 7838 22072 7894 22128
rect 7654 21120 7710 21176
rect 8114 20576 8170 20632
rect 8114 18828 8170 18864
rect 8114 18808 8116 18828
rect 8116 18808 8168 18828
rect 8168 18808 8170 18828
rect 7562 18708 7564 18728
rect 7564 18708 7616 18728
rect 7616 18708 7618 18728
rect 7562 18672 7618 18708
rect 7562 18536 7618 18592
rect 8022 17740 8078 17776
rect 8022 17720 8024 17740
rect 8024 17720 8076 17740
rect 8076 17720 8078 17740
rect 7930 17176 7986 17232
rect 7378 16768 7434 16824
rect 7010 16360 7066 16416
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9402 21392 9458 21448
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9862 23024 9918 23080
rect 10966 24792 11022 24848
rect 10690 23704 10746 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 8574 20576 8630 20632
rect 8390 17584 8446 17640
rect 9678 19352 9734 19408
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10690 20984 10746 21040
rect 10782 20460 10838 20496
rect 10782 20440 10784 20460
rect 10784 20440 10836 20460
rect 10836 20440 10838 20460
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9770 18944 9826 19000
rect 9954 18572 9956 18592
rect 9956 18572 10008 18592
rect 10008 18572 10010 18592
rect 9954 18536 10010 18572
rect 9862 17856 9918 17912
rect 9678 17176 9734 17232
rect 7562 16224 7618 16280
rect 7562 15680 7618 15736
rect 7562 15564 7618 15600
rect 7562 15544 7564 15564
rect 7564 15544 7616 15564
rect 7616 15544 7618 15564
rect 9494 15952 9550 16008
rect 7378 15272 7434 15328
rect 7838 15136 7894 15192
rect 8390 14476 8446 14512
rect 8390 14456 8392 14476
rect 8392 14456 8444 14476
rect 8444 14456 8446 14476
rect 6826 12688 6882 12744
rect 6734 11500 6736 11520
rect 6736 11500 6788 11520
rect 6788 11500 6790 11520
rect 6734 11464 6790 11500
rect 6642 11328 6698 11384
rect 7194 12144 7250 12200
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 7562 13504 7618 13560
rect 8298 13812 8300 13832
rect 8300 13812 8352 13832
rect 8352 13812 8354 13832
rect 8298 13776 8354 13812
rect 8574 13640 8630 13696
rect 7654 13368 7710 13424
rect 7838 12416 7894 12472
rect 7746 12164 7802 12200
rect 7746 12144 7748 12164
rect 7748 12144 7800 12164
rect 7800 12144 7802 12164
rect 7930 11736 7986 11792
rect 8390 11464 8446 11520
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5354 9424 5410 9480
rect 4894 9152 4950 9208
rect 4894 8880 4950 8936
rect 5078 8900 5134 8936
rect 5078 8880 5080 8900
rect 5080 8880 5132 8900
rect 5132 8880 5134 8900
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 7654 9988 7710 10024
rect 7654 9968 7656 9988
rect 7656 9968 7708 9988
rect 7708 9968 7710 9988
rect 7838 9016 7894 9072
rect 10046 16496 10102 16552
rect 9770 15816 9826 15872
rect 9678 15000 9734 15056
rect 9770 14456 9826 14512
rect 9034 9696 9090 9752
rect 9586 9424 9642 9480
rect 10046 14612 10102 14648
rect 10046 14592 10048 14612
rect 10048 14592 10100 14612
rect 10100 14592 10102 14612
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 11702 24792 11758 24848
rect 11150 24112 11206 24168
rect 12162 24112 12218 24168
rect 11794 23976 11850 24032
rect 12070 23432 12126 23488
rect 11058 21936 11114 21992
rect 11058 17040 11114 17096
rect 10966 16088 11022 16144
rect 10966 15852 10968 15872
rect 10968 15852 11020 15872
rect 11020 15852 11022 15872
rect 10966 15816 11022 15852
rect 10690 15544 10746 15600
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10322 14320 10378 14376
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10138 13524 10194 13560
rect 10138 13504 10140 13524
rect 10140 13504 10192 13524
rect 10192 13504 10194 13524
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10138 12316 10140 12336
rect 10140 12316 10192 12336
rect 10192 12316 10194 12336
rect 10138 12280 10194 12316
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10046 10376 10102 10432
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9862 10104 9918 10160
rect 10322 10104 10378 10160
rect 9862 9832 9918 9888
rect 9770 9560 9826 9616
rect 8114 8880 8170 8936
rect 8942 8916 8944 8936
rect 8944 8916 8996 8936
rect 8996 8916 8998 8936
rect 8942 8880 8998 8916
rect 4066 7928 4122 7984
rect 3974 7792 4030 7848
rect 3698 5344 3754 5400
rect 3422 4800 3478 4856
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 4066 7112 4122 7168
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 9862 9152 9918 9208
rect 9770 8336 9826 8392
rect 3974 3712 4030 3768
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 9494 3984 9550 4040
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10230 9696 10286 9752
rect 10138 9288 10194 9344
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10598 8492 10654 8528
rect 10598 8472 10600 8492
rect 10600 8472 10652 8492
rect 10652 8472 10654 8492
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11426 16788 11482 16824
rect 11426 16768 11428 16788
rect 11428 16768 11480 16788
rect 11480 16768 11482 16788
rect 12438 22500 12494 22536
rect 12438 22480 12440 22500
rect 12440 22480 12492 22500
rect 12492 22480 12494 22500
rect 12162 20712 12218 20768
rect 12530 20340 12532 20360
rect 12532 20340 12584 20360
rect 12584 20340 12586 20360
rect 12530 20304 12586 20340
rect 11702 16632 11758 16688
rect 11610 16360 11666 16416
rect 11242 15408 11298 15464
rect 11702 15136 11758 15192
rect 11426 13776 11482 13832
rect 11242 12280 11298 12336
rect 13818 21392 13874 21448
rect 14554 24792 14610 24848
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15658 24520 15714 24576
rect 15382 24248 15438 24304
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15106 23468 15108 23488
rect 15108 23468 15160 23488
rect 15160 23468 15162 23488
rect 15106 23432 15162 23468
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14738 21800 14794 21856
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14094 20848 14150 20904
rect 14278 20848 14334 20904
rect 13910 20440 13966 20496
rect 14002 18808 14058 18864
rect 13358 18672 13414 18728
rect 13450 17992 13506 18048
rect 13174 17856 13230 17912
rect 13082 17604 13138 17640
rect 13082 17584 13084 17604
rect 13084 17584 13136 17604
rect 13136 17584 13138 17604
rect 13082 16904 13138 16960
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14554 20576 14610 20632
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15290 19352 15346 19408
rect 15106 19216 15162 19272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14922 18300 14924 18320
rect 14924 18300 14976 18320
rect 14976 18300 14978 18320
rect 14922 18264 14978 18300
rect 15290 17992 15346 18048
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 12070 14728 12126 14784
rect 12162 12980 12218 13016
rect 12162 12960 12164 12980
rect 12164 12960 12216 12980
rect 12216 12960 12218 12980
rect 11150 9832 11206 9888
rect 11242 9716 11298 9752
rect 11242 9696 11244 9716
rect 11244 9696 11296 9716
rect 11296 9696 11298 9716
rect 11610 7792 11666 7848
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 14002 16496 14058 16552
rect 11978 3440 12034 3496
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12438 9424 12494 9480
rect 12806 15428 12862 15464
rect 12806 15408 12808 15428
rect 12808 15408 12860 15428
rect 12860 15408 12862 15428
rect 13082 14728 13138 14784
rect 12898 14592 12954 14648
rect 14738 16396 14740 16416
rect 14740 16396 14792 16416
rect 14792 16396 14794 16416
rect 14738 16360 14794 16396
rect 15382 16396 15384 16416
rect 15384 16396 15436 16416
rect 15436 16396 15438 16416
rect 15382 16360 15438 16396
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14646 16224 14702 16280
rect 14922 16088 14978 16144
rect 14002 15816 14058 15872
rect 14186 15816 14242 15872
rect 15290 15680 15346 15736
rect 15658 17448 15714 17504
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15198 15000 15254 15056
rect 15382 15000 15438 15056
rect 13358 12824 13414 12880
rect 13634 13776 13690 13832
rect 15290 14764 15292 14784
rect 15292 14764 15344 14784
rect 15344 14764 15346 14784
rect 15290 14728 15346 14764
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15658 14612 15714 14648
rect 15658 14592 15660 14612
rect 15660 14592 15712 14612
rect 15712 14592 15714 14612
rect 14646 13796 14702 13832
rect 14646 13776 14648 13796
rect 14648 13776 14700 13796
rect 14700 13776 14702 13796
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 13634 11736 13690 11792
rect 13358 11192 13414 11248
rect 13450 10376 13506 10432
rect 13450 7384 13506 7440
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15474 11056 15530 11112
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15842 17720 15898 17776
rect 17406 24520 17462 24576
rect 17314 24404 17370 24440
rect 17314 24384 17316 24404
rect 17316 24384 17368 24404
rect 17368 24384 17370 24404
rect 16394 23860 16450 23896
rect 16394 23840 16396 23860
rect 16396 23840 16448 23860
rect 16448 23840 16450 23860
rect 16302 23568 16358 23624
rect 17958 23840 18014 23896
rect 18418 23604 18420 23624
rect 18420 23604 18472 23624
rect 18472 23604 18474 23624
rect 18418 23568 18474 23604
rect 16762 23432 16818 23488
rect 19062 24384 19118 24440
rect 18602 23860 18658 23896
rect 18602 23840 18604 23860
rect 18604 23840 18656 23860
rect 18656 23840 18658 23860
rect 16210 20848 16266 20904
rect 16302 18128 16358 18184
rect 16486 18128 16542 18184
rect 16578 16940 16580 16960
rect 16580 16940 16632 16960
rect 16632 16940 16634 16960
rect 16578 16904 16634 16940
rect 16394 14864 16450 14920
rect 15658 10412 15660 10432
rect 15660 10412 15712 10432
rect 15712 10412 15714 10432
rect 15658 10376 15714 10412
rect 15566 7928 15622 7984
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14370 6840 14426 6896
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 13910 3984 13966 4040
rect 13082 2896 13138 2952
rect 12622 2488 12678 2544
rect 12070 1536 12126 1592
rect 9954 1264 10010 1320
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16394 12436 16450 12472
rect 16394 12416 16396 12436
rect 16396 12416 16448 12436
rect 16448 12416 16450 12436
rect 17038 12416 17094 12472
rect 16762 10648 16818 10704
rect 18510 23432 18566 23488
rect 17866 17856 17922 17912
rect 18050 17448 18106 17504
rect 17958 16768 18014 16824
rect 18050 16088 18106 16144
rect 18050 15988 18052 16008
rect 18052 15988 18104 16008
rect 18104 15988 18106 16008
rect 18050 15952 18106 15988
rect 18234 15852 18236 15872
rect 18236 15852 18288 15872
rect 18288 15852 18290 15872
rect 18234 15816 18290 15852
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19154 16652 19210 16688
rect 19154 16632 19156 16652
rect 19156 16632 19208 16652
rect 19208 16632 19210 16652
rect 19062 16360 19118 16416
rect 19246 15544 19302 15600
rect 18878 15000 18934 15056
rect 18050 12824 18106 12880
rect 17958 12416 18014 12472
rect 18142 12416 18198 12472
rect 18510 11736 18566 11792
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19430 16496 19486 16552
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19430 15408 19486 15464
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19430 13776 19486 13832
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20810 23840 20866 23896
rect 21822 24404 21878 24440
rect 21822 24384 21824 24404
rect 21824 24384 21876 24404
rect 21876 24384 21878 24404
rect 20626 16244 20682 16280
rect 20626 16224 20628 16244
rect 20628 16224 20680 16244
rect 20680 16224 20682 16244
rect 20810 12724 20812 12744
rect 20812 12724 20864 12744
rect 20864 12724 20866 12744
rect 20810 12688 20866 12724
rect 21914 23860 21970 23896
rect 21914 23840 21916 23860
rect 21916 23840 21968 23860
rect 21968 23840 21970 23860
rect 22374 23316 22430 23352
rect 22374 23296 22376 23316
rect 22376 23296 22428 23316
rect 22428 23296 22430 23316
rect 22098 16224 22154 16280
rect 22926 24520 22982 24576
rect 23662 24384 23718 24440
rect 24030 24404 24086 24440
rect 24030 24384 24032 24404
rect 24032 24384 24084 24404
rect 24084 24384 24086 24404
rect 23110 23840 23166 23896
rect 22282 12824 22338 12880
rect 23294 14864 23350 14920
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24520 24822 24576
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24950 23860 25006 23896
rect 24950 23840 24952 23860
rect 24952 23840 25004 23860
rect 25004 23840 25006 23860
rect 25962 24384 26018 24440
rect 24214 23296 24270 23352
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 27618 24656 27674 24712
rect 27066 23840 27122 23896
rect 26514 18128 26570 18184
rect 23662 17584 23718 17640
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 21086 12280 21142 12336
rect 20902 12144 20958 12200
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 21730 11192 21786 11248
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 16578 9288 16634 9344
rect 18142 9968 18198 10024
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 18050 9460 18052 9480
rect 18052 9460 18104 9480
rect 18104 9460 18106 9480
rect 18050 9424 18106 9460
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 23202 3440 23258 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 16118 1672 16174 1728
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 3054 312 3110 368
<< metal3 >>
rect 0 27706 480 27736
rect 2773 27706 2839 27709
rect 0 27704 2839 27706
rect 0 27648 2778 27704
rect 2834 27648 2839 27704
rect 0 27646 2839 27648
rect 0 27616 480 27646
rect 2773 27643 2839 27646
rect 0 27162 480 27192
rect 3877 27162 3943 27165
rect 0 27160 3943 27162
rect 0 27104 3882 27160
rect 3938 27104 3943 27160
rect 0 27102 3943 27104
rect 0 27072 480 27102
rect 3877 27099 3943 27102
rect 0 26618 480 26648
rect 2865 26618 2931 26621
rect 0 26616 2931 26618
rect 0 26560 2870 26616
rect 2926 26560 2931 26616
rect 0 26558 2931 26560
rect 0 26528 480 26558
rect 2865 26555 2931 26558
rect 0 26074 480 26104
rect 4061 26074 4127 26077
rect 0 26072 4127 26074
rect 0 26016 4066 26072
rect 4122 26016 4127 26072
rect 0 26014 4127 26016
rect 0 25984 480 26014
rect 4061 26011 4127 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 3049 25394 3115 25397
rect 0 25392 3115 25394
rect 0 25336 3054 25392
rect 3110 25336 3115 25392
rect 0 25334 3115 25336
rect 0 25304 480 25334
rect 3049 25331 3115 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 2313 24850 2379 24853
rect 6177 24850 6243 24853
rect 8201 24850 8267 24853
rect 0 24790 1410 24850
rect 0 24760 480 24790
rect 1350 24578 1410 24790
rect 2313 24848 4722 24850
rect 2313 24792 2318 24848
rect 2374 24792 4722 24848
rect 2313 24790 4722 24792
rect 2313 24787 2379 24790
rect 2037 24714 2103 24717
rect 4662 24714 4722 24790
rect 6177 24848 8267 24850
rect 6177 24792 6182 24848
rect 6238 24792 8206 24848
rect 8262 24792 8267 24848
rect 6177 24790 8267 24792
rect 6177 24787 6243 24790
rect 8201 24787 8267 24790
rect 10961 24850 11027 24853
rect 11697 24850 11763 24853
rect 14549 24850 14615 24853
rect 10961 24848 11763 24850
rect 10961 24792 10966 24848
rect 11022 24792 11702 24848
rect 11758 24792 11763 24848
rect 10961 24790 11763 24792
rect 10961 24787 11027 24790
rect 11697 24787 11763 24790
rect 11838 24848 14615 24850
rect 11838 24792 14554 24848
rect 14610 24792 14615 24848
rect 11838 24790 14615 24792
rect 6545 24714 6611 24717
rect 2037 24712 4354 24714
rect 2037 24656 2042 24712
rect 2098 24656 4354 24712
rect 2037 24654 4354 24656
rect 4662 24712 6611 24714
rect 4662 24656 6550 24712
rect 6606 24656 6611 24712
rect 4662 24654 6611 24656
rect 2037 24651 2103 24654
rect 4061 24578 4127 24581
rect 1350 24576 4127 24578
rect 1350 24520 4066 24576
rect 4122 24520 4127 24576
rect 1350 24518 4127 24520
rect 4294 24578 4354 24654
rect 6545 24651 6611 24654
rect 8201 24714 8267 24717
rect 11838 24714 11898 24790
rect 14549 24787 14615 24790
rect 27613 24714 27679 24717
rect 8201 24712 11898 24714
rect 8201 24656 8206 24712
rect 8262 24656 11898 24712
rect 8201 24654 11898 24656
rect 15518 24712 27679 24714
rect 15518 24656 27618 24712
rect 27674 24656 27679 24712
rect 15518 24654 27679 24656
rect 8201 24651 8267 24654
rect 5993 24578 6059 24581
rect 4294 24576 6059 24578
rect 4294 24520 5998 24576
rect 6054 24520 6059 24576
rect 4294 24518 6059 24520
rect 4061 24515 4127 24518
rect 5993 24515 6059 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 3693 24442 3759 24445
rect 4797 24442 4863 24445
rect 3693 24440 4863 24442
rect 3693 24384 3698 24440
rect 3754 24384 4802 24440
rect 4858 24384 4863 24440
rect 3693 24382 4863 24384
rect 3693 24379 3759 24382
rect 4797 24379 4863 24382
rect 4981 24442 5047 24445
rect 7925 24442 7991 24445
rect 4981 24440 7991 24442
rect 4981 24384 4986 24440
rect 5042 24384 7930 24440
rect 7986 24384 7991 24440
rect 4981 24382 7991 24384
rect 4981 24379 5047 24382
rect 7925 24379 7991 24382
rect 0 24306 480 24336
rect 3509 24306 3575 24309
rect 0 24304 3575 24306
rect 0 24248 3514 24304
rect 3570 24248 3575 24304
rect 0 24246 3575 24248
rect 0 24216 480 24246
rect 3509 24243 3575 24246
rect 4429 24306 4495 24309
rect 15377 24306 15443 24309
rect 4429 24304 15443 24306
rect 4429 24248 4434 24304
rect 4490 24248 15382 24304
rect 15438 24248 15443 24304
rect 4429 24246 15443 24248
rect 4429 24243 4495 24246
rect 15377 24243 15443 24246
rect 4981 24170 5047 24173
rect 5441 24170 5507 24173
rect 11145 24170 11211 24173
rect 4981 24168 11211 24170
rect 4981 24112 4986 24168
rect 5042 24112 5446 24168
rect 5502 24112 11150 24168
rect 11206 24112 11211 24168
rect 4981 24110 11211 24112
rect 4981 24107 5047 24110
rect 5441 24107 5507 24110
rect 11145 24107 11211 24110
rect 12157 24170 12223 24173
rect 15518 24170 15578 24654
rect 27613 24651 27679 24654
rect 15653 24578 15719 24581
rect 17401 24578 17467 24581
rect 15653 24576 17467 24578
rect 15653 24520 15658 24576
rect 15714 24520 17406 24576
rect 17462 24520 17467 24576
rect 15653 24518 17467 24520
rect 15653 24515 15719 24518
rect 17401 24515 17467 24518
rect 22921 24578 22987 24581
rect 24761 24578 24827 24581
rect 22921 24576 24827 24578
rect 22921 24520 22926 24576
rect 22982 24520 24766 24576
rect 24822 24520 24827 24576
rect 22921 24518 24827 24520
rect 22921 24515 22987 24518
rect 24761 24515 24827 24518
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 17309 24442 17375 24445
rect 19057 24442 19123 24445
rect 17309 24440 19123 24442
rect 17309 24384 17314 24440
rect 17370 24384 19062 24440
rect 19118 24384 19123 24440
rect 17309 24382 19123 24384
rect 17309 24379 17375 24382
rect 19057 24379 19123 24382
rect 21817 24442 21883 24445
rect 23657 24442 23723 24445
rect 21817 24440 23723 24442
rect 21817 24384 21822 24440
rect 21878 24384 23662 24440
rect 23718 24384 23723 24440
rect 21817 24382 23723 24384
rect 21817 24379 21883 24382
rect 23657 24379 23723 24382
rect 24025 24442 24091 24445
rect 25957 24442 26023 24445
rect 24025 24440 26023 24442
rect 24025 24384 24030 24440
rect 24086 24384 25962 24440
rect 26018 24384 26023 24440
rect 24025 24382 26023 24384
rect 24025 24379 24091 24382
rect 25957 24379 26023 24382
rect 12157 24168 15578 24170
rect 12157 24112 12162 24168
rect 12218 24112 15578 24168
rect 12157 24110 15578 24112
rect 12157 24107 12223 24110
rect 8109 24034 8175 24037
rect 11789 24034 11855 24037
rect 8109 24032 11855 24034
rect 8109 23976 8114 24032
rect 8170 23976 11794 24032
rect 11850 23976 11855 24032
rect 8109 23974 11855 23976
rect 8109 23971 8175 23974
rect 11789 23971 11855 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 16389 23898 16455 23901
rect 17953 23898 18019 23901
rect 16389 23896 18019 23898
rect 16389 23840 16394 23896
rect 16450 23840 17958 23896
rect 18014 23840 18019 23896
rect 16389 23838 18019 23840
rect 16389 23835 16455 23838
rect 17953 23835 18019 23838
rect 18597 23898 18663 23901
rect 20805 23898 20871 23901
rect 18597 23896 20871 23898
rect 18597 23840 18602 23896
rect 18658 23840 20810 23896
rect 20866 23840 20871 23896
rect 18597 23838 20871 23840
rect 18597 23835 18663 23838
rect 20805 23835 20871 23838
rect 21909 23898 21975 23901
rect 23105 23898 23171 23901
rect 21909 23896 23171 23898
rect 21909 23840 21914 23896
rect 21970 23840 23110 23896
rect 23166 23840 23171 23896
rect 21909 23838 23171 23840
rect 21909 23835 21975 23838
rect 23105 23835 23171 23838
rect 24945 23898 25011 23901
rect 27061 23898 27127 23901
rect 24945 23896 27127 23898
rect 24945 23840 24950 23896
rect 25006 23840 27066 23896
rect 27122 23840 27127 23896
rect 24945 23838 27127 23840
rect 24945 23835 25011 23838
rect 27061 23835 27127 23838
rect 0 23762 480 23792
rect 3233 23762 3299 23765
rect 0 23760 3299 23762
rect 0 23704 3238 23760
rect 3294 23704 3299 23760
rect 0 23702 3299 23704
rect 0 23672 480 23702
rect 3233 23699 3299 23702
rect 5349 23762 5415 23765
rect 10685 23762 10751 23765
rect 5349 23760 10751 23762
rect 5349 23704 5354 23760
rect 5410 23704 10690 23760
rect 10746 23704 10751 23760
rect 5349 23702 10751 23704
rect 5349 23699 5415 23702
rect 10685 23699 10751 23702
rect 1485 23626 1551 23629
rect 7097 23626 7163 23629
rect 1485 23624 7163 23626
rect 1485 23568 1490 23624
rect 1546 23568 7102 23624
rect 7158 23568 7163 23624
rect 1485 23566 7163 23568
rect 1485 23563 1551 23566
rect 7097 23563 7163 23566
rect 16297 23626 16363 23629
rect 18413 23626 18479 23629
rect 16297 23624 18479 23626
rect 16297 23568 16302 23624
rect 16358 23568 18418 23624
rect 18474 23568 18479 23624
rect 16297 23566 18479 23568
rect 16297 23563 16363 23566
rect 18413 23563 18479 23566
rect 3785 23490 3851 23493
rect 6545 23490 6611 23493
rect 3785 23488 6611 23490
rect 3785 23432 3790 23488
rect 3846 23432 6550 23488
rect 6606 23432 6611 23488
rect 3785 23430 6611 23432
rect 3785 23427 3851 23430
rect 6545 23427 6611 23430
rect 12065 23490 12131 23493
rect 15101 23490 15167 23493
rect 12065 23488 15167 23490
rect 12065 23432 12070 23488
rect 12126 23432 15106 23488
rect 15162 23432 15167 23488
rect 12065 23430 15167 23432
rect 12065 23427 12131 23430
rect 15101 23427 15167 23430
rect 16757 23490 16823 23493
rect 18505 23490 18571 23493
rect 16757 23488 18571 23490
rect 16757 23432 16762 23488
rect 16818 23432 18510 23488
rect 18566 23432 18571 23488
rect 16757 23430 18571 23432
rect 16757 23427 16823 23430
rect 18505 23427 18571 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 3325 23354 3391 23357
rect 5533 23354 5599 23357
rect 3325 23352 5599 23354
rect 3325 23296 3330 23352
rect 3386 23296 5538 23352
rect 5594 23296 5599 23352
rect 3325 23294 5599 23296
rect 3325 23291 3391 23294
rect 5533 23291 5599 23294
rect 7925 23354 7991 23357
rect 8845 23354 8911 23357
rect 7925 23352 8911 23354
rect 7925 23296 7930 23352
rect 7986 23296 8850 23352
rect 8906 23296 8911 23352
rect 7925 23294 8911 23296
rect 7925 23291 7991 23294
rect 8845 23291 8911 23294
rect 22369 23354 22435 23357
rect 24209 23354 24275 23357
rect 22369 23352 24275 23354
rect 22369 23296 22374 23352
rect 22430 23296 24214 23352
rect 24270 23296 24275 23352
rect 22369 23294 24275 23296
rect 22369 23291 22435 23294
rect 24209 23291 24275 23294
rect 0 23218 480 23248
rect 1577 23218 1643 23221
rect 0 23216 1643 23218
rect 0 23160 1582 23216
rect 1638 23160 1643 23216
rect 0 23158 1643 23160
rect 0 23128 480 23158
rect 1577 23155 1643 23158
rect 5993 23082 6059 23085
rect 9857 23082 9923 23085
rect 5993 23080 9923 23082
rect 5993 23024 5998 23080
rect 6054 23024 9862 23080
rect 9918 23024 9923 23080
rect 5993 23022 9923 23024
rect 5993 23019 6059 23022
rect 9857 23019 9923 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22538 480 22568
rect 1577 22538 1643 22541
rect 0 22536 1643 22538
rect 0 22480 1582 22536
rect 1638 22480 1643 22536
rect 0 22478 1643 22480
rect 0 22448 480 22478
rect 1577 22475 1643 22478
rect 5349 22538 5415 22541
rect 12433 22538 12499 22541
rect 5349 22536 12499 22538
rect 5349 22480 5354 22536
rect 5410 22480 12438 22536
rect 12494 22480 12499 22536
rect 5349 22478 12499 22480
rect 5349 22475 5415 22478
rect 12433 22475 12499 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 7557 22130 7623 22133
rect 7833 22130 7899 22133
rect 7557 22128 7899 22130
rect 7557 22072 7562 22128
rect 7618 22072 7838 22128
rect 7894 22072 7899 22128
rect 7557 22070 7899 22072
rect 7557 22067 7623 22070
rect 7833 22067 7899 22070
rect 0 21994 480 22024
rect 2773 21994 2839 21997
rect 0 21992 2839 21994
rect 0 21936 2778 21992
rect 2834 21936 2839 21992
rect 0 21934 2839 21936
rect 0 21904 480 21934
rect 2773 21931 2839 21934
rect 4245 21994 4311 21997
rect 4797 21994 4863 21997
rect 11053 21994 11119 21997
rect 4245 21992 11119 21994
rect 4245 21936 4250 21992
rect 4306 21936 4802 21992
rect 4858 21936 11058 21992
rect 11114 21936 11119 21992
rect 4245 21934 11119 21936
rect 4245 21931 4311 21934
rect 4797 21931 4863 21934
rect 11053 21931 11119 21934
rect 5993 21858 6059 21861
rect 14733 21858 14799 21861
rect 5993 21856 14799 21858
rect 5993 21800 5998 21856
rect 6054 21800 14738 21856
rect 14794 21800 14799 21856
rect 5993 21798 14799 21800
rect 5993 21795 6059 21798
rect 14733 21795 14799 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21450 480 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 480 21390
rect 1577 21387 1643 21390
rect 9397 21450 9463 21453
rect 13813 21450 13879 21453
rect 9397 21448 13879 21450
rect 9397 21392 9402 21448
rect 9458 21392 13818 21448
rect 13874 21392 13879 21448
rect 9397 21390 13879 21392
rect 9397 21387 9463 21390
rect 13813 21387 13879 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 3141 21178 3207 21181
rect 7649 21178 7715 21181
rect 3141 21176 7715 21178
rect 3141 21120 3146 21176
rect 3202 21120 7654 21176
rect 7710 21120 7715 21176
rect 3141 21118 7715 21120
rect 3141 21115 3207 21118
rect 7649 21115 7715 21118
rect 5533 21042 5599 21045
rect 10685 21042 10751 21045
rect 5533 21040 10751 21042
rect 5533 20984 5538 21040
rect 5594 20984 10690 21040
rect 10746 20984 10751 21040
rect 5533 20982 10751 20984
rect 5533 20979 5599 20982
rect 10685 20979 10751 20982
rect 0 20906 480 20936
rect 2681 20906 2747 20909
rect 0 20904 2747 20906
rect 0 20848 2686 20904
rect 2742 20848 2747 20904
rect 0 20846 2747 20848
rect 0 20816 480 20846
rect 2681 20843 2747 20846
rect 4981 20906 5047 20909
rect 14089 20906 14155 20909
rect 4981 20904 14155 20906
rect 4981 20848 4986 20904
rect 5042 20848 14094 20904
rect 14150 20848 14155 20904
rect 4981 20846 14155 20848
rect 4981 20843 5047 20846
rect 14089 20843 14155 20846
rect 14273 20906 14339 20909
rect 16205 20906 16271 20909
rect 14273 20904 16271 20906
rect 14273 20848 14278 20904
rect 14334 20848 16210 20904
rect 16266 20848 16271 20904
rect 14273 20846 16271 20848
rect 14273 20843 14339 20846
rect 16205 20843 16271 20846
rect 6453 20770 6519 20773
rect 12157 20770 12223 20773
rect 6453 20768 12223 20770
rect 6453 20712 6458 20768
rect 6514 20712 12162 20768
rect 12218 20712 12223 20768
rect 6453 20710 12223 20712
rect 6453 20707 6519 20710
rect 12157 20707 12223 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 8109 20634 8175 20637
rect 8569 20634 8635 20637
rect 14549 20634 14615 20637
rect 8109 20632 14615 20634
rect 8109 20576 8114 20632
rect 8170 20576 8574 20632
rect 8630 20576 14554 20632
rect 14610 20576 14615 20632
rect 8109 20574 14615 20576
rect 8109 20571 8175 20574
rect 8569 20571 8635 20574
rect 14549 20571 14615 20574
rect 10777 20498 10843 20501
rect 13905 20498 13971 20501
rect 10777 20496 13971 20498
rect 10777 20440 10782 20496
rect 10838 20440 13910 20496
rect 13966 20440 13971 20496
rect 10777 20438 13971 20440
rect 10777 20435 10843 20438
rect 13905 20435 13971 20438
rect 0 20362 480 20392
rect 3325 20362 3391 20365
rect 0 20360 3391 20362
rect 0 20304 3330 20360
rect 3386 20304 3391 20360
rect 0 20302 3391 20304
rect 0 20272 480 20302
rect 3325 20299 3391 20302
rect 5441 20362 5507 20365
rect 12525 20362 12591 20365
rect 5441 20360 12591 20362
rect 5441 20304 5446 20360
rect 5502 20304 12530 20360
rect 12586 20304 12591 20360
rect 5441 20302 12591 20304
rect 5441 20299 5507 20302
rect 12525 20299 12591 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19682 480 19712
rect 1577 19682 1643 19685
rect 0 19680 1643 19682
rect 0 19624 1582 19680
rect 1638 19624 1643 19680
rect 0 19622 1643 19624
rect 0 19592 480 19622
rect 1577 19619 1643 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 9673 19410 9739 19413
rect 15285 19410 15351 19413
rect 9673 19408 15351 19410
rect 9673 19352 9678 19408
rect 9734 19352 15290 19408
rect 15346 19352 15351 19408
rect 9673 19350 15351 19352
rect 9673 19347 9739 19350
rect 15285 19347 15351 19350
rect 4061 19274 4127 19277
rect 15101 19274 15167 19277
rect 4061 19272 15167 19274
rect 4061 19216 4066 19272
rect 4122 19216 15106 19272
rect 15162 19216 15167 19272
rect 4061 19214 15167 19216
rect 4061 19211 4127 19214
rect 15101 19211 15167 19214
rect 0 19138 480 19168
rect 2497 19138 2563 19141
rect 0 19136 2563 19138
rect 0 19080 2502 19136
rect 2558 19080 2563 19136
rect 0 19078 2563 19080
rect 0 19048 480 19078
rect 2497 19075 2563 19078
rect 2681 19138 2747 19141
rect 4153 19138 4219 19141
rect 2681 19136 4219 19138
rect 2681 19080 2686 19136
rect 2742 19080 4158 19136
rect 4214 19080 4219 19136
rect 2681 19078 4219 19080
rect 2681 19075 2747 19078
rect 4153 19075 4219 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 9622 18940 9628 19004
rect 9692 19002 9698 19004
rect 9765 19002 9831 19005
rect 9692 19000 9831 19002
rect 9692 18944 9770 19000
rect 9826 18944 9831 19000
rect 9692 18942 9831 18944
rect 9692 18940 9698 18942
rect 9765 18939 9831 18942
rect 8109 18866 8175 18869
rect 13997 18866 14063 18869
rect 8109 18864 14063 18866
rect 8109 18808 8114 18864
rect 8170 18808 14002 18864
rect 14058 18808 14063 18864
rect 8109 18806 14063 18808
rect 8109 18803 8175 18806
rect 13997 18803 14063 18806
rect 7557 18730 7623 18733
rect 13353 18730 13419 18733
rect 7557 18728 13419 18730
rect 7557 18672 7562 18728
rect 7618 18672 13358 18728
rect 13414 18672 13419 18728
rect 7557 18670 13419 18672
rect 7557 18667 7623 18670
rect 13353 18667 13419 18670
rect 0 18594 480 18624
rect 4245 18594 4311 18597
rect 0 18592 4311 18594
rect 0 18536 4250 18592
rect 4306 18536 4311 18592
rect 0 18534 4311 18536
rect 0 18504 480 18534
rect 4245 18531 4311 18534
rect 7557 18594 7623 18597
rect 9949 18594 10015 18597
rect 7557 18592 10015 18594
rect 7557 18536 7562 18592
rect 7618 18536 9954 18592
rect 10010 18536 10015 18592
rect 7557 18534 10015 18536
rect 7557 18531 7623 18534
rect 9949 18531 10015 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 2865 18322 2931 18325
rect 4889 18322 4955 18325
rect 14917 18322 14983 18325
rect 2865 18320 14983 18322
rect 2865 18264 2870 18320
rect 2926 18264 4894 18320
rect 4950 18264 14922 18320
rect 14978 18264 14983 18320
rect 2865 18262 14983 18264
rect 2865 18259 2931 18262
rect 4889 18259 4955 18262
rect 14917 18259 14983 18262
rect 5073 18186 5139 18189
rect 16297 18186 16363 18189
rect 5073 18184 16363 18186
rect 5073 18128 5078 18184
rect 5134 18128 16302 18184
rect 16358 18128 16363 18184
rect 5073 18126 16363 18128
rect 5073 18123 5139 18126
rect 16297 18123 16363 18126
rect 16481 18186 16547 18189
rect 26509 18186 26575 18189
rect 16481 18184 26575 18186
rect 16481 18128 16486 18184
rect 16542 18128 26514 18184
rect 26570 18128 26575 18184
rect 16481 18126 26575 18128
rect 16481 18123 16547 18126
rect 26509 18123 26575 18126
rect 0 18050 480 18080
rect 13445 18050 13511 18053
rect 15285 18050 15351 18053
rect 0 17990 1410 18050
rect 0 17960 480 17990
rect 1350 17914 1410 17990
rect 13445 18048 15351 18050
rect 13445 17992 13450 18048
rect 13506 17992 15290 18048
rect 15346 17992 15351 18048
rect 13445 17990 15351 17992
rect 13445 17987 13511 17990
rect 15285 17987 15351 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 1485 17914 1551 17917
rect 1350 17912 1551 17914
rect 1350 17856 1490 17912
rect 1546 17856 1551 17912
rect 1350 17854 1551 17856
rect 1485 17851 1551 17854
rect 3877 17914 3943 17917
rect 9857 17914 9923 17917
rect 3877 17912 9923 17914
rect 3877 17856 3882 17912
rect 3938 17856 9862 17912
rect 9918 17856 9923 17912
rect 3877 17854 9923 17856
rect 3877 17851 3943 17854
rect 9857 17851 9923 17854
rect 13169 17914 13235 17917
rect 17861 17914 17927 17917
rect 13169 17912 17927 17914
rect 13169 17856 13174 17912
rect 13230 17856 17866 17912
rect 17922 17856 17927 17912
rect 13169 17854 17927 17856
rect 13169 17851 13235 17854
rect 17861 17851 17927 17854
rect 8017 17778 8083 17781
rect 15837 17778 15903 17781
rect 8017 17776 15903 17778
rect 8017 17720 8022 17776
rect 8078 17720 15842 17776
rect 15898 17720 15903 17776
rect 8017 17718 15903 17720
rect 8017 17715 8083 17718
rect 15837 17715 15903 17718
rect 3509 17642 3575 17645
rect 8385 17642 8451 17645
rect 3509 17640 8451 17642
rect 3509 17584 3514 17640
rect 3570 17584 8390 17640
rect 8446 17584 8451 17640
rect 3509 17582 8451 17584
rect 3509 17579 3575 17582
rect 8385 17579 8451 17582
rect 13077 17642 13143 17645
rect 23657 17642 23723 17645
rect 13077 17640 23723 17642
rect 13077 17584 13082 17640
rect 13138 17584 23662 17640
rect 23718 17584 23723 17640
rect 13077 17582 23723 17584
rect 13077 17579 13143 17582
rect 23657 17579 23723 17582
rect 0 17506 480 17536
rect 1669 17506 1735 17509
rect 0 17504 1735 17506
rect 0 17448 1674 17504
rect 1730 17448 1735 17504
rect 0 17446 1735 17448
rect 0 17416 480 17446
rect 1669 17443 1735 17446
rect 15653 17506 15719 17509
rect 18045 17506 18111 17509
rect 15653 17504 18111 17506
rect 15653 17448 15658 17504
rect 15714 17448 18050 17504
rect 18106 17448 18111 17504
rect 15653 17446 18111 17448
rect 15653 17443 15719 17446
rect 18045 17443 18111 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 7925 17234 7991 17237
rect 9673 17234 9739 17237
rect 7925 17232 9739 17234
rect 7925 17176 7930 17232
rect 7986 17176 9678 17232
rect 9734 17176 9739 17232
rect 7925 17174 9739 17176
rect 7925 17171 7991 17174
rect 9673 17171 9739 17174
rect 11053 17098 11119 17101
rect 1350 17096 11119 17098
rect 1350 17040 11058 17096
rect 11114 17040 11119 17096
rect 1350 17038 11119 17040
rect 0 16826 480 16856
rect 1350 16826 1410 17038
rect 11053 17035 11119 17038
rect 2681 16962 2747 16965
rect 6177 16962 6243 16965
rect 6453 16962 6519 16965
rect 2681 16960 6519 16962
rect 2681 16904 2686 16960
rect 2742 16904 6182 16960
rect 6238 16904 6458 16960
rect 6514 16904 6519 16960
rect 2681 16902 6519 16904
rect 2681 16899 2747 16902
rect 6177 16899 6243 16902
rect 6453 16899 6519 16902
rect 13077 16962 13143 16965
rect 16573 16962 16639 16965
rect 13077 16960 16639 16962
rect 13077 16904 13082 16960
rect 13138 16904 16578 16960
rect 16634 16904 16639 16960
rect 13077 16902 16639 16904
rect 13077 16899 13143 16902
rect 16573 16899 16639 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16766 1410 16826
rect 5073 16826 5139 16829
rect 7373 16826 7439 16829
rect 5073 16824 7439 16826
rect 5073 16768 5078 16824
rect 5134 16768 7378 16824
rect 7434 16768 7439 16824
rect 5073 16766 7439 16768
rect 0 16736 480 16766
rect 5073 16763 5139 16766
rect 7373 16763 7439 16766
rect 11421 16826 11487 16829
rect 17953 16826 18019 16829
rect 11421 16824 18019 16826
rect 11421 16768 11426 16824
rect 11482 16768 17958 16824
rect 18014 16768 18019 16824
rect 11421 16766 18019 16768
rect 11421 16763 11487 16766
rect 17953 16763 18019 16766
rect 11697 16690 11763 16693
rect 19149 16690 19215 16693
rect 11697 16688 19215 16690
rect 11697 16632 11702 16688
rect 11758 16632 19154 16688
rect 19210 16632 19215 16688
rect 11697 16630 19215 16632
rect 11697 16627 11763 16630
rect 19149 16627 19215 16630
rect 1761 16554 1827 16557
rect 2681 16554 2747 16557
rect 1761 16552 2747 16554
rect 1761 16496 1766 16552
rect 1822 16496 2686 16552
rect 2742 16496 2747 16552
rect 1761 16494 2747 16496
rect 1761 16491 1827 16494
rect 2681 16491 2747 16494
rect 2957 16554 3023 16557
rect 6269 16554 6335 16557
rect 2957 16552 6335 16554
rect 2957 16496 2962 16552
rect 3018 16496 6274 16552
rect 6330 16496 6335 16552
rect 2957 16494 6335 16496
rect 2957 16491 3023 16494
rect 6269 16491 6335 16494
rect 10041 16554 10107 16557
rect 13997 16554 14063 16557
rect 19425 16554 19491 16557
rect 10041 16552 13922 16554
rect 10041 16496 10046 16552
rect 10102 16496 13922 16552
rect 10041 16494 13922 16496
rect 10041 16491 10107 16494
rect 7005 16418 7071 16421
rect 11605 16418 11671 16421
rect 7005 16416 11671 16418
rect 7005 16360 7010 16416
rect 7066 16360 11610 16416
rect 11666 16360 11671 16416
rect 7005 16358 11671 16360
rect 13862 16418 13922 16494
rect 13997 16552 19491 16554
rect 13997 16496 14002 16552
rect 14058 16496 19430 16552
rect 19486 16496 19491 16552
rect 13997 16494 19491 16496
rect 13997 16491 14063 16494
rect 19425 16491 19491 16494
rect 14733 16418 14799 16421
rect 13862 16416 14799 16418
rect 13862 16360 14738 16416
rect 14794 16360 14799 16416
rect 13862 16358 14799 16360
rect 7005 16355 7071 16358
rect 11605 16355 11671 16358
rect 14733 16355 14799 16358
rect 15377 16418 15443 16421
rect 19057 16418 19123 16421
rect 15377 16416 19123 16418
rect 15377 16360 15382 16416
rect 15438 16360 19062 16416
rect 19118 16360 19123 16416
rect 15377 16358 19123 16360
rect 15377 16355 15443 16358
rect 19057 16355 19123 16358
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 7557 16282 7623 16285
rect 14641 16282 14707 16285
rect 0 16222 5458 16282
rect 0 16192 480 16222
rect 2037 16146 2103 16149
rect 3785 16146 3851 16149
rect 4337 16146 4403 16149
rect 2037 16144 4403 16146
rect 2037 16088 2042 16144
rect 2098 16088 3790 16144
rect 3846 16088 4342 16144
rect 4398 16088 4403 16144
rect 2037 16086 4403 16088
rect 5398 16146 5458 16222
rect 7557 16280 14707 16282
rect 7557 16224 7562 16280
rect 7618 16224 14646 16280
rect 14702 16224 14707 16280
rect 7557 16222 14707 16224
rect 7557 16219 7623 16222
rect 14641 16219 14707 16222
rect 20621 16282 20687 16285
rect 22093 16282 22159 16285
rect 20621 16280 22159 16282
rect 20621 16224 20626 16280
rect 20682 16224 22098 16280
rect 22154 16224 22159 16280
rect 20621 16222 22159 16224
rect 20621 16219 20687 16222
rect 22093 16219 22159 16222
rect 10961 16146 11027 16149
rect 5398 16144 11027 16146
rect 5398 16088 10966 16144
rect 11022 16088 11027 16144
rect 5398 16086 11027 16088
rect 2037 16083 2103 16086
rect 3785 16083 3851 16086
rect 4337 16083 4403 16086
rect 10961 16083 11027 16086
rect 14917 16146 14983 16149
rect 18045 16146 18111 16149
rect 14917 16144 18111 16146
rect 14917 16088 14922 16144
rect 14978 16088 18050 16144
rect 18106 16088 18111 16144
rect 14917 16086 18111 16088
rect 14917 16083 14983 16086
rect 18045 16083 18111 16086
rect 2129 16010 2195 16013
rect 9489 16010 9555 16013
rect 18045 16010 18111 16013
rect 2129 16008 6746 16010
rect 2129 15952 2134 16008
rect 2190 15952 6746 16008
rect 2129 15950 6746 15952
rect 2129 15947 2195 15950
rect 1669 15874 1735 15877
rect 5165 15874 5231 15877
rect 5390 15874 5396 15876
rect 1669 15872 5090 15874
rect 1669 15816 1674 15872
rect 1730 15816 5090 15872
rect 1669 15814 5090 15816
rect 1669 15811 1735 15814
rect 0 15738 480 15768
rect 5030 15738 5090 15814
rect 5165 15872 5396 15874
rect 5165 15816 5170 15872
rect 5226 15816 5396 15872
rect 5165 15814 5396 15816
rect 5165 15811 5231 15814
rect 5390 15812 5396 15814
rect 5460 15812 5466 15876
rect 6686 15874 6746 15950
rect 9489 16008 18111 16010
rect 9489 15952 9494 16008
rect 9550 15952 18050 16008
rect 18106 15952 18111 16008
rect 9489 15950 18111 15952
rect 9489 15947 9555 15950
rect 18045 15947 18111 15950
rect 9765 15874 9831 15877
rect 6686 15872 9831 15874
rect 6686 15816 9770 15872
rect 9826 15816 9831 15872
rect 6686 15814 9831 15816
rect 9765 15811 9831 15814
rect 10961 15874 11027 15877
rect 13997 15874 14063 15877
rect 10961 15872 14063 15874
rect 10961 15816 10966 15872
rect 11022 15816 14002 15872
rect 14058 15816 14063 15872
rect 10961 15814 14063 15816
rect 10961 15811 11027 15814
rect 13997 15811 14063 15814
rect 14181 15874 14247 15877
rect 18229 15874 18295 15877
rect 14181 15872 18295 15874
rect 14181 15816 14186 15872
rect 14242 15816 18234 15872
rect 18290 15816 18295 15872
rect 14181 15814 18295 15816
rect 14181 15811 14247 15814
rect 18229 15811 18295 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 7557 15738 7623 15741
rect 0 15678 4170 15738
rect 5030 15736 7623 15738
rect 5030 15680 7562 15736
rect 7618 15680 7623 15736
rect 5030 15678 7623 15680
rect 0 15648 480 15678
rect 4110 15466 4170 15678
rect 7557 15675 7623 15678
rect 15285 15738 15351 15741
rect 15510 15738 15516 15740
rect 15285 15736 15516 15738
rect 15285 15680 15290 15736
rect 15346 15680 15516 15736
rect 15285 15678 15516 15680
rect 15285 15675 15351 15678
rect 15510 15676 15516 15678
rect 15580 15676 15586 15740
rect 4245 15602 4311 15605
rect 7557 15602 7623 15605
rect 4245 15600 7623 15602
rect 4245 15544 4250 15600
rect 4306 15544 7562 15600
rect 7618 15544 7623 15600
rect 4245 15542 7623 15544
rect 4245 15539 4311 15542
rect 7557 15539 7623 15542
rect 10685 15602 10751 15605
rect 19241 15602 19307 15605
rect 10685 15600 19307 15602
rect 10685 15544 10690 15600
rect 10746 15544 19246 15600
rect 19302 15544 19307 15600
rect 10685 15542 19307 15544
rect 10685 15539 10751 15542
rect 19241 15539 19307 15542
rect 11237 15466 11303 15469
rect 4110 15464 11303 15466
rect 4110 15408 11242 15464
rect 11298 15408 11303 15464
rect 4110 15406 11303 15408
rect 11237 15403 11303 15406
rect 12801 15466 12867 15469
rect 19425 15466 19491 15469
rect 12801 15464 19491 15466
rect 12801 15408 12806 15464
rect 12862 15408 19430 15464
rect 19486 15408 19491 15464
rect 12801 15406 19491 15408
rect 12801 15403 12867 15406
rect 19425 15403 19491 15406
rect 1853 15330 1919 15333
rect 4245 15330 4311 15333
rect 1853 15328 4311 15330
rect 1853 15272 1858 15328
rect 1914 15272 4250 15328
rect 4306 15272 4311 15328
rect 1853 15270 4311 15272
rect 1853 15267 1919 15270
rect 4245 15267 4311 15270
rect 7373 15330 7439 15333
rect 7373 15328 14842 15330
rect 7373 15272 7378 15328
rect 7434 15272 14842 15328
rect 7373 15270 14842 15272
rect 7373 15267 7439 15270
rect 5610 15264 5930 15265
rect 0 15194 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 7833 15194 7899 15197
rect 11697 15194 11763 15197
rect 0 15134 2698 15194
rect 0 15104 480 15134
rect 2638 15092 2698 15134
rect 7833 15192 11763 15194
rect 7833 15136 7838 15192
rect 7894 15136 11702 15192
rect 11758 15136 11763 15192
rect 7833 15134 11763 15136
rect 7833 15131 7899 15134
rect 11697 15131 11763 15134
rect 2638 15058 2882 15092
rect 9673 15058 9739 15061
rect 2638 15056 9739 15058
rect 2638 15032 9678 15056
rect 2822 15000 9678 15032
rect 9734 15000 9739 15056
rect 2822 14998 9739 15000
rect 14782 15058 14842 15270
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 15193 15058 15259 15061
rect 14782 15056 15259 15058
rect 14782 15000 15198 15056
rect 15254 15000 15259 15056
rect 14782 14998 15259 15000
rect 9673 14995 9739 14998
rect 15193 14995 15259 14998
rect 15377 15058 15443 15061
rect 18873 15058 18939 15061
rect 15377 15056 18939 15058
rect 15377 15000 15382 15056
rect 15438 15000 18878 15056
rect 18934 15000 18939 15056
rect 15377 14998 18939 15000
rect 15377 14995 15443 14998
rect 18873 14995 18939 14998
rect 197 14922 263 14925
rect 4521 14922 4587 14925
rect 197 14920 4587 14922
rect 197 14864 202 14920
rect 258 14864 4526 14920
rect 4582 14864 4587 14920
rect 197 14862 4587 14864
rect 197 14859 263 14862
rect 4521 14859 4587 14862
rect 16389 14922 16455 14925
rect 23289 14922 23355 14925
rect 16389 14920 23355 14922
rect 16389 14864 16394 14920
rect 16450 14864 23294 14920
rect 23350 14864 23355 14920
rect 16389 14862 23355 14864
rect 16389 14859 16455 14862
rect 23289 14859 23355 14862
rect 12065 14786 12131 14789
rect 13077 14786 13143 14789
rect 15285 14786 15351 14789
rect 12065 14784 15351 14786
rect 12065 14728 12070 14784
rect 12126 14728 13082 14784
rect 13138 14728 15290 14784
rect 15346 14728 15351 14784
rect 12065 14726 15351 14728
rect 12065 14723 12131 14726
rect 13077 14723 13143 14726
rect 15285 14723 15351 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 480 14590
rect 1669 14587 1735 14590
rect 3601 14650 3667 14653
rect 10041 14650 10107 14653
rect 3601 14648 10107 14650
rect 3601 14592 3606 14648
rect 3662 14592 10046 14648
rect 10102 14592 10107 14648
rect 3601 14590 10107 14592
rect 3601 14587 3667 14590
rect 10041 14587 10107 14590
rect 12893 14650 12959 14653
rect 15653 14650 15719 14653
rect 12893 14648 15719 14650
rect 12893 14592 12898 14648
rect 12954 14592 15658 14648
rect 15714 14592 15719 14648
rect 12893 14590 15719 14592
rect 12893 14587 12959 14590
rect 15653 14587 15719 14590
rect 2405 14514 2471 14517
rect 4797 14514 4863 14517
rect 2405 14512 4863 14514
rect 2405 14456 2410 14512
rect 2466 14456 4802 14512
rect 4858 14456 4863 14512
rect 2405 14454 4863 14456
rect 2405 14451 2471 14454
rect 4797 14451 4863 14454
rect 5993 14514 6059 14517
rect 8385 14514 8451 14517
rect 5993 14512 8451 14514
rect 5993 14456 5998 14512
rect 6054 14456 8390 14512
rect 8446 14456 8451 14512
rect 5993 14454 8451 14456
rect 5993 14451 6059 14454
rect 8385 14451 8451 14454
rect 9622 14452 9628 14516
rect 9692 14514 9698 14516
rect 9765 14514 9831 14517
rect 9692 14512 9831 14514
rect 9692 14456 9770 14512
rect 9826 14456 9831 14512
rect 9692 14454 9831 14456
rect 9692 14452 9698 14454
rect 9765 14451 9831 14454
rect 3693 14378 3759 14381
rect 10317 14378 10383 14381
rect 3693 14376 10383 14378
rect 3693 14320 3698 14376
rect 3754 14320 10322 14376
rect 10378 14320 10383 14376
rect 3693 14318 10383 14320
rect 3693 14315 3759 14318
rect 10317 14315 10383 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13970 480 14000
rect 5533 13970 5599 13973
rect 0 13968 5599 13970
rect 0 13912 5538 13968
rect 5594 13912 5599 13968
rect 0 13910 5599 13912
rect 0 13880 480 13910
rect 5533 13907 5599 13910
rect 4797 13834 4863 13837
rect 8293 13834 8359 13837
rect 4797 13832 8359 13834
rect 4797 13776 4802 13832
rect 4858 13776 8298 13832
rect 8354 13776 8359 13832
rect 4797 13774 8359 13776
rect 4797 13771 4863 13774
rect 8293 13771 8359 13774
rect 11421 13834 11487 13837
rect 13629 13834 13695 13837
rect 11421 13832 13695 13834
rect 11421 13776 11426 13832
rect 11482 13776 13634 13832
rect 13690 13776 13695 13832
rect 11421 13774 13695 13776
rect 11421 13771 11487 13774
rect 13629 13771 13695 13774
rect 14641 13834 14707 13837
rect 19425 13834 19491 13837
rect 14641 13832 19491 13834
rect 14641 13776 14646 13832
rect 14702 13776 19430 13832
rect 19486 13776 19491 13832
rect 14641 13774 19491 13776
rect 14641 13771 14707 13774
rect 19425 13771 19491 13774
rect 1393 13698 1459 13701
rect 4705 13698 4771 13701
rect 1393 13696 4771 13698
rect 1393 13640 1398 13696
rect 1454 13640 4710 13696
rect 4766 13640 4771 13696
rect 1393 13638 4771 13640
rect 1393 13635 1459 13638
rect 4705 13635 4771 13638
rect 6269 13698 6335 13701
rect 8569 13698 8635 13701
rect 6269 13696 8635 13698
rect 6269 13640 6274 13696
rect 6330 13640 8574 13696
rect 8630 13640 8635 13696
rect 6269 13638 8635 13640
rect 6269 13635 6335 13638
rect 8569 13635 8635 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 1853 13562 1919 13565
rect 5441 13562 5507 13565
rect 1853 13560 5507 13562
rect 1853 13504 1858 13560
rect 1914 13504 5446 13560
rect 5502 13504 5507 13560
rect 1853 13502 5507 13504
rect 1853 13499 1919 13502
rect 5441 13499 5507 13502
rect 7557 13562 7623 13565
rect 10133 13562 10199 13565
rect 7557 13560 10199 13562
rect 7557 13504 7562 13560
rect 7618 13504 10138 13560
rect 10194 13504 10199 13560
rect 7557 13502 10199 13504
rect 7557 13499 7623 13502
rect 10133 13499 10199 13502
rect 0 13426 480 13456
rect 7649 13426 7715 13429
rect 0 13424 7715 13426
rect 0 13368 7654 13424
rect 7710 13368 7715 13424
rect 0 13366 7715 13368
rect 0 13336 480 13366
rect 7649 13363 7715 13366
rect 2589 13290 2655 13293
rect 5993 13290 6059 13293
rect 2589 13288 6059 13290
rect 2589 13232 2594 13288
rect 2650 13232 5998 13288
rect 6054 13232 6059 13288
rect 2589 13230 6059 13232
rect 2589 13227 2655 13230
rect 5993 13227 6059 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6545 13018 6611 13021
rect 12157 13018 12223 13021
rect 6545 13016 12223 13018
rect 6545 12960 6550 13016
rect 6606 12960 12162 13016
rect 12218 12960 12223 13016
rect 6545 12958 12223 12960
rect 6545 12955 6611 12958
rect 12157 12955 12223 12958
rect 0 12882 480 12912
rect 4245 12882 4311 12885
rect 0 12880 4311 12882
rect 0 12824 4250 12880
rect 4306 12824 4311 12880
rect 0 12822 4311 12824
rect 0 12792 480 12822
rect 4245 12819 4311 12822
rect 5809 12882 5875 12885
rect 13353 12882 13419 12885
rect 5809 12880 13419 12882
rect 5809 12824 5814 12880
rect 5870 12824 13358 12880
rect 13414 12824 13419 12880
rect 5809 12822 13419 12824
rect 5809 12819 5875 12822
rect 13353 12819 13419 12822
rect 18045 12882 18111 12885
rect 22277 12882 22343 12885
rect 18045 12880 22343 12882
rect 18045 12824 18050 12880
rect 18106 12824 22282 12880
rect 22338 12824 22343 12880
rect 18045 12822 22343 12824
rect 18045 12819 18111 12822
rect 22277 12819 22343 12822
rect 3601 12746 3667 12749
rect 6545 12746 6611 12749
rect 3601 12744 6611 12746
rect 3601 12688 3606 12744
rect 3662 12688 6550 12744
rect 6606 12688 6611 12744
rect 3601 12686 6611 12688
rect 3601 12683 3667 12686
rect 6545 12683 6611 12686
rect 6821 12746 6887 12749
rect 20805 12746 20871 12749
rect 6821 12744 20871 12746
rect 6821 12688 6826 12744
rect 6882 12688 20810 12744
rect 20866 12688 20871 12744
rect 6821 12686 20871 12688
rect 6821 12683 6887 12686
rect 20805 12683 20871 12686
rect 4061 12610 4127 12613
rect 6177 12610 6243 12613
rect 4061 12608 6243 12610
rect 4061 12552 4066 12608
rect 4122 12552 6182 12608
rect 6238 12552 6243 12608
rect 4061 12550 6243 12552
rect 4061 12547 4127 12550
rect 6177 12547 6243 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 2681 12474 2747 12477
rect 7833 12474 7899 12477
rect 2681 12472 7899 12474
rect 2681 12416 2686 12472
rect 2742 12416 7838 12472
rect 7894 12416 7899 12472
rect 2681 12414 7899 12416
rect 2681 12411 2747 12414
rect 7833 12411 7899 12414
rect 16389 12474 16455 12477
rect 17033 12474 17099 12477
rect 17953 12474 18019 12477
rect 18137 12474 18203 12477
rect 16389 12472 18203 12474
rect 16389 12416 16394 12472
rect 16450 12416 17038 12472
rect 17094 12416 17958 12472
rect 18014 12416 18142 12472
rect 18198 12416 18203 12472
rect 16389 12414 18203 12416
rect 16389 12411 16455 12414
rect 17033 12411 17099 12414
rect 17953 12411 18019 12414
rect 18137 12411 18203 12414
rect 0 12338 480 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 480 12278
rect 1577 12275 1643 12278
rect 5257 12338 5323 12341
rect 5717 12338 5783 12341
rect 5257 12336 5783 12338
rect 5257 12280 5262 12336
rect 5318 12280 5722 12336
rect 5778 12280 5783 12336
rect 5257 12278 5783 12280
rect 5257 12275 5323 12278
rect 5717 12275 5783 12278
rect 6361 12338 6427 12341
rect 10133 12338 10199 12341
rect 6361 12336 10199 12338
rect 6361 12280 6366 12336
rect 6422 12280 10138 12336
rect 10194 12280 10199 12336
rect 6361 12278 10199 12280
rect 6361 12275 6427 12278
rect 10133 12275 10199 12278
rect 11237 12338 11303 12341
rect 21081 12338 21147 12341
rect 11237 12336 21147 12338
rect 11237 12280 11242 12336
rect 11298 12280 21086 12336
rect 21142 12280 21147 12336
rect 11237 12278 21147 12280
rect 11237 12275 11303 12278
rect 21081 12275 21147 12278
rect 5165 12202 5231 12205
rect 7189 12202 7255 12205
rect 7741 12202 7807 12205
rect 20897 12202 20963 12205
rect 5165 12200 7807 12202
rect 5165 12144 5170 12200
rect 5226 12144 7194 12200
rect 7250 12144 7746 12200
rect 7802 12144 7807 12200
rect 5165 12142 7807 12144
rect 5165 12139 5231 12142
rect 7189 12139 7255 12142
rect 7741 12139 7807 12142
rect 13494 12200 20963 12202
rect 13494 12144 20902 12200
rect 20958 12144 20963 12200
rect 13494 12142 20963 12144
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 0 11794 480 11824
rect 3969 11794 4035 11797
rect 0 11792 4035 11794
rect 0 11736 3974 11792
rect 4030 11736 4035 11792
rect 0 11734 4035 11736
rect 0 11704 480 11734
rect 3969 11731 4035 11734
rect 7925 11794 7991 11797
rect 13494 11794 13554 12142
rect 20897 12139 20963 12142
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 7925 11792 13554 11794
rect 7925 11736 7930 11792
rect 7986 11736 13554 11792
rect 7925 11734 13554 11736
rect 13629 11794 13695 11797
rect 18505 11794 18571 11797
rect 13629 11792 18571 11794
rect 13629 11736 13634 11792
rect 13690 11736 18510 11792
rect 18566 11736 18571 11792
rect 13629 11734 18571 11736
rect 7925 11731 7991 11734
rect 13629 11731 13695 11734
rect 18505 11731 18571 11734
rect 3417 11658 3483 11661
rect 6545 11658 6611 11661
rect 3417 11656 6611 11658
rect 3417 11600 3422 11656
rect 3478 11600 6550 11656
rect 6606 11600 6611 11656
rect 3417 11598 6611 11600
rect 3417 11595 3483 11598
rect 6545 11595 6611 11598
rect 6729 11522 6795 11525
rect 8385 11522 8451 11525
rect 6729 11520 8451 11522
rect 6729 11464 6734 11520
rect 6790 11464 8390 11520
rect 8446 11464 8451 11520
rect 6729 11462 8451 11464
rect 6729 11459 6795 11462
rect 8385 11459 8451 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3509 11386 3575 11389
rect 6637 11386 6703 11389
rect 3509 11384 6703 11386
rect 3509 11328 3514 11384
rect 3570 11328 6642 11384
rect 6698 11328 6703 11384
rect 3509 11326 6703 11328
rect 3509 11323 3575 11326
rect 6637 11323 6703 11326
rect 2221 11250 2287 11253
rect 4521 11250 4587 11253
rect 2221 11248 4587 11250
rect 2221 11192 2226 11248
rect 2282 11192 4526 11248
rect 4582 11192 4587 11248
rect 2221 11190 4587 11192
rect 2221 11187 2287 11190
rect 4521 11187 4587 11190
rect 13353 11250 13419 11253
rect 21725 11250 21791 11253
rect 13353 11248 21791 11250
rect 13353 11192 13358 11248
rect 13414 11192 21730 11248
rect 21786 11192 21791 11248
rect 13353 11190 21791 11192
rect 13353 11187 13419 11190
rect 21725 11187 21791 11190
rect 0 11114 480 11144
rect 2865 11114 2931 11117
rect 0 11112 2931 11114
rect 0 11056 2870 11112
rect 2926 11056 2931 11112
rect 0 11054 2931 11056
rect 0 11024 480 11054
rect 2865 11051 2931 11054
rect 4061 11114 4127 11117
rect 15469 11114 15535 11117
rect 4061 11112 15535 11114
rect 4061 11056 4066 11112
rect 4122 11056 15474 11112
rect 15530 11056 15535 11112
rect 4061 11054 15535 11056
rect 4061 11051 4127 11054
rect 15469 11051 15535 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 1761 10706 1827 10709
rect 16757 10706 16823 10709
rect 1761 10704 16823 10706
rect 1761 10648 1766 10704
rect 1822 10648 16762 10704
rect 16818 10648 16823 10704
rect 1761 10646 16823 10648
rect 1761 10643 1827 10646
rect 16757 10643 16823 10646
rect 0 10570 480 10600
rect 1853 10570 1919 10573
rect 0 10568 1919 10570
rect 0 10512 1858 10568
rect 1914 10512 1919 10568
rect 0 10510 1919 10512
rect 0 10480 480 10510
rect 1853 10507 1919 10510
rect 10041 10434 10107 10437
rect 9998 10432 10107 10434
rect 9998 10376 10046 10432
rect 10102 10376 10107 10432
rect 9998 10371 10107 10376
rect 13445 10434 13511 10437
rect 15653 10434 15719 10437
rect 13445 10432 15719 10434
rect 13445 10376 13450 10432
rect 13506 10376 15658 10432
rect 15714 10376 15719 10432
rect 13445 10374 15719 10376
rect 13445 10371 13511 10374
rect 15653 10371 15719 10374
rect 2405 10298 2471 10301
rect 4153 10298 4219 10301
rect 2405 10296 4219 10298
rect 2405 10240 2410 10296
rect 2466 10240 4158 10296
rect 4214 10240 4219 10296
rect 2405 10238 4219 10240
rect 2405 10235 2471 10238
rect 4153 10235 4219 10238
rect 9622 10100 9628 10164
rect 9692 10162 9698 10164
rect 9857 10162 9923 10165
rect 9692 10160 9923 10162
rect 9692 10104 9862 10160
rect 9918 10104 9923 10160
rect 9692 10102 9923 10104
rect 9998 10162 10058 10371
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 10317 10162 10383 10165
rect 9998 10160 10383 10162
rect 9998 10104 10322 10160
rect 10378 10104 10383 10160
rect 9998 10102 10383 10104
rect 9692 10100 9698 10102
rect 9857 10099 9923 10102
rect 10317 10099 10383 10102
rect 0 10026 480 10056
rect 2405 10026 2471 10029
rect 2865 10026 2931 10029
rect 0 10024 2931 10026
rect 0 9968 2410 10024
rect 2466 9968 2870 10024
rect 2926 9968 2931 10024
rect 0 9966 2931 9968
rect 0 9936 480 9966
rect 2405 9963 2471 9966
rect 2865 9963 2931 9966
rect 7649 10026 7715 10029
rect 18137 10026 18203 10029
rect 7649 10024 18203 10026
rect 7649 9968 7654 10024
rect 7710 9968 18142 10024
rect 18198 9968 18203 10024
rect 7649 9966 18203 9968
rect 7649 9963 7715 9966
rect 18137 9963 18203 9966
rect 9857 9890 9923 9893
rect 11145 9890 11211 9893
rect 9857 9888 11211 9890
rect 9857 9832 9862 9888
rect 9918 9832 11150 9888
rect 11206 9832 11211 9888
rect 9857 9830 11211 9832
rect 9857 9827 9923 9830
rect 11145 9827 11211 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 9029 9754 9095 9757
rect 9622 9754 9628 9756
rect 9029 9752 9628 9754
rect 9029 9696 9034 9752
rect 9090 9696 9628 9752
rect 9029 9694 9628 9696
rect 9029 9691 9095 9694
rect 9622 9692 9628 9694
rect 9692 9692 9698 9756
rect 10225 9754 10291 9757
rect 11237 9754 11303 9757
rect 10225 9752 11303 9754
rect 10225 9696 10230 9752
rect 10286 9696 11242 9752
rect 11298 9696 11303 9752
rect 10225 9694 11303 9696
rect 10225 9691 10291 9694
rect 11237 9691 11303 9694
rect 2957 9618 3023 9621
rect 9765 9618 9831 9621
rect 2957 9616 9831 9618
rect 2957 9560 2962 9616
rect 3018 9560 9770 9616
rect 9826 9560 9831 9616
rect 2957 9558 9831 9560
rect 2957 9555 3023 9558
rect 9765 9555 9831 9558
rect 0 9482 480 9512
rect 5349 9482 5415 9485
rect 0 9480 5415 9482
rect 0 9424 5354 9480
rect 5410 9424 5415 9480
rect 0 9422 5415 9424
rect 0 9392 480 9422
rect 5349 9419 5415 9422
rect 9581 9482 9647 9485
rect 12433 9482 12499 9485
rect 18045 9482 18111 9485
rect 9581 9480 10978 9482
rect 9581 9424 9586 9480
rect 9642 9424 10978 9480
rect 9581 9422 10978 9424
rect 9581 9419 9647 9422
rect 1393 9346 1459 9349
rect 10133 9346 10199 9349
rect 1393 9344 10199 9346
rect 1393 9288 1398 9344
rect 1454 9288 10138 9344
rect 10194 9288 10199 9344
rect 1393 9286 10199 9288
rect 10918 9346 10978 9422
rect 12433 9480 18111 9482
rect 12433 9424 12438 9480
rect 12494 9424 18050 9480
rect 18106 9424 18111 9480
rect 12433 9422 18111 9424
rect 12433 9419 12499 9422
rect 18045 9419 18111 9422
rect 16573 9346 16639 9349
rect 10918 9344 16639 9346
rect 10918 9288 16578 9344
rect 16634 9288 16639 9344
rect 10918 9286 16639 9288
rect 1393 9283 1459 9286
rect 10133 9283 10199 9286
rect 16573 9283 16639 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 4889 9210 4955 9213
rect 9857 9210 9923 9213
rect 4889 9208 9923 9210
rect 4889 9152 4894 9208
rect 4950 9152 9862 9208
rect 9918 9152 9923 9208
rect 4889 9150 9923 9152
rect 4889 9147 4955 9150
rect 9857 9147 9923 9150
rect 7833 9074 7899 9077
rect 2454 9072 7899 9074
rect 2454 9016 7838 9072
rect 7894 9016 7899 9072
rect 2454 9014 7899 9016
rect 0 8938 480 8968
rect 2454 8938 2514 9014
rect 7833 9011 7899 9014
rect 0 8878 2514 8938
rect 2681 8938 2747 8941
rect 4889 8938 4955 8941
rect 2681 8936 4955 8938
rect 2681 8880 2686 8936
rect 2742 8880 4894 8936
rect 4950 8880 4955 8936
rect 2681 8878 4955 8880
rect 0 8848 480 8878
rect 2681 8875 2747 8878
rect 4889 8875 4955 8878
rect 5073 8938 5139 8941
rect 8109 8938 8175 8941
rect 8937 8938 9003 8941
rect 5073 8936 9003 8938
rect 5073 8880 5078 8936
rect 5134 8880 8114 8936
rect 8170 8880 8942 8936
rect 8998 8880 9003 8936
rect 5073 8878 9003 8880
rect 5073 8875 5139 8878
rect 8109 8875 8175 8878
rect 8937 8875 9003 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 10593 8530 10659 8533
rect 2454 8528 10659 8530
rect 2454 8472 10598 8528
rect 10654 8472 10659 8528
rect 2454 8470 10659 8472
rect 0 8258 480 8288
rect 2454 8258 2514 8470
rect 10593 8467 10659 8470
rect 2589 8394 2655 8397
rect 9765 8394 9831 8397
rect 2589 8392 9831 8394
rect 2589 8336 2594 8392
rect 2650 8336 9770 8392
rect 9826 8336 9831 8392
rect 2589 8334 9831 8336
rect 2589 8331 2655 8334
rect 9765 8331 9831 8334
rect 0 8198 2514 8258
rect 0 8168 480 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 4061 7986 4127 7989
rect 15561 7986 15627 7989
rect 4061 7984 15627 7986
rect 4061 7928 4066 7984
rect 4122 7928 15566 7984
rect 15622 7928 15627 7984
rect 4061 7926 15627 7928
rect 4061 7923 4127 7926
rect 15561 7923 15627 7926
rect 3969 7850 4035 7853
rect 11605 7850 11671 7853
rect 3969 7848 11671 7850
rect 3969 7792 3974 7848
rect 4030 7792 11610 7848
rect 11666 7792 11671 7848
rect 3969 7790 11671 7792
rect 3969 7787 4035 7790
rect 11605 7787 11671 7790
rect 0 7714 480 7744
rect 0 7654 2744 7714
rect 0 7624 480 7654
rect 2684 7578 2744 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 2684 7518 2882 7578
rect 2822 7442 2882 7518
rect 13445 7442 13511 7445
rect 2822 7440 13511 7442
rect 2822 7384 13450 7440
rect 13506 7384 13511 7440
rect 2822 7382 13511 7384
rect 13445 7379 13511 7382
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 14365 6898 14431 6901
rect 2592 6896 14431 6898
rect 2592 6840 14370 6896
rect 14426 6840 14431 6896
rect 2592 6838 14431 6840
rect 0 6626 480 6656
rect 2592 6626 2652 6838
rect 14365 6835 14431 6838
rect 0 6566 2652 6626
rect 0 6536 480 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6082 480 6112
rect 3601 6082 3667 6085
rect 0 6080 3667 6082
rect 0 6024 3606 6080
rect 3662 6024 3667 6080
rect 0 6022 3667 6024
rect 0 5992 480 6022
rect 3601 6019 3667 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 3693 5402 3759 5405
rect 0 5400 3759 5402
rect 0 5344 3698 5400
rect 3754 5344 3759 5400
rect 0 5342 3759 5344
rect 0 5312 480 5342
rect 3693 5339 3759 5342
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3417 4858 3483 4861
rect 0 4856 3483 4858
rect 0 4800 3422 4856
rect 3478 4800 3483 4856
rect 0 4798 3483 4800
rect 0 4768 480 4798
rect 3417 4795 3483 4798
rect 5610 4384 5930 4385
rect 0 4314 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 565 4314 631 4317
rect 0 4312 631 4314
rect 0 4256 570 4312
rect 626 4256 631 4312
rect 0 4254 631 4256
rect 0 4224 480 4254
rect 565 4251 631 4254
rect 9489 4042 9555 4045
rect 13905 4042 13971 4045
rect 9489 4040 13971 4042
rect 9489 3984 9494 4040
rect 9550 3984 13910 4040
rect 13966 3984 13971 4040
rect 9489 3982 13971 3984
rect 9489 3979 9555 3982
rect 13905 3979 13971 3982
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 3969 3770 4035 3773
rect 0 3768 4035 3770
rect 0 3712 3974 3768
rect 4030 3712 4035 3768
rect 0 3710 4035 3712
rect 0 3680 480 3710
rect 3969 3707 4035 3710
rect 11973 3498 12039 3501
rect 23197 3498 23263 3501
rect 11973 3496 23263 3498
rect 11973 3440 11978 3496
rect 12034 3440 23202 3496
rect 23258 3440 23263 3496
rect 11973 3438 23263 3440
rect 11973 3435 12039 3438
rect 23197 3435 23263 3438
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2681 3226 2747 3229
rect 0 3224 2747 3226
rect 0 3168 2686 3224
rect 2742 3168 2747 3224
rect 0 3166 2747 3168
rect 0 3136 480 3166
rect 2681 3163 2747 3166
rect 2773 2954 2839 2957
rect 13077 2954 13143 2957
rect 2773 2952 13143 2954
rect 2773 2896 2778 2952
rect 2834 2896 13082 2952
rect 13138 2896 13143 2952
rect 2773 2894 13143 2896
rect 2773 2891 2839 2894
rect 13077 2891 13143 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2546 480 2576
rect 933 2546 999 2549
rect 12617 2546 12683 2549
rect 0 2544 999 2546
rect 0 2488 938 2544
rect 994 2488 999 2544
rect 0 2486 999 2488
rect 0 2456 480 2486
rect 933 2483 999 2486
rect 1166 2544 12683 2546
rect 1166 2488 12622 2544
rect 12678 2488 12683 2544
rect 1166 2486 12683 2488
rect 1166 2138 1226 2486
rect 12617 2483 12683 2486
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 614 2078 1226 2138
rect 0 2002 480 2032
rect 614 2002 674 2078
rect 0 1942 674 2002
rect 0 1912 480 1942
rect 933 1730 999 1733
rect 16113 1730 16179 1733
rect 933 1728 16179 1730
rect 933 1672 938 1728
rect 994 1672 16118 1728
rect 16174 1672 16179 1728
rect 933 1670 16179 1672
rect 933 1667 999 1670
rect 16113 1667 16179 1670
rect 12065 1594 12131 1597
rect 614 1592 12131 1594
rect 614 1536 12070 1592
rect 12126 1536 12131 1592
rect 614 1534 12131 1536
rect 0 1458 480 1488
rect 614 1458 674 1534
rect 12065 1531 12131 1534
rect 0 1398 674 1458
rect 0 1368 480 1398
rect 9949 1322 10015 1325
rect 614 1320 10015 1322
rect 614 1264 9954 1320
rect 10010 1264 10015 1320
rect 614 1262 10015 1264
rect 0 914 480 944
rect 614 914 674 1262
rect 9949 1259 10015 1262
rect 0 854 674 914
rect 0 824 480 854
rect 0 370 480 400
rect 3049 370 3115 373
rect 0 368 3115 370
rect 0 312 3054 368
rect 3110 312 3115 368
rect 0 310 3115 312
rect 0 280 480 310
rect 3049 307 3115 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 9628 18940 9692 19004
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 5396 15812 5460 15876
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 15516 15676 15580 15740
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 9628 14452 9692 14516
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 9628 10100 9692 10164
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 9628 9692 9692 9756
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 9627 19004 9693 19005
rect 9627 18940 9628 19004
rect 9692 18940 9693 19004
rect 9627 18939 9693 18940
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5395 15812 5396 15862
rect 5460 15812 5461 15862
rect 5395 15811 5461 15812
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 9630 14517 9690 18939
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 9627 14516 9693 14517
rect 9627 14452 9628 14516
rect 9692 14452 9693 14516
rect 9627 14451 9693 14452
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9627 10164 9693 10165
rect 9627 10100 9628 10164
rect 9692 10100 9693 10164
rect 9627 10099 9693 10100
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 9630 9757 9690 10099
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 15518 15741 15578 15862
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 15515 15740 15581 15741
rect 15515 15676 15516 15740
rect 15580 15676 15581 15740
rect 15515 15675 15581 15676
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 5310 15876 5546 16098
rect 5310 15862 5396 15876
rect 5396 15862 5460 15876
rect 5460 15862 5546 15876
rect 15430 15862 15666 16098
<< metal5 >>
rect 5268 16098 15708 16140
rect 5268 15862 5310 16098
rect 5546 15862 15430 16098
rect 15666 15862 15708 16098
rect 5268 15820 15708 15862
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604666999
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604666999
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604666999
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604666999
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604666999
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604666999
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604666999
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604666999
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604666999
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604666999
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604666999
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604666999
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604666999
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604666999
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604666999
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604666999
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604666999
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604666999
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604666999
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604666999
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604666999
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604666999
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604666999
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604666999
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604666999
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604666999
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604666999
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604666999
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604666999
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604666999
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604666999
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604666999
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604666999
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604666999
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604666999
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604666999
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604666999
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604666999
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604666999
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604666999
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604666999
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604666999
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604666999
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604666999
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604666999
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604666999
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604666999
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604666999
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604666999
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_80
timestamp 1604666999
transform 1 0 8464 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1604666999
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604666999
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604666999
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604666999
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604666999
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604666999
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604666999
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604666999
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604666999
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604666999
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604666999
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604666999
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604666999
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 9200 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_107
timestamp 1604666999
transform 1 0 10948 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1604666999
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604666999
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604666999
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604666999
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604666999
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604666999
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604666999
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604666999
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604666999
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604666999
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604666999
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604666999
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604666999
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604666999
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604666999
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604666999
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604666999
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604666999
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604666999
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604666999
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604666999
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604666999
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604666999
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604666999
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604666999
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604666999
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604666999
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604666999
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604666999
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604666999
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604666999
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604666999
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604666999
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604666999
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604666999
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604666999
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604666999
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604666999
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604666999
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604666999
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604666999
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604666999
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604666999
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604666999
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604666999
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604666999
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604666999
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604666999
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604666999
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_7
timestamp 1604666999
transform 1 0 1748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1604666999
transform 1 0 2852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1604666999
transform 1 0 3956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1604666999
transform 1 0 5060 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_55
timestamp 1604666999
transform 1 0 6164 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604666999
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _037_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 9660 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_86
timestamp 1604666999
transform 1 0 9016 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1604666999
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1604666999
transform 1 0 9936 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1604666999
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_106
timestamp 1604666999
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1604666999
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604666999
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604666999
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604666999
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604666999
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604666999
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604666999
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604666999
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604666999
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604666999
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604666999
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604666999
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_6
timestamp 1604666999
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1604666999
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_14
timestamp 1604666999
transform 1 0 2392 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_26
timestamp 1604666999
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1604666999
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604666999
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_68
timestamp 1604666999
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_76
timestamp 1604666999
transform 1 0 8096 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1604666999
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp 1604666999
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10304 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1604666999
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_123
timestamp 1604666999
transform 1 0 12420 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_127
timestamp 1604666999
transform 1 0 12788 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_130
timestamp 1604666999
transform 1 0 13064 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_142
timestamp 1604666999
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1604666999
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604666999
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604666999
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604666999
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604666999
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604666999
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604666999
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604666999
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604666999
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp 1604666999
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1604666999
transform 1 0 2024 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_14
timestamp 1604666999
transform 1 0 2392 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_17
timestamp 1604666999
transform 1 0 2668 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_29
timestamp 1604666999
transform 1 0 3772 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1604666999
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1604666999
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_49
timestamp 1604666999
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604666999
transform 1 0 6900 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 7912 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1604666999
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1604666999
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1604666999
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1604666999
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604666999
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604666999
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604666999
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12880 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604666999
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1604666999
transform 1 0 15732 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1604666999
transform 1 0 16468 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_170
timestamp 1604666999
transform 1 0 16744 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604666999
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604666999
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604666999
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604666999
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604666999
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604666999
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604666999
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _083_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1604666999
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1604666999
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1604666999
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1604666999
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_26
timestamp 1604666999
transform 1 0 3496 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_36
timestamp 1604666999
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_40
timestamp 1604666999
transform 1 0 4784 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_52
timestamp 1604666999
transform 1 0 5888 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6624 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1604666999
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_83
timestamp 1604666999
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_87
timestamp 1604666999
transform 1 0 9108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11960 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1604666999
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_116
timestamp 1604666999
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12144 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_139
timestamp 1604666999
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1604666999
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_147
timestamp 1604666999
transform 1 0 14628 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1604666999
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_161
timestamp 1604666999
transform 1 0 15916 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1604666999
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_171
timestamp 1604666999
transform 1 0 16836 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_183
timestamp 1604666999
transform 1 0 17940 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_195
timestamp 1604666999
transform 1 0 19044 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_207
timestamp 1604666999
transform 1 0 20148 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1604666999
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604666999
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604666999
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604666999
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604666999
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1604666999
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604666999
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604666999
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1604666999
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604666999
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 1604666999
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2944 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp 1604666999
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_35
timestamp 1604666999
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 3956 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1604666999
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1604666999
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1604666999
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_43
timestamp 1604666999
transform 1 0 5060 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1604666999
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1604666999
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_65
timestamp 1604666999
transform 1 0 7084 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604666999
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604666999
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604666999
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_80
timestamp 1604666999
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1604666999
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_84
timestamp 1604666999
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_28.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9568 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_108
timestamp 1604666999
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1604666999
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1604666999
transform 1 0 10764 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1604666999
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604666999
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604666999
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_30.mux_l1_in_0_
timestamp 1604666999
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604666999
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1604666999
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1604666999
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_129
timestamp 1604666999
transform 1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604666999
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604666999
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_14_147
timestamp 1604666999
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1604666999
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_140
timestamp 1604666999
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1604666999
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14352 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604666999
transform 1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15732 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1604666999
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_167
timestamp 1604666999
transform 1 0 16468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_174
timestamp 1604666999
transform 1 0 17112 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_178
timestamp 1604666999
transform 1 0 17480 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_187
timestamp 1604666999
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1604666999
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18216 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1604666999
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_189
timestamp 1604666999
transform 1 0 18492 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_195
timestamp 1604666999
transform 1 0 19044 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_207
timestamp 1604666999
transform 1 0 20148 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1604666999
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604666999
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_219
timestamp 1604666999
transform 1 0 21252 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_231
timestamp 1604666999
transform 1 0 22356 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604666999
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1604666999
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604666999
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604666999
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604666999
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604666999
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604666999
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1564 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1604666999
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1604666999
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1604666999
transform 1 0 5796 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604666999
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7268 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9752 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1604666999
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1604666999
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1604666999
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_117
timestamp 1604666999
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15180 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_142
timestamp 1604666999
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_146
timestamp 1604666999
transform 1 0 14536 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1604666999
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16744 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604666999
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1604666999
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp 1604666999
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 1604666999
transform 1 0 17388 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604666999
transform 1 0 18308 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604666999
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604666999
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1604666999
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_195
timestamp 1604666999
transform 1 0 19044 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_207
timestamp 1604666999
transform 1 0 20148 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_219
timestamp 1604666999
transform 1 0 21252 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_231
timestamp 1604666999
transform 1 0 22356 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1604666999
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604666999
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604666999
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1604666999
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp 1604666999
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604666999
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6164 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1604666999
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1604666999
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_50
timestamp 1604666999
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_54
timestamp 1604666999
transform 1 0 6072 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_74
timestamp 1604666999
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_78
timestamp 1604666999
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1604666999
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1604666999
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604666999
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_98
timestamp 1604666999
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604666999
transform 1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10856 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1604666999
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_30.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1604666999
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1604666999
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1604666999
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1604666999
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604666999
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1604666999
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1604666999
transform 1 0 17388 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604666999
transform 1 0 17756 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1604666999
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_189
timestamp 1604666999
transform 1 0 18492 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1604666999
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604666999
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604666999
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604666999
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604666999
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604666999
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2024 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1604666999
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604666999
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_29
timestamp 1604666999
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1604666999
transform 1 0 4232 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1604666999
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604666999
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604666999
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1604666999
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_75
timestamp 1604666999
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8464 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1604666999
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604666999
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_103
timestamp 1604666999
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1604666999
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604666999
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604666999
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13248 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_128
timestamp 1604666999
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1604666999
transform 1 0 14996 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_155
timestamp 1604666999
transform 1 0 15364 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1604666999
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16008 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1604666999
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604666999
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1604666999
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_197
timestamp 1604666999
transform 1 0 19228 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_209
timestamp 1604666999
transform 1 0 20332 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1604666999
transform 1 0 21436 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_226
timestamp 1604666999
transform 1 0 21896 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_238
timestamp 1604666999
transform 1 0 23000 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604666999
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604666999
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1604666999
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1604666999
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1604666999
transform 1 0 3312 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1604666999
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1604666999
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5428 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1604666999
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_46
timestamp 1604666999
transform 1 0 5336 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 1604666999
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_70
timestamp 1604666999
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_83
timestamp 1604666999
transform 1 0 8740 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_87
timestamp 1604666999
transform 1 0 9108 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1604666999
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_28.mux_l2_in_0_
timestamp 1604666999
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_102
timestamp 1604666999
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1604666999
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_125
timestamp 1604666999
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_129
timestamp 1604666999
transform 1 0 12972 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1604666999
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 15640 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1604666999
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16652 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_161
timestamp 1604666999
transform 1 0 15916 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_165
timestamp 1604666999
transform 1 0 16284 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1604666999
transform 1 0 16560 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_188
timestamp 1604666999
transform 1 0 18400 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_200
timestamp 1604666999
transform 1 0 19504 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1604666999
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21712 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_223
timestamp 1604666999
transform 1 0 21620 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604666999
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604666999
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604666999
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604666999
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1604666999
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_7
timestamp 1604666999
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604666999
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1604666999
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 2576 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1604666999
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1604666999
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_20
timestamp 1604666999
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1604666999
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_35
timestamp 1604666999
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_49
timestamp 1604666999
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1604666999
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1604666999
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604666999
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604666999
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5888 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1604666999
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1604666999
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604666999
transform 1 0 7452 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_77
timestamp 1604666999
transform 1 0 8188 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_73
timestamp 1604666999
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_75
timestamp 1604666999
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1604666999
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604666999
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_84
timestamp 1604666999
transform 1 0 8832 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_84
timestamp 1604666999
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1604666999
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604666999
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_97
timestamp 1604666999
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1604666999
transform 1 0 11040 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604666999
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604666999
transform 1 0 10764 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1604666999
transform 1 0 11592 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_102
timestamp 1604666999
transform 1 0 10488 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11960 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604666999
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_136
timestamp 1604666999
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1604666999
transform 1 0 13708 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_142
timestamp 1604666999
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_150
timestamp 1604666999
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1604666999
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1604666999
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15548 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1604666999
transform 1 0 15732 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_163
timestamp 1604666999
transform 1 0 16100 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604666999
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_176
timestamp 1604666999
transform 1 0 17296 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18032 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1604666999
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_187
timestamp 1604666999
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_191
timestamp 1604666999
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_195
timestamp 1604666999
transform 1 0 19044 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_207
timestamp 1604666999
transform 1 0 20148 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_203
timestamp 1604666999
transform 1 0 19780 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1604666999
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_218
timestamp 1604666999
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_220
timestamp 1604666999
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_224
timestamp 1604666999
transform 1 0 21712 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_233
timestamp 1604666999
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_237
timestamp 1604666999
transform 1 0 22908 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_230
timestamp 1604666999
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_243
timestamp 1604666999
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604666999
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_242
timestamp 1604666999
transform 1 0 23368 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_254
timestamp 1604666999
transform 1 0 24472 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604666999
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_266
timestamp 1604666999
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1604666999
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604666999
transform 1 0 2760 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_7
timestamp 1604666999
transform 1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_11
timestamp 1604666999
transform 1 0 2116 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1604666999
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4324 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_31
timestamp 1604666999
transform 1 0 3956 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_34
timestamp 1604666999
transform 1 0 4232 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp 1604666999
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1604666999
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_52
timestamp 1604666999
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_56
timestamp 1604666999
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7544 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604666999
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1604666999
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1604666999
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9108 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1604666999
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1604666999
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1604666999
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604666999
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604666999
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13800 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_126
timestamp 1604666999
transform 1 0 12696 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1604666999
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1604666999
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_34.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16284 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1604666999
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_174
timestamp 1604666999
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1604666999
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604666999
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604666999
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604666999
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604666999
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604666999
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604666999
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604666999
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604666999
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1604666999
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1604666999
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604666999
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604666999
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6072 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604666999
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1604666999
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_45
timestamp 1604666999
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_49
timestamp 1604666999
transform 1 0 5612 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1604666999
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1604666999
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604666999
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_84
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1604666999
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11776 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1604666999
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_106
timestamp 1604666999
transform 1 0 10856 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1604666999
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1604666999
transform 1 0 13524 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1604666999
transform 1 0 14076 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604666999
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604666999
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1604666999
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1604666999
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_174
timestamp 1604666999
transform 1 0 17112 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_186
timestamp 1604666999
transform 1 0 18216 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_198
timestamp 1604666999
transform 1 0 19320 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1604666999
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604666999
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604666999
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604666999
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604666999
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2852 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1604666999
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1604666999
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp 1604666999
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1604666999
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604666999
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1604666999
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_50
timestamp 1604666999
transform 1 0 5704 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_54
timestamp 1604666999
transform 1 0 6072 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604666999
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 9752 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1604666999
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_85
timestamp 1604666999
transform 1 0 8924 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1604666999
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1604666999
transform 1 0 11500 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1604666999
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604666999
transform 1 0 12880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1604666999
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1604666999
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13892 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1604666999
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_34.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1604666999
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604666999
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604666999
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_196
timestamp 1604666999
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1604666999
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_206
timestamp 1604666999
transform 1 0 20056 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_218
timestamp 1604666999
transform 1 0 21160 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_230
timestamp 1604666999
transform 1 0 22264 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_242
timestamp 1604666999
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604666999
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604666999
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1472 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4692 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604666999
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_36
timestamp 1604666999
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_58
timestamp 1604666999
transform 1 0 6440 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7176 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_62
timestamp 1604666999
transform 1 0 6808 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_65
timestamp 1604666999
transform 1 0 7084 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1604666999
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1604666999
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_83
timestamp 1604666999
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_87
timestamp 1604666999
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_97
timestamp 1604666999
transform 1 0 10028 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10304 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1604666999
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12788 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_123
timestamp 1604666999
transform 1 0 12420 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1604666999
transform 1 0 13616 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604666999
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_140
timestamp 1604666999
transform 1 0 13984 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_143
timestamp 1604666999
transform 1 0 14260 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1604666999
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1604666999
transform 1 0 15548 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16376 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 15732 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_161
timestamp 1604666999
transform 1 0 15916 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_165
timestamp 1604666999
transform 1 0 16284 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_185
timestamp 1604666999
transform 1 0 18124 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1604666999
transform 1 0 19228 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1604666999
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1604666999
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604666999
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604666999
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604666999
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604666999
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1656 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_19
timestamp 1604666999
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 3220 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_32
timestamp 1604666999
transform 1 0 4048 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_37
timestamp 1604666999
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_41
timestamp 1604666999
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604666999
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604666999
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_72
timestamp 1604666999
transform 1 0 7728 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_77
timestamp 1604666999
transform 1 0 8188 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604666999
transform 1 0 8464 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 9476 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1604666999
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1604666999
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604666999
transform 1 0 11040 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604666999
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604666999
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1604666999
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1604666999
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1604666999
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1604666999
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_36.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13064 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_127
timestamp 1604666999
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14628 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1604666999
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1604666999
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_166
timestamp 1604666999
transform 1 0 16376 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1604666999
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1604666999
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19044 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_187
timestamp 1604666999
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_191
timestamp 1604666999
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_198
timestamp 1604666999
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604666999
transform 1 0 20424 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604666999
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_202
timestamp 1604666999
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1604666999
transform 1 0 20056 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_214
timestamp 1604666999
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_218
timestamp 1604666999
transform 1 0 21160 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_230
timestamp 1604666999
transform 1 0 22264 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_242
timestamp 1604666999
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604666999
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604666999
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604666999
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_6
timestamp 1604666999
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_19
timestamp 1604666999
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1604666999
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_10
timestamp 1604666999
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604666999
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1604666999
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1604666999
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604666999
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604666999
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_31
timestamp 1604666999
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_36
timestamp 1604666999
transform 1 0 4416 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4232 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 4692 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_47
timestamp 1604666999
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1604666999
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_48
timestamp 1604666999
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_55
timestamp 1604666999
transform 1 0 6164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_51
timestamp 1604666999
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_52
timestamp 1604666999
transform 1 0 5888 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_66
timestamp 1604666999
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1604666999
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1604666999
transform 1 0 7268 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_79
timestamp 1604666999
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_73
timestamp 1604666999
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7544 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1604666999
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_89
timestamp 1604666999
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_84
timestamp 1604666999
transform 1 0 8832 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1604666999
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9108 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1604666999
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1604666999
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1604666999
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604666999
transform 1 0 10764 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_114
timestamp 1604666999
transform 1 0 11592 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1604666999
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_117
timestamp 1604666999
transform 1 0 11868 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1604666999
transform 1 0 11500 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604666999
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1604666999
transform 1 0 11960 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_127
timestamp 1604666999
transform 1 0 12788 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1604666999
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp 1604666999
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12788 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1604666999
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_145
timestamp 1604666999
transform 1 0 14444 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_140
timestamp 1604666999
transform 1 0 13984 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604666999
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_150
timestamp 1604666999
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1604666999
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15272 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16652 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_161
timestamp 1604666999
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1604666999
transform 1 0 16284 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1604666999
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_177
timestamp 1604666999
transform 1 0 17388 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19136 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1604666999
transform 1 0 18400 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_187
timestamp 1604666999
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_191
timestamp 1604666999
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_199
timestamp 1604666999
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1604666999
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_203
timestamp 1604666999
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_215
timestamp 1604666999
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604666999
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_227
timestamp 1604666999
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604666999
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604666999
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1604666999
transform 1 0 23092 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_243
timestamp 1604666999
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604666999
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604666999
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604666999
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2300 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1604666999
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1604666999
transform 1 0 3496 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_22
timestamp 1604666999
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604666999
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_36
timestamp 1604666999
transform 1 0 4416 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604666999
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604666999
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4692 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1604666999
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7636 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_64
timestamp 1604666999
transform 1 0 6992 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_68
timestamp 1604666999
transform 1 0 7360 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_84
timestamp 1604666999
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_80
timestamp 1604666999
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604666999
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_88
timestamp 1604666999
transform 1 0 9200 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1604666999
transform 1 0 10028 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10580 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13064 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_122
timestamp 1604666999
transform 1 0 12328 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_126
timestamp 1604666999
transform 1 0 12696 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_129
timestamp 1604666999
transform 1 0 12972 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_36.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_139
timestamp 1604666999
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_143
timestamp 1604666999
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1604666999
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16836 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_163
timestamp 1604666999
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_174
timestamp 1604666999
transform 1 0 17112 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 17848 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_185
timestamp 1604666999
transform 1 0 18124 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1604666999
transform 1 0 19228 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1604666999
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1604666999
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604666999
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604666999
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604666999
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604666999
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2208 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1604666999
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1604666999
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1604666999
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_48
timestamp 1604666999
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_52
timestamp 1604666999
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_56
timestamp 1604666999
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9292 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_81
timestamp 1604666999
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_85
timestamp 1604666999
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 1604666999
transform 1 0 10120 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604666999
transform 1 0 10856 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_104
timestamp 1604666999
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1604666999
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13524 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_126
timestamp 1604666999
transform 1 0 12696 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1604666999
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_154
timestamp 1604666999
transform 1 0 15272 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604666999
transform 1 0 16284 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604666999
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_162
timestamp 1604666999
transform 1 0 16008 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1604666999
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1604666999
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1604666999
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604666999
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604666999
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604666999
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_248
timestamp 1604666999
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_252
timestamp 1604666999
transform 1 0 24288 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_264
timestamp 1604666999
transform 1 0 25392 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604666999
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 1748 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_16
timestamp 1604666999
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_20
timestamp 1604666999
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_24
timestamp 1604666999
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_28
timestamp 1604666999
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604666999
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5152 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1604666999
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7636 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_63
timestamp 1604666999
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604666999
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604666999
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_97
timestamp 1604666999
transform 1 0 10028 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10488 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1604666999
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1604666999
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1604666999
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_142
timestamp 1604666999
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1604666999
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_157
timestamp 1604666999
transform 1 0 15548 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1604666999
transform 1 0 16284 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1604666999
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1604666999
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_192
timestamp 1604666999
transform 1 0 18768 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1604666999
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604666999
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604666999
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604666999
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604666999
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604666999
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1564 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_14
timestamp 1604666999
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 1604666999
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 3128 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_31
timestamp 1604666999
transform 1 0 3956 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1604666999
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4784 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1604666999
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604666999
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604666999
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7452 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_66
timestamp 1604666999
transform 1 0 7176 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_78
timestamp 1604666999
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1604666999
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_105
timestamp 1604666999
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1604666999
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1604666999
transform 1 0 11500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604666999
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14904 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_142
timestamp 1604666999
transform 1 0 14168 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_153
timestamp 1604666999
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1604666999
transform 1 0 15548 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604666999
transform 1 0 15916 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_164
timestamp 1604666999
transform 1 0 16192 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_176
timestamp 1604666999
transform 1 0 17296 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1604666999
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604666999
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604666999
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604666999
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604666999
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604666999
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604666999
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1472 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604666999
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_38
timestamp 1604666999
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 4968 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_51
timestamp 1604666999
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_55
timestamp 1604666999
transform 1 0 6164 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_59
timestamp 1604666999
transform 1 0 6532 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6624 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_32_79
timestamp 1604666999
transform 1 0 8372 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_87
timestamp 1604666999
transform 1 0 9108 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_96
timestamp 1604666999
transform 1 0 9936 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10764 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_102
timestamp 1604666999
transform 1 0 10488 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1604666999
transform 1 0 11592 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_118
timestamp 1604666999
transform 1 0 11960 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12328 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12144 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1604666999
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_145
timestamp 1604666999
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_157
timestamp 1604666999
transform 1 0 15548 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_169
timestamp 1604666999
transform 1 0 16652 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_181
timestamp 1604666999
transform 1 0 17756 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_193
timestamp 1604666999
transform 1 0 18860 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_205
timestamp 1604666999
transform 1 0 19964 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604666999
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604666999
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604666999
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604666999
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604666999
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_7
timestamp 1604666999
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604666999
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 1932 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604666999
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_19
timestamp 1604666999
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_11
timestamp 1604666999
transform 1 0 2116 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 2300 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604666999
transform 1 0 2484 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 1932 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604666999
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_28
timestamp 1604666999
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604666999
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_32
timestamp 1604666999
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 4416 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1604666999
transform 1 0 5612 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_45
timestamp 1604666999
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_55
timestamp 1604666999
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_51
timestamp 1604666999
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604666999
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6348 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6532 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7820 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp 1604666999
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1604666999
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_78
timestamp 1604666999
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_86
timestamp 1604666999
transform 1 0 9016 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1604666999
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_92
timestamp 1604666999
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1604666999
transform 1 0 9936 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_96
timestamp 1604666999
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_106
timestamp 1604666999
transform 1 0 10856 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_102
timestamp 1604666999
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_109
timestamp 1604666999
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10304 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10304 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604666999
transform 1 0 11132 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1604666999
transform 1 0 11960 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604666999
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1604666999
transform 1 0 11500 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1604666999
transform 1 0 12604 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_122
timestamp 1604666999
transform 1 0 12328 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1604666999
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604666999
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12696 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13984 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_149
timestamp 1604666999
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_153
timestamp 1604666999
transform 1 0 15180 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_145
timestamp 1604666999
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_165
timestamp 1604666999
transform 1 0 16284 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1604666999
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604666999
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604666999
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604666999
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604666999
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604666999
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604666999
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604666999
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604666999
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604666999
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604666999
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604666999
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604666999
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604666999
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1604666999
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_11
timestamp 1604666999
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_19
timestamp 1604666999
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 3220 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3036 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_32
timestamp 1604666999
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_36
timestamp 1604666999
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_40
timestamp 1604666999
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_53
timestamp 1604666999
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1604666999
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_71
timestamp 1604666999
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1604666999
transform 1 0 8004 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8556 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604666999
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_100
timestamp 1604666999
transform 1 0 10304 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1604666999
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_110
timestamp 1604666999
transform 1 0 11224 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604666999
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13156 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12972 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12604 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_127
timestamp 1604666999
transform 1 0 12788 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_150
timestamp 1604666999
transform 1 0 14904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_162
timestamp 1604666999
transform 1 0 16008 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_174
timestamp 1604666999
transform 1 0 17112 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1604666999
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604666999
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604666999
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604666999
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604666999
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604666999
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604666999
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604666999
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604666999
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1748 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_16
timestamp 1604666999
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_20
timestamp 1604666999
transform 1 0 2944 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_25
timestamp 1604666999
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1604666999
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_36
timestamp 1604666999
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4968 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6532 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5980 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6348 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_40
timestamp 1604666999
transform 1 0 4784 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_51
timestamp 1604666999
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_55
timestamp 1604666999
transform 1 0 6164 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 8096 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7544 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 7912 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_68
timestamp 1604666999
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1604666999
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_79
timestamp 1604666999
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_83
timestamp 1604666999
transform 1 0 8740 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1604666999
transform 1 0 9292 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_96
timestamp 1604666999
transform 1 0 9936 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10672 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10396 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_100
timestamp 1604666999
transform 1 0 10304 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_103
timestamp 1604666999
transform 1 0 10580 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_113
timestamp 1604666999
transform 1 0 11500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12512 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13524 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_121
timestamp 1604666999
transform 1 0 12236 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_133
timestamp 1604666999
transform 1 0 13340 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_137
timestamp 1604666999
transform 1 0 13708 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1604666999
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604666999
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604666999
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604666999
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604666999
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604666999
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604666999
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604666999
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604666999
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604666999
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604666999
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604666999
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2208 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604666999
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1604666999
transform 1 0 2116 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_31
timestamp 1604666999
transform 1 0 3956 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_36
timestamp 1604666999
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_40
timestamp 1604666999
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604666999
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604666999
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 7636 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 7452 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_62
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_67
timestamp 1604666999
transform 1 0 7268 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_90
timestamp 1604666999
transform 1 0 9384 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1604666999
transform 1 0 9844 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10396 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1604666999
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604666999
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604666999
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13524 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_126
timestamp 1604666999
transform 1 0 12696 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_131
timestamp 1604666999
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604666999
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_154
timestamp 1604666999
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_158
timestamp 1604666999
transform 1 0 15640 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16100 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604666999
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_162
timestamp 1604666999
transform 1 0 16008 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1604666999
transform 1 0 16376 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_170
timestamp 1604666999
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_174
timestamp 1604666999
transform 1 0 17112 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1604666999
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1604666999
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_188
timestamp 1604666999
transform 1 0 18400 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_192
timestamp 1604666999
transform 1 0 18768 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_195
timestamp 1604666999
transform 1 0 19044 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_207
timestamp 1604666999
transform 1 0 20148 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_217
timestamp 1604666999
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604666999
transform 1 0 22172 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_231
timestamp 1604666999
transform 1 0 22356 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23276 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_239
timestamp 1604666999
transform 1 0 23092 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1604666999
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604666999
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604666999
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604666999
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 1932 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 1748 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_18
timestamp 1604666999
transform 1 0 2760 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4600 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1604666999
transform 1 0 3128 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_28
timestamp 1604666999
transform 1 0 3680 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_57
timestamp 1604666999
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7084 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_61
timestamp 1604666999
transform 1 0 6716 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_84
timestamp 1604666999
transform 1 0 8832 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11776 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_102
timestamp 1604666999
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_106
timestamp 1604666999
transform 1 0 10856 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_114
timestamp 1604666999
transform 1 0 11592 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13708 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_135
timestamp 1604666999
transform 1 0 13524 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604666999
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_139
timestamp 1604666999
transform 1 0 13892 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_151
timestamp 1604666999
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_158
timestamp 1604666999
transform 1 0 15640 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604666999
transform 1 0 16560 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_166
timestamp 1604666999
transform 1 0 16376 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_172
timestamp 1604666999
transform 1 0 16928 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 17848 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18860 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_180
timestamp 1604666999
transform 1 0 17664 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1604666999
transform 1 0 18124 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_196
timestamp 1604666999
transform 1 0 19136 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_208
timestamp 1604666999
transform 1 0 20240 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_218
timestamp 1604666999
transform 1 0 21160 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604666999
transform 1 0 22172 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_226
timestamp 1604666999
transform 1 0 21896 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_233
timestamp 1604666999
transform 1 0 22540 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23276 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_244
timestamp 1604666999
transform 1 0 23552 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_256
timestamp 1604666999
transform 1 0 24656 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604666999
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_268
timestamp 1604666999
transform 1 0 25760 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604666999
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604666999
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604666999
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604666999
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2116 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2116 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_40_28
timestamp 1604666999
transform 1 0 3680 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1604666999
transform 1 0 3312 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_20
timestamp 1604666999
transform 1 0 2944 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_36
timestamp 1604666999
transform 1 0 4416 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_37
timestamp 1604666999
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_34
timestamp 1604666999
transform 1 0 4232 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_30
timestamp 1604666999
transform 1 0 3864 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4232 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4692 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4876 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5888 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_50
timestamp 1604666999
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_54
timestamp 1604666999
transform 1 0 6072 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_58
timestamp 1604666999
transform 1 0 6440 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_58
timestamp 1604666999
transform 1 0 6440 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_65
timestamp 1604666999
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_62
timestamp 1604666999
transform 1 0 6808 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_62
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6900 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7084 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7452 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_39_78
timestamp 1604666999
transform 1 0 8280 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_74
timestamp 1604666999
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_78
timestamp 1604666999
transform 1 0 8280 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_86
timestamp 1604666999
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604666999
transform 1 0 8740 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_90
timestamp 1604666999
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9752 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11316 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12052 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1604666999
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_117
timestamp 1604666999
transform 1 0 11868 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_102
timestamp 1604666999
transform 1 0 10488 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_110
timestamp 1604666999
transform 1 0 11224 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604666999
transform 1 0 12696 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13708 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1604666999
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_123
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_129
timestamp 1604666999
transform 1 0 12972 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_130
timestamp 1604666999
transform 1 0 13064 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604666999
transform 1 0 15456 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604666999
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604666999
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_156
timestamp 1604666999
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_142
timestamp 1604666999
transform 1 0 14168 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_150
timestamp 1604666999
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1604666999
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_168
timestamp 1604666999
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_160
timestamp 1604666999
transform 1 0 15824 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604666999
transform 1 0 16192 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_172
timestamp 1604666999
transform 1 0 16928 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_176
timestamp 1604666999
transform 1 0 17296 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_172
timestamp 1604666999
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604666999
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604666999
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604666999
transform 1 0 17112 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604666999
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_160
timestamp 1604666999
transform 1 0 15824 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604666999
transform 1 0 18400 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604666999
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604666999
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_182
timestamp 1604666999
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_184
timestamp 1604666999
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1604666999
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_196
timestamp 1604666999
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604666999
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_208
timestamp 1604666999
transform 1 0 20240 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1604666999
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604666999
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604666999
transform 1 0 19504 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_215
timestamp 1604666999
transform 1 0 20884 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_216
timestamp 1604666999
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604666999
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604666999
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604666999
transform 1 0 20608 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604666999
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_227
timestamp 1604666999
transform 1 0 21988 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_220
timestamp 1604666999
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604666999
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604666999
transform 1 0 21712 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604666999
transform 1 0 21620 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_232
timestamp 1604666999
transform 1 0 22448 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_228
timestamp 1604666999
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604666999
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604666999
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604666999
transform 1 0 22724 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_237
timestamp 1604666999
transform 1 0 22908 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_239
timestamp 1604666999
transform 1 0 23092 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1604666999
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604666999
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604666999
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604666999
transform 1 0 23828 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1604666999
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_249
timestamp 1604666999
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604666999
transform 1 0 24564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604666999
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604666999
transform 1 0 24748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1604666999
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604666999
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604666999
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_261
timestamp 1604666999
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1604666999
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604666999
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604666999
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 2392 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604666999
transform 1 0 1840 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604666999
transform 1 0 2208 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_6
timestamp 1604666999
transform 1 0 1656 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_10
timestamp 1604666999
transform 1 0 2024 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 3956 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1604666999
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_27
timestamp 1604666999
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604666999
transform 1 0 5520 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604666999
transform 1 0 6072 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5336 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_40
timestamp 1604666999
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_44
timestamp 1604666999
transform 1 0 5152 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_52
timestamp 1604666999
transform 1 0 5888 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_56
timestamp 1604666999
transform 1 0 6256 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7728 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_60
timestamp 1604666999
transform 1 0 6624 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_68
timestamp 1604666999
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9660 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_81
timestamp 1604666999
transform 1 0 8556 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_89
timestamp 1604666999
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_112
timestamp 1604666999
transform 1 0 11408 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604666999
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_132
timestamp 1604666999
transform 1 0 13248 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_144
timestamp 1604666999
transform 1 0 14352 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_156
timestamp 1604666999
transform 1 0 15456 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_168
timestamp 1604666999
transform 1 0 16560 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604666999
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1604666999
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604666999
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604666999
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604666999
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604666999
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604666999
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604666999
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604666999
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604666999
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604666999
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604666999
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 2300 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1932 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_7
timestamp 1604666999
transform 1 0 1748 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_11
timestamp 1604666999
transform 1 0 2116 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_19
timestamp 1604666999
transform 1 0 2852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4232 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 3036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_23
timestamp 1604666999
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_32
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604666999
transform 1 0 5796 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_43
timestamp 1604666999
transform 1 0 5060 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_54
timestamp 1604666999
transform 1 0 6072 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604666999
transform 1 0 7912 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1604666999
transform 1 0 6900 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_66
timestamp 1604666999
transform 1 0 7176 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_77
timestamp 1604666999
transform 1 0 8188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1604666999
transform 1 0 9292 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604666999
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604666999
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604666999
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604666999
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_125
timestamp 1604666999
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_129
timestamp 1604666999
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604666999
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1604666999
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_153
timestamp 1604666999
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604666999
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604666999
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604666999
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604666999
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604666999
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604666999
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604666999
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604666999
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604666999
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604666999
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604666999
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604666999
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604666999
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604666999
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604666999
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 13910 0 13966 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 23202 0 23258 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21904 480 22024 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 82 nsew default input
rlabel metal3 s 0 23672 480 23792 6 left_top_grid_pin_42_
port 83 nsew default input
rlabel metal3 s 0 24216 480 24336 6 left_top_grid_pin_43_
port 84 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 85 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 86 nsew default input
rlabel metal3 s 0 25984 480 26104 6 left_top_grid_pin_46_
port 87 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 88 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 89 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 90 nsew default input
rlabel metal2 s 4618 0 4674 480 6 prog_clk
port 91 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 92 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 93 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 94 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_37_
port 95 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_38_
port 96 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 97 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_40_
port 98 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_41_
port 99 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 100 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 101 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 102 nsew default input
<< properties >>
string FIXED_BBOX 0 0 27679 28000
<< end >>
