* NGSPICE file created from cbx_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

.subckt cbx_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_14_ top_grid_pin_2_ top_grid_pin_6_ vpwr vgnd
XFILLER_22_133 vpwr vgnd scs8hd_fill_2
XFILLER_22_144 vgnd vpwr scs8hd_decap_6
XFILLER_26_52 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_148 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__113__B _111_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_129 vgnd vpwr scs8hd_decap_4
XFILLER_10_125 vpwr vgnd scs8hd_fill_2
XFILLER_10_169 vgnd vpwr scs8hd_decap_4
XFILLER_12_21 vpwr vgnd scs8hd_fill_2
XFILLER_12_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__108__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vpwr vgnd scs8hd_fill_2
XFILLER_5_151 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_3_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA__124__A _052_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _041_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_062_ address[4] _122_/B _076_/C _068_/B vgnd vpwr scs8hd_or3_4
X_131_ _131_/HI _131_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_2_143 vgnd vpwr scs8hd_decap_4
XFILLER_2_121 vpwr vgnd scs8hd_fill_2
XFILLER_2_110 vpwr vgnd scs8hd_fill_2
XFILLER_0_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _056_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_20 vpwr vgnd scs8hd_fill_2
XFILLER_18_42 vpwr vgnd scs8hd_fill_2
XFILLER_18_86 vgnd vpwr scs8hd_decap_6
X_045_ address[6] _049_/B vgnd vpwr scs8hd_inv_8
Xmem_top_ipin_5.LATCH_0_.latch data_in mem_top_ipin_5.LATCH_0_.latch/Q _090_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__105__C address[5] vgnd vpwr scs8hd_diode_2
X_114_ _121_/A _111_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _136_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_117 vgnd vpwr scs8hd_decap_4
XFILLER_29_106 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_10 vpwr vgnd scs8hd_fill_2
XFILLER_20_54 vpwr vgnd scs8hd_fill_2
XFILLER_29_30 vpwr vgnd scs8hd_fill_2
XFILLER_28_150 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_7.LATCH_3_.latch data_in mem_top_ipin_7.LATCH_3_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__116__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _129_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB _053_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__042__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_54 vpwr vgnd scs8hd_fill_2
XFILLER_15_76 vpwr vgnd scs8hd_fill_2
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_156 vgnd vpwr scs8hd_decap_12
XFILLER_31_112 vgnd vpwr scs8hd_decap_12
XFILLER_31_101 vgnd vpwr scs8hd_decap_4
XANTENNA__127__A _058_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_75 vpwr vgnd scs8hd_fill_2
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_4
XFILLER_13_167 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_193 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__C _122_/C vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _122_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__140__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA__050__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _130_/HI _130_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_10 vpwr vgnd scs8hd_fill_2
X_061_ _051_/B _121_/A _061_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_87 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_9_12 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_56 vgnd vpwr scs8hd_decap_3
XANTENNA__045__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_fill_1
XFILLER_18_65 vpwr vgnd scs8hd_fill_2
X_113_ _058_/X _111_/B _113_/Y vgnd vpwr scs8hd_nor2_4
X_044_ enable _098_/C vgnd vpwr scs8hd_inv_8
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_140 vgnd vpwr scs8hd_decap_3
XFILLER_19_173 vpwr vgnd scs8hd_fill_2
XFILLER_25_198 vpwr vgnd scs8hd_fill_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_3.LATCH_3_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_15_99 vpwr vgnd scs8hd_fill_2
XFILLER_31_168 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _122_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XANTENNA__143__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__053__A _051_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _124_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_87 vgnd vpwr scs8hd_decap_3
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_25 vpwr vgnd scs8hd_fill_2
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XFILLER_12_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__048__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_10_105 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_ipin_7.LATCH_4_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__050__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_4
XFILLER_3_3 vgnd vpwr scs8hd_decap_3
X_060_ address[1] address[2] address[0] _121_/A vgnd vpwr scs8hd_or3_4
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XANTENNA__151__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__061__A _051_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_043_ address[2] _052_/B vgnd vpwr scs8hd_inv_8
XFILLER_7_204 vpwr vgnd scs8hd_fill_2
XFILLER_11_200 vgnd vpwr scs8hd_fill_1
X_112_ _056_/X _111_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _137_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__056__A _054_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB _077_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_4
XFILLER_29_87 vgnd vpwr scs8hd_decap_6
XFILLER_29_43 vpwr vgnd scs8hd_fill_2
XFILLER_6_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_0_.latch data_in mem_top_ipin_1.LATCH_0_.latch/Q _061_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_152 vpwr vgnd scs8hd_fill_2
XFILLER_25_111 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_122 vpwr vgnd scs8hd_fill_2
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_ipin_3.LATCH_3_.latch data_in mem_top_ipin_3.LATCH_3_.latch/Q _072_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_103 vgnd vpwr scs8hd_decap_4
XANTENNA__053__B _052_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_90 vgnd vpwr scs8hd_decap_3
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_21_191 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__048__B _052_/B vgnd vpwr scs8hd_diode_2
XANTENNA__064__A _052_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_13 vpwr vgnd scs8hd_fill_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_4
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_0_.latch data_in _041_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__050__C _076_/C vgnd vpwr scs8hd_diode_2
XANTENNA__059__A _051_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XFILLER_2_168 vgnd vpwr scs8hd_decap_3
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_3_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA__061__B _121_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_78 vpwr vgnd scs8hd_fill_2
X_042_ address[1] _054_/A vgnd vpwr scs8hd_inv_8
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_111_ _054_/X _111_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_81 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__056__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _054_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_35 vgnd vpwr scs8hd_decap_4
XFILLER_29_99 vgnd vpwr scs8hd_decap_4
XFILLER_29_66 vpwr vgnd scs8hd_fill_2
XFILLER_29_55 vgnd vpwr scs8hd_decap_4
XFILLER_28_142 vgnd vpwr scs8hd_decap_8
XFILLER_28_131 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__157__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_197 vpwr vgnd scs8hd_fill_2
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XFILLER_25_178 vpwr vgnd scs8hd_fill_2
XFILLER_25_167 vpwr vgnd scs8hd_fill_2
XFILLER_25_156 vgnd vpwr scs8hd_decap_4
XFILLER_25_134 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A _058_/X vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_6.LATCH_2_.latch data_in mem_top_ipin_6.LATCH_2_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_13 vpwr vgnd scs8hd_fill_2
XFILLER_31_56 vgnd vpwr scs8hd_decap_4
XFILLER_31_45 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_4_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_0_200 vgnd vpwr scs8hd_decap_12
XFILLER_16_189 vpwr vgnd scs8hd_fill_2
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _040_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_137 vpwr vgnd scs8hd_fill_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_13_148 vpwr vgnd scs8hd_fill_2
XFILLER_3_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB _075_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__048__C _054_/C vgnd vpwr scs8hd_diode_2
XANTENNA__064__B _068_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_118 vgnd vpwr scs8hd_decap_4
XFILLER_10_129 vpwr vgnd scs8hd_fill_2
XFILLER_12_25 vgnd vpwr scs8hd_decap_4
XANTENNA__080__A _056_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_177 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__059__B _058_/X vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_68 vpwr vgnd scs8hd_fill_2
XFILLER_2_125 vgnd vpwr scs8hd_decap_4
XFILLER_0_39 vpwr vgnd scs8hd_fill_2
XFILLER_9_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_24 vpwr vgnd scs8hd_fill_2
XFILLER_18_46 vpwr vgnd scs8hd_fill_2
X_110_ _052_/X _111_/B _110_/Y vgnd vpwr scs8hd_nor2_4
X_041_ _041_/A _041_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _129_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _138_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__056__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_209 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _059_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__072__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_58 vpwr vgnd scs8hd_fill_2
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_6_49 vpwr vgnd scs8hd_fill_2
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _049_/B vgnd vpwr scs8hd_diode_2
XANTENNA__067__B _068_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_116 vgnd vpwr scs8hd_decap_6
XFILLER_26_79 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__078__A _052_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_1.LATCH_3_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_8_131 vpwr vgnd scs8hd_fill_2
XFILLER_8_142 vpwr vgnd scs8hd_fill_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__080__B _079_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_5_156 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XFILLER_4_71 vpwr vgnd scs8hd_fill_2
XANTENNA__075__B _074_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_211 vgnd vpwr scs8hd_fill_1
XFILLER_9_16 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_4_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA__086__A _052_/X vgnd vpwr scs8hd_diode_2
X_040_ _040_/A _040_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_177 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__083__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_16_103 vgnd vpwr scs8hd_decap_8
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_139 vpwr vgnd scs8hd_fill_2
XFILLER_31_128 vpwr vgnd scs8hd_fill_2
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_158 vgnd vpwr scs8hd_decap_4
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__078__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_36 vgnd vpwr scs8hd_fill_1
XANTENNA__094__A _054_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_2_.latch data_in mem_top_ipin_2.LATCH_2_.latch/Q _066_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_194 vgnd vpwr scs8hd_decap_4
XFILLER_8_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__089__A _058_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_209 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_4.LATCH_5_.latch data_in mem_top_ipin_4.LATCH_5_.latch/Q _077_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_168 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__091__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_81 vgnd vpwr scs8hd_fill_1
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
XANTENNA__086__B _088_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_204 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_24_80 vgnd vpwr scs8hd_fill_1
X_099_ _051_/A _101_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _139_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_29_47 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_18 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_10_60 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XFILLER_19_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_115 vgnd vpwr scs8hd_fill_1
XFILLER_15_49 vgnd vpwr scs8hd_decap_3
XFILLER_16_126 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_140 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_5.LATCH_1_.latch data_in mem_top_ipin_5.LATCH_1_.latch/Q _089_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_48 vpwr vgnd scs8hd_fill_2
XANTENNA__094__B _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_129 vpwr vgnd scs8hd_fill_2
XFILLER_8_111 vgnd vpwr scs8hd_decap_3
XFILLER_8_166 vgnd vpwr scs8hd_fill_1
XFILLER_12_140 vgnd vpwr scs8hd_fill_1
XFILLER_12_173 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_4_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_4_.latch data_in mem_top_ipin_7.LATCH_4_.latch/Q _100_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB _065_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_17 vpwr vgnd scs8hd_fill_2
XANTENNA__089__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_210 vpwr vgnd scs8hd_fill_2
XFILLER_5_103 vpwr vgnd scs8hd_fill_2
XFILLER_5_136 vpwr vgnd scs8hd_fill_2
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_4_180 vgnd vpwr scs8hd_decap_4
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XFILLER_23_202 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_6
XFILLER_3_8 vpwr vgnd scs8hd_fill_2
XFILLER_2_106 vpwr vgnd scs8hd_fill_2
XANTENNA__091__C _098_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_93 vpwr vgnd scs8hd_fill_2
XFILLER_29_7 vgnd vpwr scs8hd_decap_3
XFILLER_1_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_098_ _122_/A address[3] _098_/C _098_/D _101_/B vgnd vpwr scs8hd_or4_4
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_26 vpwr vgnd scs8hd_fill_2
XFILLER_28_168 vgnd vpwr scs8hd_decap_12
XFILLER_28_157 vgnd vpwr scs8hd_decap_8
XFILLER_28_113 vgnd vpwr scs8hd_decap_12
XFILLER_28_102 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XANTENNA__097__B _091_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_92 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_138 vgnd vpwr scs8hd_decap_3
XFILLER_15_17 vpwr vgnd scs8hd_fill_2
XFILLER_31_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_108 vpwr vgnd scs8hd_fill_2
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_193 vpwr vgnd scs8hd_fill_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XFILLER_21_82 vpwr vgnd scs8hd_fill_2
XFILLER_11_7 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vgnd vpwr scs8hd_decap_4
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_7_95 vgnd vpwr scs8hd_decap_3
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_71 vgnd vpwr scs8hd_decap_3
XFILLER_16_93 vgnd vpwr scs8hd_fill_1
XFILLER_8_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_129 vgnd vpwr scs8hd_fill_1
XANTENNA__091__D _098_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_097_ _121_/A _091_/X _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_97 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _131_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
XFILLER_29_16 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_3.LATCH_4_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_136 vpwr vgnd scs8hd_fill_2
XFILLER_19_169 vpwr vgnd scs8hd_fill_2
X_149_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_180 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_139 vgnd vpwr scs8hd_decap_12
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_172 vgnd vpwr scs8hd_decap_4
XFILLER_7_41 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _139_/HI mem_top_ipin_7.LATCH_5_.latch/Q
+ mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_12_120 vgnd vpwr scs8hd_fill_1
XFILLER_16_83 vgnd vpwr scs8hd_decap_6
XFILLER_8_146 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_12_ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_1.LATCH_1_.latch data_in mem_top_ipin_1.LATCH_1_.latch/Q _059_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_82 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_42 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_3.LATCH_4_.latch data_in mem_top_ipin_3.LATCH_4_.latch/Q _071_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_73 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _052_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_83 vgnd vpwr scs8hd_decap_6
X_096_ _058_/X _091_/X _096_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_21 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_1.LATCH_1_.latch data_in _040_/A _106_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XFILLER_10_85 vgnd vpwr scs8hd_decap_6
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_148_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
X_079_ _054_/X _079_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_25_107 vpwr vgnd scs8hd_fill_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XFILLER_21_154 vpwr vgnd scs8hd_fill_2
XFILLER_21_187 vpwr vgnd scs8hd_fill_2
XFILLER_21_198 vpwr vgnd scs8hd_fill_2
XFILLER_12_132 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XFILLER_8_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_0_.latch data_in mem_top_ipin_4.LATCH_0_.latch/Q _082_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__103__A _058_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_202 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_94 vpwr vgnd scs8hd_fill_2
XFILLER_27_50 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_6.LATCH_3_.latch data_in mem_top_ipin_6.LATCH_3_.latch/Q _094_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_54 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_fill_1
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_4_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_1_131 vpwr vgnd scs8hd_fill_2
XANTENNA__100__B _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_197 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_095_ _056_/X _091_/X _095_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _054_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_77 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _138_/HI mem_top_ipin_6.LATCH_5_.latch/Q
+ mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_204 vpwr vgnd scs8hd_fill_2
XFILLER_10_64 vpwr vgnd scs8hd_fill_2
XFILLER_19_95 vpwr vgnd scs8hd_fill_2
XFILLER_19_116 vgnd vpwr scs8hd_decap_4
X_147_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
X_078_ _052_/X _079_/B _078_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_31_19 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_185 vgnd vpwr scs8hd_decap_8
XFILLER_24_174 vgnd vpwr scs8hd_decap_8
XFILLER_24_163 vgnd vpwr scs8hd_decap_8
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_41 vgnd vpwr scs8hd_decap_3
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_26_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _068_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vpwr vgnd scs8hd_fill_2
XFILLER_12_177 vpwr vgnd scs8hd_fill_2
XFILLER_16_63 vpwr vgnd scs8hd_fill_2
XANTENNA__103__B _101_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XFILLER_4_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_206 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_97 vgnd vpwr scs8hd_decap_4
XFILLER_1_154 vpwr vgnd scs8hd_fill_2
XFILLER_1_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _051_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_209 vgnd vpwr scs8hd_decap_3
XFILLER_24_63 vpwr vgnd scs8hd_fill_2
XFILLER_24_41 vgnd vpwr scs8hd_decap_3
XFILLER_24_30 vgnd vpwr scs8hd_fill_1
X_094_ _054_/X _091_/X _094_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_106 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_30 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _122_/B vgnd vpwr scs8hd_diode_2
X_146_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
X_077_ _051_/A _079_/B _077_/Y vgnd vpwr scs8hd_nor2_4
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
XFILLER_21_86 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_1.LATCH_4_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XANTENNA__117__A _052_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_129_ _129_/HI _129_/LO vgnd vpwr scs8hd_conb_1
XFILLER_21_123 vgnd vpwr scs8hd_fill_1
XFILLER_8_127 vpwr vgnd scs8hd_fill_2
XFILLER_12_112 vgnd vpwr scs8hd_decap_8
XFILLER_12_145 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_17_204 vpwr vgnd scs8hd_fill_2
XFILLER_27_74 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_67 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _137_/HI mem_top_ipin_5.LATCH_5_.latch/Q
+ mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _128_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__040__A _040_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_177 vgnd vpwr scs8hd_decap_4
XANTENNA__109__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _054_/X vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_3_.latch data_in mem_top_ipin_2.LATCH_3_.latch/Q _065_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_093_ _052_/X _091_/X _093_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_13 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_22 vpwr vgnd scs8hd_fill_2
XFILLER_10_77 vpwr vgnd scs8hd_fill_2
XFILLER_10_99 vgnd vpwr scs8hd_decap_4
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_173 vpwr vgnd scs8hd_fill_2
XFILLER_27_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_145_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__106__C _122_/C vgnd vpwr scs8hd_diode_2
XANTENNA__122__B _122_/B vgnd vpwr scs8hd_diode_2
X_076_ _122_/A _122_/B _076_/C _079_/B vgnd vpwr scs8hd_or3_4
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_132 vpwr vgnd scs8hd_fill_2
XFILLER_24_121 vgnd vpwr scs8hd_decap_4
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XFILLER_15_176 vgnd vpwr scs8hd_fill_1
XANTENNA__117__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
X_128_ _121_/A _122_/X _128_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_059_ _051_/B _058_/X _059_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_113 vgnd vpwr scs8hd_decap_3
XFILLER_21_135 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vgnd vpwr scs8hd_decap_4
XANTENNA__043__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_142 vgnd vpwr scs8hd_decap_4
XFILLER_4_197 vgnd vpwr scs8hd_decap_12
XFILLER_4_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_22 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_5.LATCH_2_.latch data_in mem_top_ipin_5.LATCH_2_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_44 vpwr vgnd scs8hd_fill_2
XFILLER_13_77 vgnd vpwr scs8hd_decap_4
XFILLER_1_167 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA__141__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__051__A _051_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_5_.latch data_in mem_top_ipin_7.LATCH_5_.latch/Q _099_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_24_76 vgnd vpwr scs8hd_decap_4
XFILLER_10_211 vgnd vpwr scs8hd_fill_1
X_092_ _051_/A _091_/X _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__046__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_45 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_27_141 vgnd vpwr scs8hd_decap_3
X_075_ _121_/A _074_/B _075_/Y vgnd vpwr scs8hd_nor2_4
X_144_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__106__D _054_/C vgnd vpwr scs8hd_diode_2
XANTENNA__122__C _122_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_22 vgnd vpwr scs8hd_decap_3
XPHY_8 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _136_/HI mem_top_ipin_4.LATCH_5_.latch/Q
+ mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_155 vpwr vgnd scs8hd_fill_2
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
X_058_ address[1] address[2] _054_/C _058_/X vgnd vpwr scs8hd_or3_4
X_127_ _058_/X _122_/X _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_24 vpwr vgnd scs8hd_fill_2
XFILLER_7_46 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_79 vpwr vgnd scs8hd_fill_2
XFILLER_21_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB _055_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vpwr vgnd scs8hd_fill_2
XFILLER_12_136 vgnd vpwr scs8hd_decap_4
XFILLER_12_158 vgnd vpwr scs8hd_decap_6
XFILLER_20_180 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__144__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_173 vgnd vpwr scs8hd_decap_4
XANTENNA__054__A _054_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_98 vpwr vgnd scs8hd_fill_2
XFILLER_27_54 vgnd vpwr scs8hd_fill_1
XFILLER_4_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__049__A enable vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_135 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__051__B _051_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_22 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_091_ address[4] _122_/B _098_/C _098_/D _091_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__152__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_109 vgnd vpwr scs8hd_fill_1
XFILLER_3_208 vgnd vpwr scs8hd_decap_4
XANTENNA__062__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_19_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_074_ _058_/X _074_/B _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_186 vpwr vgnd scs8hd_fill_2
XFILLER_18_197 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
XANTENNA__057__A _051_/B vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_057_ _051_/B _056_/X _057_/Y vgnd vpwr scs8hd_nor2_4
X_126_ _056_/X _122_/X _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_6 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_45 vgnd vpwr scs8hd_decap_4
XFILLER_16_67 vpwr vgnd scs8hd_fill_2
XFILLER_16_89 vgnd vpwr scs8hd_fill_1
XFILLER_7_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_109_ _051_/A _111_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__054__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_11 vpwr vgnd scs8hd_fill_2
XANTENNA__070__A _051_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__155__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__049__B _049_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_210 vpwr vgnd scs8hd_fill_2
XANTENNA__065__A _054_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _135_/HI mem_top_ipin_3.LATCH_5_.latch/Q
+ mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_24_89 vgnd vpwr scs8hd_fill_1
X_090_ _121_/A _088_/B _090_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_ipin_1.LATCH_2_.latch data_in mem_top_ipin_1.LATCH_2_.latch/Q _057_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__062__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_14 vpwr vgnd scs8hd_fill_2
XFILLER_10_36 vgnd vpwr scs8hd_decap_3
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_34 vpwr vgnd scs8hd_fill_2
X_142_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_3.LATCH_5_.latch data_in mem_top_ipin_3.LATCH_5_.latch/Q _070_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_073_ _056_/X _074_/B _073_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__057__B _056_/X vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__073__A _056_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_125_ _054_/X _122_/X _125_/Y vgnd vpwr scs8hd_nor2_4
X_056_ _054_/A address[2] address[0] _056_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_105 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_197 vgnd vpwr scs8hd_decap_4
XFILLER_11_193 vgnd vpwr scs8hd_decap_4
X_108_ address[4] address[3] _122_/C _111_/B vgnd vpwr scs8hd_or3_4
X_039_ address[0] _054_/C vgnd vpwr scs8hd_inv_8
XANTENNA__054__C _054_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
XANTENNA__070__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_34 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_208 vgnd vpwr scs8hd_decap_4
XFILLER_27_78 vgnd vpwr scs8hd_decap_4
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XFILLER_31_211 vgnd vpwr scs8hd_fill_1
XANTENNA__049__C address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__065__B _068_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_14 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A _058_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB _063_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_1_.latch data_in mem_top_ipin_4.LATCH_1_.latch/Q _081_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__076__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_46 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_6.LATCH_4_.latch data_in mem_top_ipin_6.LATCH_4_.latch/Q _093_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__062__C _076_/C vgnd vpwr scs8hd_diode_2
XFILLER_10_26 vpwr vgnd scs8hd_fill_2
XFILLER_19_13 vpwr vgnd scs8hd_fill_2
XFILLER_27_177 vgnd vpwr scs8hd_decap_6
XFILLER_27_111 vpwr vgnd scs8hd_fill_2
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_141_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
X_072_ _054_/X _074_/B _072_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_111 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_125 vgnd vpwr scs8hd_fill_1
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_14 vpwr vgnd scs8hd_fill_2
XANTENNA__073__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_36 vgnd vpwr scs8hd_decap_3
XFILLER_15_103 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
X_055_ _051_/B _054_/X _055_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_16 vpwr vgnd scs8hd_fill_2
X_124_ _052_/X _122_/X _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_191 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_139 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__068__B _068_/B vgnd vpwr scs8hd_diode_2
XANTENNA__084__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
X_107_ address[4] _122_/B _122_/C address[0] _107_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _134_/HI mem_top_ipin_2.LATCH_5_.latch/Q
+ mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_81 vgnd vpwr scs8hd_decap_4
XANTENNA__079__A _054_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_46 vpwr vgnd scs8hd_fill_2
XFILLER_27_24 vpwr vgnd scs8hd_fill_2
XFILLER_4_146 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_26 vgnd vpwr scs8hd_fill_1
XFILLER_13_48 vpwr vgnd scs8hd_fill_2
XANTENNA__081__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_7.LATCH_0_.latch data_in mem_top_ipin_7.LATCH_0_.latch/Q _104_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XANTENNA__076__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_36 vgnd vpwr scs8hd_decap_3
XFILLER_24_14 vpwr vgnd scs8hd_fill_2
XANTENNA__092__A _051_/A vgnd vpwr scs8hd_diode_2
XANTENNA__087__A _054_/X vgnd vpwr scs8hd_diode_2
X_071_ _052_/X _074_/B _071_/Y vgnd vpwr scs8hd_nor2_4
X_140_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XFILLER_18_167 vgnd vpwr scs8hd_decap_4
XFILLER_25_90 vgnd vpwr scs8hd_decap_3
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_8
XFILLER_30_118 vgnd vpwr scs8hd_decap_8
XFILLER_30_107 vgnd vpwr scs8hd_decap_8
XFILLER_15_159 vpwr vgnd scs8hd_fill_2
X_054_ _054_/A address[2] _054_/C _054_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_28 vpwr vgnd scs8hd_fill_2
X_123_ _051_/A _122_/X _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _061_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_92 vgnd vpwr scs8hd_decap_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__084__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_111 vgnd vpwr scs8hd_decap_3
XFILLER_11_162 vpwr vgnd scs8hd_fill_2
X_106_ address[4] _122_/B _122_/C _054_/C _106_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__079__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_210 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _056_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_202 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_1_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__076__C _076_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_59 vpwr vgnd scs8hd_fill_2
XFILLER_24_26 vgnd vpwr scs8hd_decap_4
XANTENNA__092__B _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_209 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_26 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _088_/B vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ _051_/A _074_/B _070_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _133_/HI mem_top_ipin_1.LATCH_5_.latch/Q
+ mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_124 vpwr vgnd scs8hd_fill_2
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_2.LATCH_4_.latch data_in mem_top_ipin_2.LATCH_4_.latch/Q _064_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__098__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_149 vgnd vpwr scs8hd_decap_4
X_122_ _122_/A _122_/B _122_/C _122_/X vgnd vpwr scs8hd_or3_4
X_053_ _051_/B _052_/X _053_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
XFILLER_14_182 vpwr vgnd scs8hd_fill_2
XANTENNA__084__C _098_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_49 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_156 vpwr vgnd scs8hd_fill_2
X_105_ _098_/C address[6] address[5] _122_/C vgnd vpwr scs8hd_or3_4
XFILLER_22_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__095__B _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_91 vgnd vpwr scs8hd_fill_1
XFILLER_0_173 vgnd vpwr scs8hd_fill_1
XFILLER_5_40 vpwr vgnd scs8hd_fill_2
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_3.LATCH_0_.latch data_in mem_top_ipin_3.LATCH_0_.latch/Q _075_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_18 vpwr vgnd scs8hd_fill_2
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_27_147 vgnd vpwr scs8hd_decap_8
XFILLER_27_136 vgnd vpwr scs8hd_decap_3
XFILLER_19_38 vgnd vpwr scs8hd_decap_4
XFILLER_27_169 vpwr vgnd scs8hd_fill_2
XFILLER_18_114 vgnd vpwr scs8hd_fill_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_ipin_5.LATCH_3_.latch data_in mem_top_ipin_5.LATCH_3_.latch/Q _087_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_63 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XFILLER_24_128 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__098__B address[3] vgnd vpwr scs8hd_diode_2
X_121_ _121_/A _121_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_150 vpwr vgnd scs8hd_fill_2
X_052_ address[1] _052_/B address[0] _052_/X vgnd vpwr scs8hd_or3_4
XFILLER_14_150 vgnd vpwr scs8hd_decap_3
XFILLER_21_109 vpwr vgnd scs8hd_fill_2
XFILLER_29_209 vgnd vpwr scs8hd_decap_3
XANTENNA__084__D _098_/D vgnd vpwr scs8hd_diode_2
XFILLER_20_142 vgnd vpwr scs8hd_fill_1
XFILLER_20_197 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vgnd vpwr scs8hd_fill_1
X_104_ _121_/A _101_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_93 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XFILLER_4_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_201 vgnd vpwr scs8hd_decap_8
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_18 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _132_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB _066_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_208 vgnd vpwr scs8hd_decap_4
XFILLER_13_204 vpwr vgnd scs8hd_fill_2
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XFILLER_0_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_18 vpwr vgnd scs8hd_fill_2
XANTENNA__098__C _098_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_107 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_051_ _051_/A _051_/B _051_/Y vgnd vpwr scs8hd_nor2_4
X_120_ _058_/X _121_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_121 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
X_103_ _058_/X _101_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_136 vgnd vpwr scs8hd_decap_3
XFILLER_7_169 vpwr vgnd scs8hd_fill_2
XFILLER_22_50 vpwr vgnd scs8hd_fill_2
XFILLER_8_41 vgnd vpwr scs8hd_decap_4
XFILLER_6_180 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_28 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_202 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _040_/A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_75 vgnd vpwr scs8hd_decap_3
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_24_18 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _054_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_43 vpwr vgnd scs8hd_fill_2
XFILLER_2_10 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_108 vpwr vgnd scs8hd_fill_2
XFILLER_17_160 vpwr vgnd scs8hd_fill_2
XFILLER_17_171 vpwr vgnd scs8hd_fill_2
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__D _098_/D vgnd vpwr scs8hd_diode_2
XFILLER_23_130 vgnd vpwr scs8hd_decap_3
XFILLER_23_163 vpwr vgnd scs8hd_fill_2
XFILLER_23_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_050_ address[4] address[3] _076_/C _051_/B vgnd vpwr scs8hd_or3_4
XFILLER_11_30 vpwr vgnd scs8hd_fill_2
XFILLER_11_96 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_3_.latch data_in mem_top_ipin_1.LATCH_3_.latch/Q _055_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_155 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
X_102_ _056_/X _101_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_62 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_40 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_162 vpwr vgnd scs8hd_fill_2
XFILLER_3_140 vgnd vpwr scs8hd_decap_4
XANTENNA__104__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_121 vgnd vpwr scs8hd_decap_3
XFILLER_28_83 vgnd vpwr scs8hd_decap_8
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XFILLER_30_62 vgnd vpwr scs8hd_fill_1
XANTENNA__101__B _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_128 vgnd vpwr scs8hd_decap_4
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_95 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA__112__A _056_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_4.LATCH_2_.latch data_in mem_top_ipin_4.LATCH_2_.latch/Q _080_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_142 vgnd vpwr scs8hd_decap_8
XFILLER_14_186 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XFILLER_20_167 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_6.LATCH_5_.latch data_in mem_top_ipin_6.LATCH_5_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_101_ _054_/X _101_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_116 vgnd vpwr scs8hd_decap_4
XFILLER_22_85 vgnd vpwr scs8hd_decap_6
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_87 vpwr vgnd scs8hd_fill_2
XFILLER_4_108 vpwr vgnd scs8hd_fill_2
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XANTENNA__104__B _101_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _058_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB _051_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_44 vgnd vpwr scs8hd_decap_4
XANTENNA__115__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_53 vpwr vgnd scs8hd_fill_2
XFILLER_30_41 vgnd vpwr scs8hd_decap_8
XFILLER_14_64 vpwr vgnd scs8hd_fill_2
XFILLER_14_75 vpwr vgnd scs8hd_fill_2
XFILLER_30_96 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_107 vgnd vpwr scs8hd_decap_4
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_41 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XANTENNA__112__B _111_/B vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_1_.latch data_in mem_top_ipin_7.LATCH_1_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XFILLER_23_198 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_21 vgnd vpwr scs8hd_decap_3
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
XFILLER_14_165 vpwr vgnd scs8hd_fill_2
XANTENNA__107__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _051_/A vgnd vpwr scs8hd_diode_2
X_100_ _052_/X _101_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _054_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_77 vpwr vgnd scs8hd_fill_2
XFILLER_17_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vgnd vpwr scs8hd_decap_4
XFILLER_3_197 vgnd vpwr scs8hd_decap_4
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_208 vgnd vpwr scs8hd_decap_4
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_89 vgnd vpwr scs8hd_decap_4
XFILLER_5_23 vgnd vpwr scs8hd_decap_4
XANTENNA__115__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__041__A _041_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_87 vgnd vpwr scs8hd_decap_3
XFILLER_30_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_204 vpwr vgnd scs8hd_fill_2
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _056_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_119 vgnd vpwr scs8hd_fill_1
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vgnd vpwr scs8hd_decap_6
XFILLER_25_20 vpwr vgnd scs8hd_fill_2
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_6 vpwr vgnd scs8hd_fill_2
XFILLER_11_44 vgnd vpwr scs8hd_decap_3
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
XFILLER_11_99 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_199 vgnd vpwr scs8hd_decap_12
XANTENNA__107__C _122_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_158 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_4
XFILLER_22_54 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _126_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_23 vgnd vpwr scs8hd_decap_6
XFILLER_8_45 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__118__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA__044__A enable vgnd vpwr scs8hd_diode_2
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_2.LATCH_5_.latch data_in mem_top_ipin_2.LATCH_5_.latch/Q _063_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__039__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_113 vpwr vgnd scs8hd_fill_2
XFILLER_28_64 vgnd vpwr scs8hd_fill_1
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA__115__C _122_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_22 vpwr vgnd scs8hd_fill_2
XFILLER_30_65 vgnd vpwr scs8hd_fill_1
XFILLER_30_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _122_/X vgnd vpwr scs8hd_diode_2
XANTENNA__142__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__052__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_54 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_2_47 vgnd vpwr scs8hd_decap_3
XFILLER_17_164 vpwr vgnd scs8hd_fill_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_197 vgnd vpwr scs8hd_decap_4
XANTENNA__047__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_167 vpwr vgnd scs8hd_fill_2
XFILLER_23_178 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_34 vgnd vpwr scs8hd_fill_1
XANTENNA__107__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_28_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XFILLER_20_104 vpwr vgnd scs8hd_fill_2
XFILLER_20_126 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_3.LATCH_1_.latch data_in mem_top_ipin_3.LATCH_1_.latch/Q _074_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _041_/A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XFILLER_22_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_204 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_089_ _058_/X _088_/B _089_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_163 vgnd vpwr scs8hd_decap_4
XFILLER_26_3 vgnd vpwr scs8hd_decap_4
XANTENNA__150__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_5.LATCH_4_.latch data_in mem_top_ipin_5.LATCH_4_.latch/Q _086_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__060__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_44 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_144 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_210 vpwr vgnd scs8hd_fill_2
XANTENNA__145__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__055__A _051_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_43 vpwr vgnd scs8hd_fill_2
XFILLER_28_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_169 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_14_45 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__052__B _052_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_209 vgnd vpwr scs8hd_decap_3
XFILLER_26_121 vpwr vgnd scs8hd_fill_2
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XFILLER_25_33 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_143 vpwr vgnd scs8hd_fill_2
XANTENNA__153__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_146 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A _051_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_6.LATCH_0_.latch data_in mem_top_ipin_6.LATCH_0_.latch/Q _097_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__148__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_138 vgnd vpwr scs8hd_decap_4
XFILLER_20_149 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_149 vgnd vpwr scs8hd_decap_6
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
XFILLER_10_182 vpwr vgnd scs8hd_fill_2
X_157_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_186 vpwr vgnd scs8hd_fill_2
XFILLER_6_197 vgnd vpwr scs8hd_decap_12
X_088_ _056_/X _088_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__060__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB _057_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_70 vpwr vgnd scs8hd_fill_2
XANTENNA__055__B _054_/X vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _052_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_148 vgnd vpwr scs8hd_decap_4
XFILLER_5_15 vpwr vgnd scs8hd_fill_2
XFILLER_8_204 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__156__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__066__A _056_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_23 vgnd vpwr scs8hd_decap_8
XFILLER_14_79 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_163 vgnd vpwr scs8hd_decap_12
XFILLER_29_152 vgnd vpwr scs8hd_decap_4
XFILLER_29_141 vpwr vgnd scs8hd_fill_2
XFILLER_29_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__052__C address[0] vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_31_180 vgnd vpwr scs8hd_decap_6
XANTENNA__063__B _068_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
XFILLER_14_169 vpwr vgnd scs8hd_fill_2
XFILLER_22_180 vgnd vpwr scs8hd_decap_8
XFILLER_22_191 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_3_92 vgnd vpwr scs8hd_decap_3
XANTENNA__058__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _058_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
X_156_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_087_ _054_/X _088_/B _087_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_48 vgnd vpwr scs8hd_fill_1
XANTENNA__069__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA__060__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_209 vgnd vpwr scs8hd_decap_3
XFILLER_17_24 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _130_/HI _040_/Y mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
X_139_ _139_/HI _139_/LO vgnd vpwr scs8hd_conb_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_4
XANTENNA__071__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_67 vgnd vpwr scs8hd_decap_3
XFILLER_28_56 vgnd vpwr scs8hd_decap_8
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_1.LATCH_4_.latch data_in mem_top_ipin_1.LATCH_4_.latch/Q _053_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _132_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__066__B _068_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_14 vpwr vgnd scs8hd_fill_2
XFILLER_14_58 vgnd vpwr scs8hd_decap_4
XFILLER_30_79 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vgnd vpwr scs8hd_decap_4
XANTENNA__082__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_197 vgnd vpwr scs8hd_decap_12
XFILLER_29_175 vgnd vpwr scs8hd_decap_8
XFILLER_20_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_70 vgnd vpwr scs8hd_decap_3
XFILLER_26_145 vgnd vpwr scs8hd_decap_8
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _051_/A vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _130_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_126 vpwr vgnd scs8hd_fill_2
XFILLER_11_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__058__C _054_/C vgnd vpwr scs8hd_diode_2
XANTENNA__074__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_22_36 vgnd vpwr scs8hd_fill_1
XFILLER_22_58 vgnd vpwr scs8hd_fill_1
XANTENNA__090__A _121_/A vgnd vpwr scs8hd_diode_2
X_155_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_086_ _052_/X _088_/B _086_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_ipin_2.LATCH_0_.latch data_in mem_top_ipin_2.LATCH_0_.latch/Q _068_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__069__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__085__A _051_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_158 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vpwr vgnd scs8hd_fill_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_138_ _138_/HI _138_/LO vgnd vpwr scs8hd_conb_1
X_069_ _122_/A address[3] _076_/C _074_/B vgnd vpwr scs8hd_or3_4
Xmem_top_ipin_4.LATCH_3_.latch data_in mem_top_ipin_4.LATCH_3_.latch/Q _079_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_180 vgnd vpwr scs8hd_decap_4
XFILLER_0_94 vpwr vgnd scs8hd_fill_2
XFILLER_21_202 vpwr vgnd scs8hd_fill_2
XFILLER_9_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_117 vpwr vgnd scs8hd_fill_2
XFILLER_28_79 vpwr vgnd scs8hd_fill_2
XFILLER_28_35 vpwr vgnd scs8hd_fill_2
XFILLER_12_202 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_26 vpwr vgnd scs8hd_fill_2
XFILLER_30_58 vgnd vpwr scs8hd_decap_4
XANTENNA__082__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XFILLER_29_110 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_179 vgnd vpwr scs8hd_decap_8
XFILLER_26_168 vgnd vpwr scs8hd_decap_8
XFILLER_26_157 vgnd vpwr scs8hd_decap_8
XFILLER_26_135 vgnd vpwr scs8hd_decap_8
XFILLER_26_113 vgnd vpwr scs8hd_decap_8
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _079_/B vgnd vpwr scs8hd_diode_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _052_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_80 vpwr vgnd scs8hd_fill_2
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _041_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_49 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _056_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_116 vgnd vpwr scs8hd_decap_3
XFILLER_14_138 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_20_108 vgnd vpwr scs8hd_decap_4
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XANTENNA__090__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_208 vgnd vpwr scs8hd_decap_4
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
X_085_ _051_/A _088_/B _085_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_112 vpwr vgnd scs8hd_fill_2
X_154_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_81 vgnd vpwr scs8hd_decap_3
XFILLER_26_7 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_211 vgnd vpwr scs8hd_fill_1
XANTENNA__069__C _076_/C vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_2_.latch data_in mem_top_ipin_7.LATCH_2_.latch/Q _102_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__085__B _088_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_137_ _137_/HI _137_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
X_068_ _121_/A _068_/B _068_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_129 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _058_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _133_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_49 vpwr vgnd scs8hd_fill_2
XFILLER_29_188 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_125 vgnd vpwr scs8hd_fill_1
XFILLER_25_37 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _091_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_103 vpwr vgnd scs8hd_fill_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_191 vpwr vgnd scs8hd_fill_2
XFILLER_31_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
XANTENNA__088__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_150 vgnd vpwr scs8hd_fill_1
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_9_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_73 vpwr vgnd scs8hd_fill_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A _051_/A vgnd vpwr scs8hd_diode_2
X_153_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_135 vgnd vpwr scs8hd_decap_6
XFILLER_10_142 vpwr vgnd scs8hd_fill_2
XFILLER_10_186 vpwr vgnd scs8hd_fill_2
X_084_ address[4] address[3] _098_/C _098_/D _088_/B vgnd vpwr scs8hd_or4_4
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_7 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_136_ _136_/HI _136_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_81 vgnd vpwr scs8hd_decap_4
X_067_ _058_/X _068_/B _067_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_ipin_7.LATCH_3_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_119_ _056_/X _121_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _125_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_71 vgnd vpwr scs8hd_decap_8
XFILLER_20_82 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_31_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_23_118 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_100 vgnd vpwr scs8hd_decap_3
XFILLER_9_144 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__099__B _101_/B vgnd vpwr scs8hd_diode_2
X_152_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_083_ _049_/B address[5] _098_/D vgnd vpwr scs8hd_or2_4
XFILLER_10_165 vpwr vgnd scs8hd_fill_2
XFILLER_6_169 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_28 vgnd vpwr scs8hd_decap_3
XFILLER_3_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_135_ _135_/HI _135_/LO vgnd vpwr scs8hd_conb_1
X_066_ _056_/X _068_/B _066_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_7 vgnd vpwr scs8hd_fill_1
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_3.LATCH_2_.latch data_in mem_top_ipin_3.LATCH_2_.latch/Q _073_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_82 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _134_/HI vgnd vpwr
+ scs8hd_diode_2
X_049_ enable _049_/B address[5] _076_/C vgnd vpwr scs8hd_nand3_4
X_118_ _054_/X _121_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XFILLER_14_18 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_5.LATCH_5_.latch data_in mem_top_ipin_5.LATCH_5_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_204 vpwr vgnd scs8hd_fill_2
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_193 vgnd vpwr scs8hd_decap_4
XFILLER_23_108 vgnd vpwr scs8hd_decap_4
XFILLER_14_108 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _041_/Y mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_163 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_3_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_26_60 vpwr vgnd scs8hd_fill_2
XFILLER_13_163 vpwr vgnd scs8hd_fill_2
XFILLER_3_97 vgnd vpwr scs8hd_decap_3
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_151_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
Xmux_top_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_122 vgnd vpwr scs8hd_fill_1
XFILLER_10_199 vgnd vpwr scs8hd_decap_12
X_082_ _121_/A _079_/B _082_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
X_065_ _054_/X _068_/B _065_/Y vgnd vpwr scs8hd_nor2_4
X_134_ _134_/HI _134_/LO vgnd vpwr scs8hd_conb_1
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
XFILLER_21_206 vgnd vpwr scs8hd_decap_6
Xmem_top_ipin_6.LATCH_1_.latch data_in mem_top_ipin_6.LATCH_1_.latch/Q _096_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_52 vpwr vgnd scs8hd_fill_2
XFILLER_9_96 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _040_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _131_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_61 vpwr vgnd scs8hd_fill_2
X_117_ _052_/X _121_/B _117_/Y vgnd vpwr scs8hd_nor2_4
X_048_ address[1] _052_/B _054_/C _051_/A vgnd vpwr scs8hd_or3_4
XFILLER_15_3 vgnd vpwr scs8hd_fill_1
XFILLER_29_114 vgnd vpwr scs8hd_fill_1
XFILLER_29_103 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_93 vgnd vpwr scs8hd_fill_1
XFILLER_28_180 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _067_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_64 vgnd vpwr scs8hd_decap_4
XFILLER_6_97 vpwr vgnd scs8hd_fill_2
XFILLER_26_106 vgnd vpwr scs8hd_decap_4
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XFILLER_15_84 vgnd vpwr scs8hd_decap_4
XFILLER_17_128 vpwr vgnd scs8hd_fill_2
XFILLER_31_72 vgnd vpwr scs8hd_decap_8
XANTENNA__102__A _056_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_142 vgnd vpwr scs8hd_decap_4
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_21 vpwr vgnd scs8hd_fill_2
XFILLER_22_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_150_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_116 vgnd vpwr scs8hd_decap_4
X_081_ _058_/X _079_/B _081_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_204 vpwr vgnd scs8hd_fill_2
X_133_ _133_/HI _133_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XFILLER_2_163 vgnd vpwr scs8hd_decap_3
X_064_ _052_/X _068_/B _064_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__110__A _052_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_66 vpwr vgnd scs8hd_fill_2
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_14_ vgnd vpwr scs8hd_inv_1
X_116_ _051_/A _121_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _098_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_047_ address[3] _122_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _135_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_3_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_29_159 vpwr vgnd scs8hd_fill_2
XFILLER_29_148 vpwr vgnd scs8hd_fill_2
XFILLER_29_137 vpwr vgnd scs8hd_fill_2
XFILLER_29_126 vpwr vgnd scs8hd_fill_2
XFILLER_20_41 vpwr vgnd scs8hd_fill_2
XFILLER_29_83 vpwr vgnd scs8hd_fill_2
XFILLER_28_192 vgnd vpwr scs8hd_decap_12
XFILLER_6_43 vgnd vpwr scs8hd_decap_4
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_107 vpwr vgnd scs8hd_fill_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_84 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_1.LATCH_5_.latch data_in mem_top_ipin_1.LATCH_5_.latch/Q _051_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__102__B _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_162 vgnd vpwr scs8hd_fill_1
XFILLER_31_187 vgnd vpwr scs8hd_decap_12
XFILLER_31_143 vgnd vpwr scs8hd_decap_12
XFILLER_31_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_9_169 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__113__A _058_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_180 vgnd vpwr scs8hd_decap_4
XFILLER_10_146 vgnd vpwr scs8hd_decap_6
X_080_ _056_/X _079_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_3 vgnd vpwr scs8hd_decap_3
XFILLER_12_64 vpwr vgnd scs8hd_fill_2
XFILLER_12_86 vgnd vpwr scs8hd_decap_6
XFILLER_12_97 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
X_063_ _051_/A _068_/B _063_/Y vgnd vpwr scs8hd_nor2_4
X_132_ _132_/HI _132_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_197 vgnd vpwr scs8hd_decap_12
XFILLER_2_186 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_23 vgnd vpwr scs8hd_decap_4
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__105__B address[6] vgnd vpwr scs8hd_diode_2
X_115_ _122_/A address[3] _122_/C _121_/B vgnd vpwr scs8hd_or3_4
X_046_ address[4] _122_/A vgnd vpwr scs8hd_inv_8
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_2.LATCH_1_.latch data_in mem_top_ipin_2.LATCH_1_.latch/Q _067_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_fill_1
XFILLER_29_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__116__A _051_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_22 vgnd vpwr scs8hd_decap_3
XFILLER_6_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_4.LATCH_4_.latch data_in mem_top_ipin_4.LATCH_4_.latch/Q _078_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_25_174 vpwr vgnd scs8hd_fill_2
XFILLER_25_163 vpwr vgnd scs8hd_fill_2
XFILLER_25_152 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_52 vpwr vgnd scs8hd_fill_2
XFILLER_31_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_199 vgnd vpwr scs8hd_decap_12
.ends

