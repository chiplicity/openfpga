magic
tech EFS8A
magscale 1 2
timestamp 1604430969
<< locali >>
rect 26249 17051 26283 17289
rect 7757 12631 7791 12733
rect 21741 12699 21775 12937
rect 21189 11543 21223 11781
<< viali >>
rect 24317 21097 24351 21131
rect 25329 21097 25363 21131
rect 24133 20961 24167 20995
rect 25145 20961 25179 20995
rect 15577 20757 15611 20791
rect 19257 20757 19291 20791
rect 25697 20757 25731 20791
rect 26065 20757 26099 20791
rect 1593 20553 1627 20587
rect 7113 20553 7147 20587
rect 9505 20553 9539 20587
rect 12633 20553 12667 20587
rect 14289 20553 14323 20587
rect 17141 20553 17175 20587
rect 18245 20553 18279 20587
rect 20913 20553 20947 20587
rect 24409 20553 24443 20587
rect 4997 20485 5031 20519
rect 15669 20417 15703 20451
rect 19717 20417 19751 20451
rect 25421 20417 25455 20451
rect 26157 20417 26191 20451
rect 1409 20349 1443 20383
rect 4813 20349 4847 20383
rect 5273 20349 5307 20383
rect 6929 20349 6963 20383
rect 9321 20349 9355 20383
rect 12449 20349 12483 20383
rect 12909 20349 12943 20383
rect 14105 20349 14139 20383
rect 15485 20349 15519 20383
rect 16957 20349 16991 20383
rect 18061 20349 18095 20383
rect 18521 20349 18555 20383
rect 20729 20349 20763 20383
rect 21189 20349 21223 20383
rect 24225 20349 24259 20383
rect 14565 20281 14599 20315
rect 15577 20281 15611 20315
rect 19073 20281 19107 20315
rect 25973 20281 26007 20315
rect 1961 20213 1995 20247
rect 7481 20213 7515 20247
rect 9873 20213 9907 20247
rect 14013 20213 14047 20247
rect 14933 20213 14967 20247
rect 15117 20213 15151 20247
rect 17509 20213 17543 20247
rect 19165 20213 19199 20247
rect 19533 20213 19567 20247
rect 19625 20213 19659 20247
rect 23489 20213 23523 20247
rect 24133 20213 24167 20247
rect 24961 20213 24995 20247
rect 25513 20213 25547 20247
rect 25881 20213 25915 20247
rect 15761 20009 15795 20043
rect 17785 20009 17819 20043
rect 24041 19941 24075 19975
rect 12357 19873 12391 19907
rect 15669 19873 15703 19907
rect 18153 19873 18187 19907
rect 25237 19873 25271 19907
rect 12449 19805 12483 19839
rect 12541 19805 12575 19839
rect 15853 19805 15887 19839
rect 18245 19805 18279 19839
rect 18429 19805 18463 19839
rect 25329 19805 25363 19839
rect 25513 19805 25547 19839
rect 26525 19805 26559 19839
rect 24409 19737 24443 19771
rect 24869 19737 24903 19771
rect 1685 19669 1719 19703
rect 8677 19669 8711 19703
rect 10885 19669 10919 19703
rect 11805 19669 11839 19703
rect 11989 19669 12023 19703
rect 13001 19669 13035 19703
rect 15025 19669 15059 19703
rect 15301 19669 15335 19703
rect 19165 19669 19199 19703
rect 24777 19669 24811 19703
rect 25881 19669 25915 19703
rect 14933 19465 14967 19499
rect 24593 19465 24627 19499
rect 26341 19465 26375 19499
rect 10701 19397 10735 19431
rect 8493 19329 8527 19363
rect 9137 19329 9171 19363
rect 11345 19329 11379 19363
rect 13001 19329 13035 19363
rect 15485 19329 15519 19363
rect 25053 19329 25087 19363
rect 25145 19329 25179 19363
rect 26985 19329 27019 19363
rect 2789 19261 2823 19295
rect 3617 19261 3651 19295
rect 11253 19261 11287 19295
rect 12817 19261 12851 19295
rect 14841 19261 14875 19295
rect 15301 19261 15335 19295
rect 17509 19261 17543 19295
rect 19073 19261 19107 19295
rect 21833 19261 21867 19295
rect 22293 19261 22327 19295
rect 24133 19261 24167 19295
rect 24961 19261 24995 19295
rect 25881 19261 25915 19295
rect 26709 19261 26743 19295
rect 1685 19193 1719 19227
rect 8125 19193 8159 19227
rect 8953 19193 8987 19227
rect 10333 19193 10367 19227
rect 11161 19193 11195 19227
rect 14473 19193 14507 19227
rect 17141 19193 17175 19227
rect 19318 19193 19352 19227
rect 1777 19125 1811 19159
rect 2237 19125 2271 19159
rect 2973 19125 3007 19159
rect 3249 19125 3283 19159
rect 8585 19125 8619 19159
rect 9045 19125 9079 19159
rect 10793 19125 10827 19159
rect 11989 19125 12023 19159
rect 12449 19125 12483 19159
rect 12909 19125 12943 19159
rect 13553 19125 13587 19159
rect 13921 19125 13955 19159
rect 15393 19125 15427 19159
rect 15945 19125 15979 19159
rect 17877 19125 17911 19159
rect 18521 19125 18555 19159
rect 18981 19125 19015 19159
rect 20453 19125 20487 19159
rect 22017 19125 22051 19159
rect 24409 19125 24443 19159
rect 26157 19125 26191 19159
rect 26801 19125 26835 19159
rect 27353 19125 27387 19159
rect 1593 18921 1627 18955
rect 8769 18921 8803 18955
rect 10333 18921 10367 18955
rect 11345 18921 11379 18955
rect 11805 18921 11839 18955
rect 15485 18921 15519 18955
rect 19809 18921 19843 18955
rect 22477 18921 22511 18955
rect 25329 18921 25363 18955
rect 26525 18921 26559 18955
rect 26985 18921 27019 18955
rect 12142 18853 12176 18887
rect 16773 18853 16807 18887
rect 23857 18853 23891 18887
rect 24216 18853 24250 18887
rect 1961 18785 1995 18819
rect 5273 18785 5307 18819
rect 5365 18785 5399 18819
rect 8585 18785 8619 18819
rect 10701 18785 10735 18819
rect 16681 18785 16715 18819
rect 17785 18785 17819 18819
rect 18144 18785 18178 18819
rect 22385 18785 22419 18819
rect 23949 18785 23983 18819
rect 26893 18785 26927 18819
rect 2053 18717 2087 18751
rect 2145 18717 2179 18751
rect 2605 18717 2639 18751
rect 5457 18717 5491 18751
rect 10241 18717 10275 18751
rect 10793 18717 10827 18751
rect 10977 18717 11011 18751
rect 11897 18717 11931 18751
rect 16957 18717 16991 18751
rect 17877 18717 17911 18751
rect 20913 18717 20947 18751
rect 22569 18717 22603 18751
rect 27169 18717 27203 18751
rect 22017 18649 22051 18683
rect 2973 18581 3007 18615
rect 3341 18581 3375 18615
rect 3709 18581 3743 18615
rect 4905 18581 4939 18615
rect 13277 18581 13311 18615
rect 15025 18581 15059 18615
rect 16313 18581 16347 18615
rect 19257 18581 19291 18615
rect 20269 18581 20303 18615
rect 21833 18581 21867 18615
rect 23489 18581 23523 18615
rect 3065 18377 3099 18411
rect 9965 18377 9999 18411
rect 10609 18377 10643 18411
rect 11897 18377 11931 18411
rect 16497 18377 16531 18411
rect 17785 18377 17819 18411
rect 18705 18377 18739 18411
rect 19809 18377 19843 18411
rect 21465 18377 21499 18411
rect 23121 18377 23155 18411
rect 26893 18377 26927 18411
rect 27813 18377 27847 18411
rect 1501 18309 1535 18343
rect 1961 18241 1995 18275
rect 2145 18241 2179 18275
rect 3617 18241 3651 18275
rect 4169 18241 4203 18275
rect 5549 18241 5583 18275
rect 11253 18241 11287 18275
rect 19165 18241 19199 18275
rect 19349 18241 19383 18275
rect 20821 18241 20855 18275
rect 22569 18241 22603 18275
rect 24501 18241 24535 18275
rect 1869 18173 1903 18207
rect 3433 18173 3467 18207
rect 4537 18173 4571 18207
rect 6009 18173 6043 18207
rect 8585 18173 8619 18207
rect 12449 18173 12483 18207
rect 15025 18173 15059 18207
rect 15117 18173 15151 18207
rect 20177 18173 20211 18207
rect 20637 18173 20671 18207
rect 22477 18173 22511 18207
rect 25513 18173 25547 18207
rect 5365 18105 5399 18139
rect 8830 18105 8864 18139
rect 12716 18105 12750 18139
rect 14657 18105 14691 18139
rect 15384 18105 15418 18139
rect 19073 18105 19107 18139
rect 20729 18105 20763 18139
rect 21833 18105 21867 18139
rect 23489 18105 23523 18139
rect 24409 18105 24443 18139
rect 25758 18105 25792 18139
rect 27445 18105 27479 18139
rect 2513 18037 2547 18071
rect 2881 18037 2915 18071
rect 3525 18037 3559 18071
rect 4813 18037 4847 18071
rect 4997 18037 5031 18071
rect 5457 18037 5491 18071
rect 6469 18037 6503 18071
rect 7665 18037 7699 18071
rect 8125 18037 8159 18071
rect 8493 18037 8527 18071
rect 11345 18037 11379 18071
rect 13829 18037 13863 18071
rect 17049 18037 17083 18071
rect 17417 18037 17451 18071
rect 18337 18037 18371 18071
rect 20269 18037 20303 18071
rect 22017 18037 22051 18071
rect 22385 18037 22419 18071
rect 23949 18037 23983 18071
rect 24317 18037 24351 18071
rect 24961 18037 24995 18071
rect 25329 18037 25363 18071
rect 28181 18037 28215 18071
rect 2881 17833 2915 17867
rect 4261 17833 4295 17867
rect 4905 17833 4939 17867
rect 9045 17833 9079 17867
rect 9505 17833 9539 17867
rect 11713 17833 11747 17867
rect 12081 17833 12115 17867
rect 13277 17833 13311 17867
rect 13645 17833 13679 17867
rect 14933 17833 14967 17867
rect 17785 17833 17819 17867
rect 18889 17833 18923 17867
rect 19993 17833 20027 17867
rect 20361 17833 20395 17867
rect 21097 17833 21131 17867
rect 22017 17833 22051 17867
rect 1768 17765 1802 17799
rect 3433 17765 3467 17799
rect 10701 17765 10735 17799
rect 11529 17765 11563 17799
rect 16650 17765 16684 17799
rect 18613 17765 18647 17799
rect 24777 17765 24811 17799
rect 25237 17765 25271 17799
rect 5253 17697 5287 17731
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 13737 17697 13771 17731
rect 19257 17697 19291 17731
rect 22376 17697 22410 17731
rect 25329 17697 25363 17731
rect 26893 17697 26927 17731
rect 26985 17697 27019 17731
rect 1501 17629 1535 17663
rect 4997 17629 5031 17663
rect 8493 17629 8527 17663
rect 8585 17629 8619 17663
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 12173 17629 12207 17663
rect 12357 17629 12391 17663
rect 13921 17629 13955 17663
rect 15301 17629 15335 17663
rect 16405 17629 16439 17663
rect 19349 17629 19383 17663
rect 19441 17629 19475 17663
rect 22109 17629 22143 17663
rect 25513 17629 25547 17663
rect 27169 17629 27203 17663
rect 3801 17561 3835 17595
rect 8033 17561 8067 17595
rect 11069 17561 11103 17595
rect 23489 17561 23523 17595
rect 26525 17561 26559 17595
rect 6377 17493 6411 17527
rect 6929 17493 6963 17527
rect 7941 17493 7975 17527
rect 9689 17493 9723 17527
rect 12817 17493 12851 17527
rect 13093 17493 13127 17527
rect 21557 17493 21591 17527
rect 24041 17493 24075 17527
rect 24869 17493 24903 17527
rect 25881 17493 25915 17527
rect 26341 17493 26375 17527
rect 2973 17289 3007 17323
rect 5457 17289 5491 17323
rect 7941 17289 7975 17323
rect 10517 17289 10551 17323
rect 13921 17289 13955 17323
rect 14749 17289 14783 17323
rect 17141 17289 17175 17323
rect 20453 17289 20487 17323
rect 21373 17289 21407 17323
rect 21833 17289 21867 17323
rect 25973 17289 26007 17323
rect 26249 17289 26283 17323
rect 26525 17289 26559 17323
rect 17877 17221 17911 17255
rect 22845 17221 22879 17255
rect 23857 17221 23891 17255
rect 1593 17153 1627 17187
rect 7021 17153 7055 17187
rect 10977 17153 11011 17187
rect 11069 17153 11103 17187
rect 13093 17153 13127 17187
rect 13553 17153 13587 17187
rect 14841 17153 14875 17187
rect 21741 17153 21775 17187
rect 22477 17153 22511 17187
rect 24041 17153 24075 17187
rect 1860 17085 1894 17119
rect 4077 17085 4111 17119
rect 4344 17085 4378 17119
rect 8033 17085 8067 17119
rect 10333 17085 10367 17119
rect 15108 17085 15142 17119
rect 18521 17085 18555 17119
rect 18788 17085 18822 17119
rect 27077 17153 27111 17187
rect 27905 17153 27939 17187
rect 26985 17085 27019 17119
rect 7481 17017 7515 17051
rect 8300 17017 8334 17051
rect 10885 17017 10919 17051
rect 12817 17017 12851 17051
rect 21005 17017 21039 17051
rect 22293 17017 22327 17051
rect 24286 17017 24320 17051
rect 26249 17017 26283 17051
rect 26893 17017 26927 17051
rect 28273 17017 28307 17051
rect 3525 16949 3559 16983
rect 3893 16949 3927 16983
rect 6009 16949 6043 16983
rect 6561 16949 6595 16983
rect 9413 16949 9447 16983
rect 9965 16949 9999 16983
rect 11805 16949 11839 16983
rect 12173 16949 12207 16983
rect 12449 16949 12483 16983
rect 12909 16949 12943 16983
rect 14289 16949 14323 16983
rect 16221 16949 16255 16983
rect 16865 16949 16899 16983
rect 18429 16949 18463 16983
rect 19901 16949 19935 16983
rect 22201 16949 22235 16983
rect 23489 16949 23523 16983
rect 25421 16949 25455 16983
rect 26433 16949 26467 16983
rect 27629 16949 27663 16983
rect 1685 16745 1719 16779
rect 4077 16745 4111 16779
rect 4445 16745 4479 16779
rect 5549 16745 5583 16779
rect 6469 16745 6503 16779
rect 6837 16745 6871 16779
rect 8033 16745 8067 16779
rect 8401 16745 8435 16779
rect 10425 16745 10459 16779
rect 12817 16745 12851 16779
rect 13093 16745 13127 16779
rect 14105 16745 14139 16779
rect 15301 16745 15335 16779
rect 17233 16745 17267 16779
rect 17325 16745 17359 16779
rect 17969 16745 18003 16779
rect 18521 16745 18555 16779
rect 19533 16745 19567 16779
rect 24133 16745 24167 16779
rect 24869 16745 24903 16779
rect 26157 16745 26191 16779
rect 26525 16745 26559 16779
rect 2053 16677 2087 16711
rect 7481 16677 7515 16711
rect 8493 16677 8527 16711
rect 10854 16677 10888 16711
rect 13553 16677 13587 16711
rect 15761 16677 15795 16711
rect 18981 16677 19015 16711
rect 21557 16677 21591 16711
rect 25237 16677 25271 16711
rect 27629 16677 27663 16711
rect 2145 16609 2179 16643
rect 2789 16609 2823 16643
rect 5273 16609 5307 16643
rect 5917 16609 5951 16643
rect 13461 16609 13495 16643
rect 15669 16609 15703 16643
rect 18889 16609 18923 16643
rect 21905 16609 21939 16643
rect 24777 16609 24811 16643
rect 26893 16609 26927 16643
rect 26985 16609 27019 16643
rect 2329 16541 2363 16575
rect 3433 16541 3467 16575
rect 3801 16541 3835 16575
rect 4537 16541 4571 16575
rect 4629 16541 4663 16575
rect 6929 16541 6963 16575
rect 7113 16541 7147 16575
rect 8585 16541 8619 16575
rect 9873 16541 9907 16575
rect 10609 16541 10643 16575
rect 13737 16541 13771 16575
rect 15853 16541 15887 16575
rect 17417 16541 17451 16575
rect 19073 16541 19107 16575
rect 21649 16541 21683 16575
rect 25329 16541 25363 16575
rect 25421 16541 25455 16575
rect 27077 16541 27111 16575
rect 3065 16473 3099 16507
rect 6377 16473 6411 16507
rect 11989 16473 12023 16507
rect 16865 16473 16899 16507
rect 7941 16405 7975 16439
rect 9045 16405 9079 16439
rect 15117 16405 15151 16439
rect 18429 16405 18463 16439
rect 21189 16405 21223 16439
rect 23029 16405 23063 16439
rect 23765 16405 23799 16439
rect 1593 16201 1627 16235
rect 3157 16201 3191 16235
rect 4537 16201 4571 16235
rect 5181 16201 5215 16235
rect 6837 16201 6871 16235
rect 8125 16201 8159 16235
rect 9873 16201 9907 16235
rect 11069 16201 11103 16235
rect 11529 16201 11563 16235
rect 16313 16201 16347 16235
rect 17233 16201 17267 16235
rect 18245 16201 18279 16235
rect 21833 16201 21867 16235
rect 25053 16201 25087 16235
rect 27537 16201 27571 16235
rect 14105 16133 14139 16167
rect 14657 16133 14691 16167
rect 16957 16133 16991 16167
rect 21005 16133 21039 16167
rect 25605 16133 25639 16167
rect 2237 16065 2271 16099
rect 2605 16065 2639 16099
rect 3709 16065 3743 16099
rect 5825 16065 5859 16099
rect 7389 16065 7423 16099
rect 10701 16065 10735 16099
rect 12725 16065 12759 16099
rect 15761 16065 15795 16099
rect 22385 16065 22419 16099
rect 2053 15997 2087 16031
rect 6193 15997 6227 16031
rect 7297 15997 7331 16031
rect 8493 15997 8527 16031
rect 12992 15997 13026 16031
rect 15669 15997 15703 16031
rect 18429 15997 18463 16031
rect 18685 15997 18719 16031
rect 22293 15997 22327 16031
rect 22845 15997 22879 16031
rect 23673 15997 23707 16031
rect 23929 15997 23963 16031
rect 26157 15997 26191 16031
rect 3617 15929 3651 15963
rect 5089 15929 5123 15963
rect 5549 15929 5583 15963
rect 8738 15929 8772 15963
rect 11897 15929 11931 15963
rect 15577 15929 15611 15963
rect 17877 15929 17911 15963
rect 23397 15929 23431 15963
rect 25973 15929 26007 15963
rect 26402 15929 26436 15963
rect 28089 15929 28123 15963
rect 1961 15861 1995 15895
rect 3065 15861 3099 15895
rect 3525 15861 3559 15895
rect 4261 15861 4295 15895
rect 5641 15861 5675 15895
rect 6561 15861 6595 15895
rect 7205 15861 7239 15895
rect 12173 15861 12207 15895
rect 15025 15861 15059 15895
rect 15209 15861 15243 15895
rect 19809 15861 19843 15895
rect 21373 15861 21407 15895
rect 21741 15861 21775 15895
rect 22201 15861 22235 15895
rect 1777 15657 1811 15691
rect 2789 15657 2823 15691
rect 3617 15657 3651 15691
rect 4261 15657 4295 15691
rect 6837 15657 6871 15691
rect 8033 15657 8067 15691
rect 13185 15657 13219 15691
rect 14657 15657 14691 15691
rect 15117 15657 15151 15691
rect 18429 15657 18463 15691
rect 21741 15657 21775 15691
rect 23305 15657 23339 15691
rect 24869 15657 24903 15691
rect 27629 15657 27663 15691
rect 5080 15589 5114 15623
rect 23857 15589 23891 15623
rect 24777 15589 24811 15623
rect 26985 15589 27019 15623
rect 2145 15521 2179 15555
rect 8401 15521 8435 15555
rect 8493 15521 8527 15555
rect 9413 15521 9447 15555
rect 10609 15521 10643 15555
rect 10701 15521 10735 15555
rect 12061 15521 12095 15555
rect 14105 15521 14139 15555
rect 15568 15521 15602 15555
rect 18797 15521 18831 15555
rect 21465 15521 21499 15555
rect 22192 15521 22226 15555
rect 25237 15521 25271 15555
rect 26893 15521 26927 15555
rect 2237 15453 2271 15487
rect 2421 15453 2455 15487
rect 4813 15453 4847 15487
rect 8585 15453 8619 15487
rect 10885 15453 10919 15487
rect 11805 15453 11839 15487
rect 15301 15453 15335 15487
rect 18889 15453 18923 15487
rect 18981 15453 19015 15487
rect 21925 15453 21959 15487
rect 25329 15453 25363 15487
rect 25513 15453 25547 15487
rect 27169 15453 27203 15487
rect 10241 15385 10275 15419
rect 1593 15317 1627 15351
rect 3157 15317 3191 15351
rect 4721 15317 4755 15351
rect 6193 15317 6227 15351
rect 7481 15317 7515 15351
rect 7849 15317 7883 15351
rect 9045 15317 9079 15351
rect 9873 15317 9907 15351
rect 13737 15317 13771 15351
rect 16681 15317 16715 15351
rect 17233 15317 17267 15351
rect 18337 15317 18371 15351
rect 24225 15317 24259 15351
rect 26249 15317 26283 15351
rect 26525 15317 26559 15351
rect 3157 15113 3191 15147
rect 6653 15113 6687 15147
rect 8033 15113 8067 15147
rect 11621 15113 11655 15147
rect 13185 15113 13219 15147
rect 18429 15113 18463 15147
rect 21741 15113 21775 15147
rect 25973 15113 26007 15147
rect 4077 15045 4111 15079
rect 11989 15045 12023 15079
rect 14473 15045 14507 15079
rect 22753 15045 22787 15079
rect 25697 15045 25731 15079
rect 4261 14977 4295 15011
rect 7573 14977 7607 15011
rect 8677 14977 8711 15011
rect 13829 14977 13863 15011
rect 14013 14977 14047 15011
rect 15485 14977 15519 15011
rect 18981 14977 19015 15011
rect 19073 14977 19107 15011
rect 22385 14977 22419 15011
rect 24133 14977 24167 15011
rect 24225 14977 24259 15011
rect 1777 14909 1811 14943
rect 9597 14909 9631 14943
rect 13737 14909 13771 14943
rect 21281 14909 21315 14943
rect 22109 14909 22143 14943
rect 24041 14909 24075 14943
rect 26157 14909 26191 14943
rect 2044 14841 2078 14875
rect 4528 14841 4562 14875
rect 7849 14841 7883 14875
rect 8493 14841 8527 14875
rect 9864 14841 9898 14875
rect 15301 14841 15335 14875
rect 16313 14841 16347 14875
rect 19340 14841 19374 14875
rect 21649 14841 21683 14875
rect 22201 14841 22235 14875
rect 24961 14841 24995 14875
rect 26402 14841 26436 14875
rect 1593 14773 1627 14807
rect 3709 14773 3743 14807
rect 5641 14773 5675 14807
rect 6193 14773 6227 14807
rect 6837 14773 6871 14807
rect 8401 14773 8435 14807
rect 9045 14773 9079 14807
rect 9413 14773 9447 14807
rect 10977 14773 11011 14807
rect 12909 14773 12943 14807
rect 13369 14773 13403 14807
rect 14841 14773 14875 14807
rect 14933 14773 14967 14807
rect 15393 14773 15427 14807
rect 16037 14773 16071 14807
rect 17877 14773 17911 14807
rect 20453 14773 20487 14807
rect 23489 14773 23523 14807
rect 23673 14773 23707 14807
rect 25237 14773 25271 14807
rect 27537 14773 27571 14807
rect 28089 14773 28123 14807
rect 2881 14569 2915 14603
rect 3525 14569 3559 14603
rect 4905 14569 4939 14603
rect 7297 14569 7331 14603
rect 8033 14569 8067 14603
rect 10425 14569 10459 14603
rect 11713 14569 11747 14603
rect 13185 14569 13219 14603
rect 15485 14569 15519 14603
rect 18337 14569 18371 14603
rect 20361 14569 20395 14603
rect 24041 14569 24075 14603
rect 25789 14569 25823 14603
rect 26525 14569 26559 14603
rect 5632 14501 5666 14535
rect 8493 14501 8527 14535
rect 16396 14501 16430 14535
rect 19717 14501 19751 14535
rect 24409 14501 24443 14535
rect 25513 14501 25547 14535
rect 1501 14433 1535 14467
rect 1768 14433 1802 14467
rect 4077 14433 4111 14467
rect 5365 14433 5399 14467
rect 8401 14433 8435 14467
rect 9505 14433 9539 14467
rect 10517 14433 10551 14467
rect 11161 14433 11195 14467
rect 12072 14433 12106 14467
rect 16129 14433 16163 14467
rect 19625 14433 19659 14467
rect 21813 14433 21847 14467
rect 26893 14433 26927 14467
rect 8677 14365 8711 14399
rect 10609 14365 10643 14399
rect 11805 14365 11839 14399
rect 19901 14365 19935 14399
rect 21557 14365 21591 14399
rect 24501 14365 24535 14399
rect 24593 14365 24627 14399
rect 26157 14365 26191 14399
rect 26985 14365 27019 14399
rect 27169 14365 27203 14399
rect 9045 14297 9079 14331
rect 10057 14297 10091 14331
rect 19165 14297 19199 14331
rect 3893 14229 3927 14263
rect 4261 14229 4295 14263
rect 5273 14229 5307 14263
rect 6745 14229 6779 14263
rect 7941 14229 7975 14263
rect 9873 14229 9907 14263
rect 13829 14229 13863 14263
rect 15117 14229 15151 14263
rect 17509 14229 17543 14263
rect 18705 14229 18739 14263
rect 19257 14229 19291 14263
rect 21373 14229 21407 14263
rect 22937 14229 22971 14263
rect 23857 14229 23891 14263
rect 25053 14229 25087 14263
rect 1869 14025 1903 14059
rect 3065 14025 3099 14059
rect 3617 14025 3651 14059
rect 4721 14025 4755 14059
rect 6561 14025 6595 14059
rect 9781 14025 9815 14059
rect 10425 14025 10459 14059
rect 11253 14025 11287 14059
rect 11897 14025 11931 14059
rect 14841 14025 14875 14059
rect 15025 14025 15059 14059
rect 16497 14025 16531 14059
rect 17785 14025 17819 14059
rect 18429 14025 18463 14059
rect 18613 14025 18647 14059
rect 19625 14025 19659 14059
rect 20177 14025 20211 14059
rect 21557 14025 21591 14059
rect 21741 14025 21775 14059
rect 22845 14025 22879 14059
rect 23489 14025 23523 14059
rect 24041 14025 24075 14059
rect 27905 14025 27939 14059
rect 6837 13957 6871 13991
rect 12449 13957 12483 13991
rect 28273 13957 28307 13991
rect 2513 13889 2547 13923
rect 4261 13889 4295 13923
rect 4997 13889 5031 13923
rect 5825 13889 5859 13923
rect 7389 13889 7423 13923
rect 7849 13889 7883 13923
rect 8309 13889 8343 13923
rect 8401 13889 8435 13923
rect 13093 13889 13127 13923
rect 13461 13889 13495 13923
rect 15577 13889 15611 13923
rect 19165 13889 19199 13923
rect 20729 13889 20763 13923
rect 22201 13889 22235 13923
rect 22385 13889 22419 13923
rect 26801 13889 26835 13923
rect 27353 13889 27387 13923
rect 27537 13889 27571 13923
rect 2421 13821 2455 13855
rect 4077 13821 4111 13855
rect 6285 13821 6319 13855
rect 7205 13821 7239 13855
rect 7297 13821 7331 13855
rect 8668 13821 8702 13855
rect 10701 13821 10735 13855
rect 12909 13821 12943 13855
rect 13829 13821 13863 13855
rect 15485 13821 15519 13855
rect 16221 13821 16255 13855
rect 19073 13821 19107 13855
rect 20085 13821 20119 13855
rect 20637 13821 20671 13855
rect 24409 13821 24443 13855
rect 5549 13753 5583 13787
rect 11345 13753 11379 13787
rect 21189 13753 21223 13787
rect 24654 13753 24688 13787
rect 26433 13753 26467 13787
rect 27261 13753 27295 13787
rect 1961 13685 1995 13719
rect 2329 13685 2363 13719
rect 3341 13685 3375 13719
rect 3985 13685 4019 13719
rect 5181 13685 5215 13719
rect 5641 13685 5675 13719
rect 12265 13685 12299 13719
rect 12817 13685 12851 13719
rect 15393 13685 15427 13719
rect 16957 13685 16991 13719
rect 18981 13685 19015 13719
rect 20545 13685 20579 13719
rect 22109 13685 22143 13719
rect 25789 13685 25823 13719
rect 26893 13685 26927 13719
rect 4813 13481 4847 13515
rect 5181 13481 5215 13515
rect 5825 13481 5859 13515
rect 6193 13481 6227 13515
rect 8493 13481 8527 13515
rect 8861 13481 8895 13515
rect 9229 13481 9263 13515
rect 10241 13481 10275 13515
rect 12725 13481 12759 13515
rect 13093 13481 13127 13515
rect 15025 13481 15059 13515
rect 15761 13481 15795 13515
rect 19349 13481 19383 13515
rect 20361 13481 20395 13515
rect 23213 13481 23247 13515
rect 23857 13481 23891 13515
rect 25329 13481 25363 13515
rect 26341 13481 26375 13515
rect 26525 13481 26559 13515
rect 26985 13481 27019 13515
rect 27629 13481 27663 13515
rect 1676 13413 1710 13447
rect 3709 13413 3743 13447
rect 6644 13413 6678 13447
rect 11529 13413 11563 13447
rect 17316 13413 17350 13447
rect 19717 13413 19751 13447
rect 1409 13345 1443 13379
rect 4353 13345 4387 13379
rect 14749 13345 14783 13379
rect 15669 13345 15703 13379
rect 17049 13345 17083 13379
rect 21189 13345 21223 13379
rect 21548 13345 21582 13379
rect 23949 13345 23983 13379
rect 24216 13345 24250 13379
rect 26893 13345 26927 13379
rect 5273 13277 5307 13311
rect 5457 13277 5491 13311
rect 6377 13277 6411 13311
rect 11621 13277 11655 13311
rect 11713 13277 11747 13311
rect 13185 13277 13219 13311
rect 13369 13277 13403 13311
rect 15853 13277 15887 13311
rect 19809 13277 19843 13311
rect 21281 13277 21315 13311
rect 27077 13277 27111 13311
rect 4721 13209 4755 13243
rect 15301 13209 15335 13243
rect 2789 13141 2823 13175
rect 3341 13141 3375 13175
rect 7757 13141 7791 13175
rect 9965 13141 9999 13175
rect 11069 13141 11103 13175
rect 11161 13141 11195 13175
rect 12541 13141 12575 13175
rect 18429 13141 18463 13175
rect 20729 13141 20763 13175
rect 22661 13141 22695 13175
rect 2053 12937 2087 12971
rect 4077 12937 4111 12971
rect 4721 12937 4755 12971
rect 6377 12937 6411 12971
rect 8309 12937 8343 12971
rect 9689 12937 9723 12971
rect 11253 12937 11287 12971
rect 13461 12937 13495 12971
rect 14841 12937 14875 12971
rect 15025 12937 15059 12971
rect 16037 12937 16071 12971
rect 17141 12937 17175 12971
rect 17509 12937 17543 12971
rect 18613 12937 18647 12971
rect 20453 12937 20487 12971
rect 21741 12937 21775 12971
rect 21833 12937 21867 12971
rect 22017 12937 22051 12971
rect 23029 12937 23063 12971
rect 23857 12937 23891 12971
rect 24225 12937 24259 12971
rect 28089 12937 28123 12971
rect 2513 12869 2547 12903
rect 2697 12801 2731 12835
rect 5825 12801 5859 12835
rect 7573 12801 7607 12835
rect 7941 12801 7975 12835
rect 9873 12801 9907 12835
rect 13093 12801 13127 12835
rect 13921 12801 13955 12835
rect 14197 12801 14231 12835
rect 15485 12801 15519 12835
rect 15669 12801 15703 12835
rect 17785 12801 17819 12835
rect 19165 12801 19199 12835
rect 19625 12801 19659 12835
rect 20361 12801 20395 12835
rect 21005 12801 21039 12835
rect 1409 12733 1443 12767
rect 2964 12733 2998 12767
rect 7757 12733 7791 12767
rect 8953 12733 8987 12767
rect 10129 12733 10163 12767
rect 12265 12733 12299 12767
rect 12817 12733 12851 12767
rect 18981 12733 19015 12767
rect 20913 12733 20947 12767
rect 21557 12733 21591 12767
rect 5641 12665 5675 12699
rect 7297 12665 7331 12699
rect 23489 12869 23523 12903
rect 24593 12869 24627 12903
rect 27445 12869 27479 12903
rect 22569 12801 22603 12835
rect 27077 12801 27111 12835
rect 27629 12801 27663 12835
rect 24041 12733 24075 12767
rect 25145 12733 25179 12767
rect 25412 12733 25446 12767
rect 9321 12665 9355 12699
rect 12909 12665 12943 12699
rect 15393 12665 15427 12699
rect 18521 12665 18555 12699
rect 19073 12665 19107 12699
rect 21741 12665 21775 12699
rect 24961 12665 24995 12699
rect 1593 12597 1627 12631
rect 4997 12597 5031 12631
rect 5181 12597 5215 12631
rect 5549 12597 5583 12631
rect 6929 12597 6963 12631
rect 7389 12597 7423 12631
rect 7757 12597 7791 12631
rect 8493 12597 8527 12631
rect 11805 12597 11839 12631
rect 12449 12597 12483 12631
rect 16497 12597 16531 12631
rect 20821 12597 20855 12631
rect 22385 12597 22419 12631
rect 22477 12597 22511 12631
rect 26525 12597 26559 12631
rect 1685 12393 1719 12427
rect 3709 12393 3743 12427
rect 7113 12393 7147 12427
rect 9781 12393 9815 12427
rect 12725 12393 12759 12427
rect 15025 12393 15059 12427
rect 15485 12393 15519 12427
rect 16773 12393 16807 12427
rect 22293 12393 22327 12427
rect 22845 12393 22879 12427
rect 24685 12393 24719 12427
rect 25697 12393 25731 12427
rect 2789 12325 2823 12359
rect 5181 12325 5215 12359
rect 8125 12325 8159 12359
rect 11590 12325 11624 12359
rect 14749 12325 14783 12359
rect 18144 12325 18178 12359
rect 25053 12325 25087 12359
rect 2145 12257 2179 12291
rect 2697 12257 2731 12291
rect 4077 12257 4111 12291
rect 5917 12257 5951 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 9413 12257 9447 12291
rect 10149 12257 10183 12291
rect 11345 12257 11379 12291
rect 16681 12257 16715 12291
rect 17877 12257 17911 12291
rect 20913 12257 20947 12291
rect 21180 12257 21214 12291
rect 23581 12257 23615 12291
rect 24133 12257 24167 12291
rect 26893 12257 26927 12291
rect 2973 12189 3007 12223
rect 6009 12189 6043 12223
rect 6193 12189 6227 12223
rect 7757 12189 7791 12223
rect 10241 12189 10275 12223
rect 10333 12189 10367 12223
rect 16957 12189 16991 12223
rect 25145 12189 25179 12223
rect 25329 12189 25363 12223
rect 26985 12189 27019 12223
rect 27169 12189 27203 12223
rect 3433 12121 3467 12155
rect 5549 12121 5583 12155
rect 16313 12121 16347 12155
rect 26249 12121 26283 12155
rect 2329 12053 2363 12087
rect 4261 12053 4295 12087
rect 4721 12053 4755 12087
rect 6653 12053 6687 12087
rect 7021 12053 7055 12087
rect 8677 12053 8711 12087
rect 9045 12053 9079 12087
rect 11161 12053 11195 12087
rect 13277 12053 13311 12087
rect 16129 12053 16163 12087
rect 19257 12053 19291 12087
rect 20545 12053 20579 12087
rect 23765 12053 23799 12087
rect 24501 12053 24535 12087
rect 26525 12053 26559 12087
rect 1869 11849 1903 11883
rect 2329 11849 2363 11883
rect 3893 11849 3927 11883
rect 5457 11849 5491 11883
rect 8217 11849 8251 11883
rect 10057 11849 10091 11883
rect 10977 11849 11011 11883
rect 11345 11849 11379 11883
rect 11713 11849 11747 11883
rect 14657 11849 14691 11883
rect 15853 11849 15887 11883
rect 17877 11849 17911 11883
rect 21465 11849 21499 11883
rect 23121 11849 23155 11883
rect 23489 11849 23523 11883
rect 25053 11849 25087 11883
rect 28089 11849 28123 11883
rect 10609 11781 10643 11815
rect 16313 11781 16347 11815
rect 18245 11781 18279 11815
rect 18797 11781 18831 11815
rect 20913 11781 20947 11815
rect 21189 11781 21223 11815
rect 25973 11781 26007 11815
rect 2145 11713 2179 11747
rect 2789 11713 2823 11747
rect 2973 11713 3007 11747
rect 4077 11713 4111 11747
rect 7665 11713 7699 11747
rect 15485 11713 15519 11747
rect 17049 11713 17083 11747
rect 18981 11713 19015 11747
rect 2697 11645 2731 11679
rect 3341 11645 3375 11679
rect 8677 11645 8711 11679
rect 8933 11645 8967 11679
rect 15209 11645 15243 11679
rect 16865 11645 16899 11679
rect 4344 11577 4378 11611
rect 7573 11577 7607 11611
rect 14381 11577 14415 11611
rect 16773 11577 16807 11611
rect 19226 11577 19260 11611
rect 22017 11713 22051 11747
rect 24409 11713 24443 11747
rect 24501 11713 24535 11747
rect 26157 11713 26191 11747
rect 21925 11645 21959 11679
rect 22477 11645 22511 11679
rect 24317 11645 24351 11679
rect 26424 11645 26458 11679
rect 21833 11577 21867 11611
rect 25605 11577 25639 11611
rect 6009 11509 6043 11543
rect 6469 11509 6503 11543
rect 7113 11509 7147 11543
rect 7481 11509 7515 11543
rect 8493 11509 8527 11543
rect 14841 11509 14875 11543
rect 15301 11509 15335 11543
rect 16405 11509 16439 11543
rect 17509 11509 17543 11543
rect 20361 11509 20395 11543
rect 21189 11509 21223 11543
rect 21281 11509 21315 11543
rect 23949 11509 23983 11543
rect 27537 11509 27571 11543
rect 3709 11305 3743 11339
rect 4261 11305 4295 11339
rect 5825 11305 5859 11339
rect 6929 11305 6963 11339
rect 9321 11305 9355 11339
rect 10149 11305 10183 11339
rect 10517 11305 10551 11339
rect 10977 11305 11011 11339
rect 11437 11305 11471 11339
rect 14933 11305 14967 11339
rect 16037 11305 16071 11339
rect 16497 11305 16531 11339
rect 17049 11305 17083 11339
rect 17601 11305 17635 11339
rect 19257 11305 19291 11339
rect 19625 11305 19659 11339
rect 21373 11305 21407 11339
rect 22109 11305 22143 11339
rect 22753 11305 22787 11339
rect 23673 11305 23707 11339
rect 24317 11305 24351 11339
rect 24961 11305 24995 11339
rect 25329 11305 25363 11339
rect 26157 11305 26191 11339
rect 26985 11305 27019 11339
rect 2697 11237 2731 11271
rect 3433 11237 3467 11271
rect 4629 11237 4663 11271
rect 7288 11237 7322 11271
rect 11345 11237 11379 11271
rect 18981 11237 19015 11271
rect 19717 11237 19751 11271
rect 24225 11237 24259 11271
rect 25421 11237 25455 11271
rect 26893 11237 26927 11271
rect 2605 11169 2639 11203
rect 4077 11169 4111 11203
rect 5733 11169 5767 11203
rect 16405 11169 16439 11203
rect 17969 11169 18003 11203
rect 21189 11169 21223 11203
rect 22661 11169 22695 11203
rect 23305 11169 23339 11203
rect 1777 11101 1811 11135
rect 2145 11101 2179 11135
rect 2881 11101 2915 11135
rect 5917 11101 5951 11135
rect 7021 11101 7055 11135
rect 9689 11101 9723 11135
rect 11621 11101 11655 11135
rect 16681 11101 16715 11135
rect 18061 11101 18095 11135
rect 18245 11101 18279 11135
rect 19901 11101 19935 11135
rect 22937 11101 22971 11135
rect 24409 11101 24443 11135
rect 27077 11101 27111 11135
rect 2237 11033 2271 11067
rect 4997 11033 5031 11067
rect 5365 11033 5399 11067
rect 6469 11033 6503 11067
rect 8401 11033 8435 11067
rect 22293 11033 22327 11067
rect 23857 11033 23891 11067
rect 26525 11033 26559 11067
rect 8953 10965 8987 10999
rect 21833 10965 21867 10999
rect 2881 10761 2915 10795
rect 4721 10761 4755 10795
rect 5457 10761 5491 10795
rect 7113 10761 7147 10795
rect 8677 10761 8711 10795
rect 11253 10761 11287 10795
rect 11529 10761 11563 10795
rect 16037 10761 16071 10795
rect 16405 10761 16439 10795
rect 17233 10761 17267 10795
rect 18245 10761 18279 10795
rect 19073 10761 19107 10795
rect 19533 10761 19567 10795
rect 21281 10761 21315 10795
rect 23121 10761 23155 10795
rect 23489 10761 23523 10795
rect 27169 10761 27203 10795
rect 27905 10761 27939 10795
rect 17693 10693 17727 10727
rect 21189 10693 21223 10727
rect 26157 10693 26191 10727
rect 2237 10625 2271 10659
rect 2329 10625 2363 10659
rect 3341 10625 3375 10659
rect 7665 10625 7699 10659
rect 8125 10625 8159 10659
rect 9229 10625 9263 10659
rect 18705 10625 18739 10659
rect 20177 10625 20211 10659
rect 21833 10625 21867 10659
rect 23673 10625 23707 10659
rect 26709 10625 26743 10659
rect 27537 10625 27571 10659
rect 6285 10557 6319 10591
rect 7481 10557 7515 10591
rect 8585 10557 8619 10591
rect 9045 10557 9079 10591
rect 10241 10557 10275 10591
rect 10793 10557 10827 10591
rect 19993 10557 20027 10591
rect 25973 10557 26007 10591
rect 26525 10557 26559 10591
rect 1685 10489 1719 10523
rect 2145 10489 2179 10523
rect 3586 10489 3620 10523
rect 5825 10489 5859 10523
rect 19441 10489 19475 10523
rect 19901 10489 19935 10523
rect 21649 10489 21683 10523
rect 22661 10489 22695 10523
rect 23918 10489 23952 10523
rect 25605 10489 25639 10523
rect 26617 10489 26651 10523
rect 1777 10421 1811 10455
rect 3249 10421 3283 10455
rect 6653 10421 6687 10455
rect 7573 10421 7607 10455
rect 9137 10421 9171 10455
rect 9689 10421 9723 10455
rect 10425 10421 10459 10455
rect 16865 10421 16899 10455
rect 20637 10421 20671 10455
rect 21741 10421 21775 10455
rect 22385 10421 22419 10455
rect 25053 10421 25087 10455
rect 1593 10217 1627 10251
rect 2421 10217 2455 10251
rect 6745 10217 6779 10251
rect 7665 10217 7699 10251
rect 7849 10217 7883 10251
rect 11069 10217 11103 10251
rect 17969 10217 18003 10251
rect 18429 10217 18463 10251
rect 19349 10217 19383 10251
rect 19809 10217 19843 10251
rect 20085 10217 20119 10251
rect 21373 10217 21407 10251
rect 22017 10217 22051 10251
rect 22753 10217 22787 10251
rect 23397 10217 23431 10251
rect 26249 10217 26283 10251
rect 27077 10217 27111 10251
rect 2789 10149 2823 10183
rect 4629 10149 4663 10183
rect 8861 10149 8895 10183
rect 22109 10149 22143 10183
rect 1409 10081 1443 10115
rect 2329 10081 2363 10115
rect 2881 10081 2915 10115
rect 3801 10081 3835 10115
rect 4077 10081 4111 10115
rect 5621 10081 5655 10115
rect 8217 10081 8251 10115
rect 18337 10081 18371 10115
rect 23489 10081 23523 10115
rect 23756 10081 23790 10115
rect 26525 10081 26559 10115
rect 2973 10013 3007 10047
rect 5365 10013 5399 10047
rect 8309 10013 8343 10047
rect 8493 10013 8527 10047
rect 18521 10013 18555 10047
rect 22293 10013 22327 10047
rect 3433 9945 3467 9979
rect 20729 9945 20763 9979
rect 21649 9945 21683 9979
rect 1961 9877 1995 9911
rect 4261 9877 4295 9911
rect 5181 9877 5215 9911
rect 7297 9877 7331 9911
rect 24869 9877 24903 9911
rect 26709 9877 26743 9911
rect 19165 9673 19199 9707
rect 21649 9673 21683 9707
rect 26985 9673 27019 9707
rect 2697 9605 2731 9639
rect 4169 9605 4203 9639
rect 4813 9605 4847 9639
rect 5457 9605 5491 9639
rect 5825 9605 5859 9639
rect 6837 9605 6871 9639
rect 8401 9605 8435 9639
rect 9413 9605 9447 9639
rect 17141 9605 17175 9639
rect 18153 9605 18187 9639
rect 19717 9605 19751 9639
rect 23121 9605 23155 9639
rect 23857 9605 23891 9639
rect 26341 9605 26375 9639
rect 6653 9537 6687 9571
rect 7297 9537 7331 9571
rect 7481 9537 7515 9571
rect 8953 9537 8987 9571
rect 17785 9537 17819 9571
rect 18613 9537 18647 9571
rect 18797 9537 18831 9571
rect 20269 9537 20303 9571
rect 20821 9537 20855 9571
rect 22293 9537 22327 9571
rect 22661 9537 22695 9571
rect 23489 9537 23523 9571
rect 24501 9537 24535 9571
rect 1409 9469 1443 9503
rect 1961 9469 1995 9503
rect 2789 9469 2823 9503
rect 5273 9469 5307 9503
rect 7205 9469 7239 9503
rect 17509 9469 17543 9503
rect 20085 9469 20119 9503
rect 21189 9469 21223 9503
rect 22109 9469 22143 9503
rect 26433 9469 26467 9503
rect 27537 9469 27571 9503
rect 28089 9469 28123 9503
rect 3056 9401 3090 9435
rect 8309 9401 8343 9435
rect 8769 9401 8803 9435
rect 21465 9401 21499 9435
rect 22017 9401 22051 9435
rect 24225 9401 24259 9435
rect 1593 9333 1627 9367
rect 5089 9333 5123 9367
rect 6193 9333 6227 9367
rect 7849 9333 7883 9367
rect 8861 9333 8895 9367
rect 18521 9333 18555 9367
rect 19625 9333 19659 9367
rect 20177 9333 20211 9367
rect 24317 9333 24351 9367
rect 26617 9333 26651 9367
rect 27721 9333 27755 9367
rect 1961 9129 1995 9163
rect 2329 9129 2363 9163
rect 2881 9129 2915 9163
rect 4077 9129 4111 9163
rect 5457 9129 5491 9163
rect 8125 9129 8159 9163
rect 8953 9129 8987 9163
rect 17877 9129 17911 9163
rect 18521 9129 18555 9163
rect 18981 9129 19015 9163
rect 19809 9129 19843 9163
rect 21741 9129 21775 9163
rect 22109 9129 22143 9163
rect 23949 9129 23983 9163
rect 24501 9129 24535 9163
rect 24869 9129 24903 9163
rect 24961 9129 24995 9163
rect 18153 9061 18187 9095
rect 24225 9061 24259 9095
rect 2789 8993 2823 9027
rect 3893 8993 3927 9027
rect 4445 8993 4479 9027
rect 5908 8993 5942 9027
rect 18889 8993 18923 9027
rect 26525 8993 26559 9027
rect 3065 8925 3099 8959
rect 4537 8925 4571 8959
rect 4721 8925 4755 8959
rect 5641 8925 5675 8959
rect 19165 8925 19199 8959
rect 23581 8925 23615 8959
rect 25145 8925 25179 8959
rect 3433 8857 3467 8891
rect 2421 8789 2455 8823
rect 5089 8789 5123 8823
rect 7021 8789 7055 8823
rect 7849 8789 7883 8823
rect 8585 8789 8619 8823
rect 26709 8789 26743 8823
rect 2605 8585 2639 8619
rect 6837 8585 6871 8619
rect 18613 8585 18647 8619
rect 18889 8585 18923 8619
rect 19257 8585 19291 8619
rect 24133 8585 24167 8619
rect 25237 8585 25271 8619
rect 25513 8585 25547 8619
rect 27353 8585 27387 8619
rect 27721 8585 27755 8619
rect 4629 8517 4663 8551
rect 24409 8517 24443 8551
rect 26617 8517 26651 8551
rect 27077 8517 27111 8551
rect 1961 8449 1995 8483
rect 2053 8449 2087 8483
rect 3617 8449 3651 8483
rect 4169 8449 4203 8483
rect 4537 8449 4571 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 7389 8449 7423 8483
rect 24869 8449 24903 8483
rect 1869 8381 1903 8415
rect 2973 8381 3007 8415
rect 3433 8381 3467 8415
rect 4997 8381 5031 8415
rect 7205 8381 7239 8415
rect 8217 8381 8251 8415
rect 24225 8381 24259 8415
rect 25329 8381 25363 8415
rect 25881 8381 25915 8415
rect 26433 8381 26467 8415
rect 27537 8381 27571 8415
rect 28089 8381 28123 8415
rect 3525 8313 3559 8347
rect 5733 8313 5767 8347
rect 6101 8313 6135 8347
rect 7297 8313 7331 8347
rect 7849 8313 7883 8347
rect 1501 8245 1535 8279
rect 3065 8245 3099 8279
rect 6561 8245 6595 8279
rect 1685 8041 1719 8075
rect 2145 8041 2179 8075
rect 2789 8041 2823 8075
rect 3525 8041 3559 8075
rect 3893 8041 3927 8075
rect 4261 8041 4295 8075
rect 5273 8041 5307 8075
rect 5641 8041 5675 8075
rect 24593 8041 24627 8075
rect 25513 8041 25547 8075
rect 3157 7973 3191 8007
rect 2053 7905 2087 7939
rect 4077 7905 4111 7939
rect 5733 7905 5767 7939
rect 7205 7905 7239 7939
rect 25329 7905 25363 7939
rect 26525 7905 26559 7939
rect 2237 7837 2271 7871
rect 5825 7837 5859 7871
rect 7297 7837 7331 7871
rect 7481 7837 7515 7871
rect 4813 7769 4847 7803
rect 5089 7701 5123 7735
rect 6837 7701 6871 7735
rect 26709 7701 26743 7735
rect 3065 7497 3099 7531
rect 4169 7497 4203 7531
rect 4905 7497 4939 7531
rect 5917 7497 5951 7531
rect 6561 7497 6595 7531
rect 6837 7497 6871 7531
rect 25329 7497 25363 7531
rect 27353 7497 27387 7531
rect 1593 7429 1627 7463
rect 2329 7429 2363 7463
rect 27721 7429 27755 7463
rect 2973 7361 3007 7395
rect 3617 7361 3651 7395
rect 5365 7361 5399 7395
rect 5457 7361 5491 7395
rect 7297 7361 7331 7395
rect 7481 7361 7515 7395
rect 1409 7293 1443 7327
rect 1961 7293 1995 7327
rect 3525 7293 3559 7327
rect 4813 7293 4847 7327
rect 5273 7293 5307 7327
rect 26433 7293 26467 7327
rect 26985 7293 27019 7327
rect 27537 7293 27571 7327
rect 28089 7293 28123 7327
rect 3433 7157 3467 7191
rect 7205 7157 7239 7191
rect 7849 7157 7883 7191
rect 8309 7157 8343 7191
rect 26617 7157 26651 7191
rect 3433 6953 3467 6987
rect 3801 6953 3835 6987
rect 4997 6953 5031 6987
rect 5457 6953 5491 6987
rect 7205 6953 7239 6987
rect 7665 6885 7699 6919
rect 1409 6817 1443 6851
rect 1961 6817 1995 6851
rect 2513 6817 2547 6851
rect 4077 6817 4111 6851
rect 5365 6817 5399 6851
rect 5825 6817 5859 6851
rect 26525 6817 26559 6851
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 5917 6749 5951 6783
rect 6101 6749 6135 6783
rect 1593 6681 1627 6715
rect 2697 6681 2731 6715
rect 4261 6613 4295 6647
rect 6929 6613 6963 6647
rect 26709 6613 26743 6647
rect 2421 6409 2455 6443
rect 3157 6409 3191 6443
rect 4261 6409 4295 6443
rect 5549 6409 5583 6443
rect 6285 6409 6319 6443
rect 26617 6409 26651 6443
rect 1593 6341 1627 6375
rect 2053 6341 2087 6375
rect 26985 6341 27019 6375
rect 26341 6273 26375 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 3525 6205 3559 6239
rect 3617 6205 3651 6239
rect 26433 6205 26467 6239
rect 2697 6069 2731 6103
rect 3801 6069 3835 6103
rect 5825 6069 5859 6103
rect 2053 5865 2087 5899
rect 2421 5865 2455 5899
rect 3617 5865 3651 5899
rect 3065 5797 3099 5831
rect 1409 5729 1443 5763
rect 2513 5729 2547 5763
rect 26525 5729 26559 5763
rect 1593 5593 1627 5627
rect 26709 5593 26743 5627
rect 2697 5525 2731 5559
rect 2513 5321 2547 5355
rect 27353 5321 27387 5355
rect 2053 5185 2087 5219
rect 1409 5117 1443 5151
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 1593 4981 1627 5015
rect 26617 4981 26651 5015
rect 1685 4777 1719 4811
rect 2053 3145 2087 3179
rect 1409 2941 1443 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 1593 2805 1627 2839
rect 26617 2805 26651 2839
rect 8309 2601 8343 2635
rect 6745 2465 6779 2499
rect 7196 2465 7230 2499
rect 6929 2397 6963 2431
rect 6285 2261 6319 2295
<< metal1 >>
rect 3326 22516 3332 22568
rect 3384 22556 3390 22568
rect 7926 22556 7932 22568
rect 3384 22528 7932 22556
rect 3384 22516 3390 22528
rect 7926 22516 7932 22528
rect 7984 22516 7990 22568
rect 2958 22108 2964 22160
rect 3016 22148 3022 22160
rect 13630 22148 13636 22160
rect 3016 22120 13636 22148
rect 3016 22108 3022 22120
rect 13630 22108 13636 22120
rect 13688 22108 13694 22160
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 24305 21131 24363 21137
rect 24305 21097 24317 21131
rect 24351 21097 24363 21131
rect 24305 21091 24363 21097
rect 25317 21131 25375 21137
rect 25317 21097 25329 21131
rect 25363 21128 25375 21131
rect 27154 21128 27160 21140
rect 25363 21100 27160 21128
rect 25363 21097 25375 21100
rect 25317 21091 25375 21097
rect 24320 21060 24348 21091
rect 27154 21088 27160 21100
rect 27212 21088 27218 21140
rect 28994 21060 29000 21072
rect 24320 21032 29000 21060
rect 28994 21020 29000 21032
rect 29052 21020 29058 21072
rect 23842 20952 23848 21004
rect 23900 20992 23906 21004
rect 24121 20995 24179 21001
rect 24121 20992 24133 20995
rect 23900 20964 24133 20992
rect 23900 20952 23906 20964
rect 24121 20961 24133 20964
rect 24167 20961 24179 20995
rect 24121 20955 24179 20961
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20992 25191 20995
rect 25179 20964 26096 20992
rect 25179 20961 25191 20964
rect 25133 20955 25191 20961
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 5718 20788 5724 20800
rect 4120 20760 5724 20788
rect 4120 20748 4126 20760
rect 5718 20748 5724 20760
rect 5776 20748 5782 20800
rect 15562 20788 15568 20800
rect 15523 20760 15568 20788
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 19242 20788 19248 20800
rect 19203 20760 19248 20788
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 21266 20748 21272 20800
rect 21324 20788 21330 20800
rect 25498 20788 25504 20800
rect 21324 20760 25504 20788
rect 21324 20748 21330 20760
rect 25498 20748 25504 20760
rect 25556 20748 25562 20800
rect 25685 20791 25743 20797
rect 25685 20757 25697 20791
rect 25731 20788 25743 20791
rect 25774 20788 25780 20800
rect 25731 20760 25780 20788
rect 25731 20757 25743 20760
rect 25685 20751 25743 20757
rect 25774 20748 25780 20760
rect 25832 20748 25838 20800
rect 26068 20797 26096 20964
rect 26053 20791 26111 20797
rect 26053 20757 26065 20791
rect 26099 20788 26111 20791
rect 26602 20788 26608 20800
rect 26099 20760 26608 20788
rect 26099 20757 26111 20760
rect 26053 20751 26111 20757
rect 26602 20748 26608 20760
rect 26660 20748 26666 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 992 20556 1593 20584
rect 992 20544 998 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 7101 20587 7159 20593
rect 7101 20553 7113 20587
rect 7147 20584 7159 20587
rect 8202 20584 8208 20596
rect 7147 20556 8208 20584
rect 7147 20553 7159 20556
rect 7101 20547 7159 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 9493 20587 9551 20593
rect 9493 20553 9505 20587
rect 9539 20584 9551 20587
rect 10226 20584 10232 20596
rect 9539 20556 10232 20584
rect 9539 20553 9551 20556
rect 9493 20547 9551 20553
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 12621 20587 12679 20593
rect 12621 20553 12633 20587
rect 12667 20584 12679 20587
rect 13998 20584 14004 20596
rect 12667 20556 14004 20584
rect 12667 20553 12679 20556
rect 12621 20547 12679 20553
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 15838 20584 15844 20596
rect 14323 20556 15844 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 17129 20587 17187 20593
rect 17129 20553 17141 20587
rect 17175 20584 17187 20587
rect 17770 20584 17776 20596
rect 17175 20556 17776 20584
rect 17175 20553 17187 20556
rect 17129 20547 17187 20553
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 19610 20584 19616 20596
rect 18279 20556 19616 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 19610 20544 19616 20556
rect 19668 20544 19674 20596
rect 20901 20587 20959 20593
rect 20901 20553 20913 20587
rect 20947 20584 20959 20587
rect 21542 20584 21548 20596
rect 20947 20556 21548 20584
rect 20947 20553 20959 20556
rect 20901 20547 20959 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 24397 20587 24455 20593
rect 24397 20553 24409 20587
rect 24443 20584 24455 20587
rect 25222 20584 25228 20596
rect 24443 20556 25228 20584
rect 24443 20553 24455 20556
rect 24397 20547 24455 20553
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 4982 20516 4988 20528
rect 4943 20488 4988 20516
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 15620 20420 15669 20448
rect 15620 20408 15626 20420
rect 15657 20417 15669 20420
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 19242 20408 19248 20460
rect 19300 20448 19306 20460
rect 19702 20448 19708 20460
rect 19300 20420 19708 20448
rect 19300 20408 19306 20420
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 25409 20451 25467 20457
rect 25409 20417 25421 20451
rect 25455 20448 25467 20451
rect 26142 20448 26148 20460
rect 25455 20420 26148 20448
rect 25455 20417 25467 20420
rect 25409 20411 25467 20417
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1443 20352 1992 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1964 20253 1992 20352
rect 4154 20340 4160 20392
rect 4212 20380 4218 20392
rect 4801 20383 4859 20389
rect 4801 20380 4813 20383
rect 4212 20352 4813 20380
rect 4212 20340 4218 20352
rect 4801 20349 4813 20352
rect 4847 20380 4859 20383
rect 5261 20383 5319 20389
rect 5261 20380 5273 20383
rect 4847 20352 5273 20380
rect 4847 20349 4859 20352
rect 4801 20343 4859 20349
rect 5261 20349 5273 20352
rect 5307 20349 5319 20383
rect 5261 20343 5319 20349
rect 6917 20383 6975 20389
rect 6917 20349 6929 20383
rect 6963 20380 6975 20383
rect 9309 20383 9367 20389
rect 6963 20352 7512 20380
rect 6963 20349 6975 20352
rect 6917 20343 6975 20349
rect 1949 20247 2007 20253
rect 1949 20213 1961 20247
rect 1995 20244 2007 20247
rect 2406 20244 2412 20256
rect 1995 20216 2412 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 7484 20253 7512 20352
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 9355 20352 9904 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 7469 20247 7527 20253
rect 7469 20213 7481 20247
rect 7515 20244 7527 20247
rect 7834 20244 7840 20256
rect 7515 20216 7840 20244
rect 7515 20213 7527 20216
rect 7469 20207 7527 20213
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 9876 20253 9904 20352
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 12897 20383 12955 20389
rect 12897 20380 12909 20383
rect 12492 20352 12909 20380
rect 12492 20340 12498 20352
rect 12897 20349 12909 20352
rect 12943 20349 12955 20383
rect 14093 20383 14151 20389
rect 14093 20380 14105 20383
rect 12897 20343 12955 20349
rect 14016 20352 14105 20380
rect 14016 20256 14044 20352
rect 14093 20349 14105 20352
rect 14139 20349 14151 20383
rect 14093 20343 14151 20349
rect 14918 20340 14924 20392
rect 14976 20380 14982 20392
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 14976 20352 15485 20380
rect 14976 20340 14982 20352
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 15473 20343 15531 20349
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20380 17003 20383
rect 18046 20380 18052 20392
rect 16991 20352 17540 20380
rect 18007 20352 18052 20380
rect 16991 20349 17003 20352
rect 16945 20343 17003 20349
rect 14550 20312 14556 20324
rect 14511 20284 14556 20312
rect 14550 20272 14556 20284
rect 14608 20312 14614 20324
rect 15565 20315 15623 20321
rect 15565 20312 15577 20315
rect 14608 20284 15577 20312
rect 14608 20272 14614 20284
rect 15565 20281 15577 20284
rect 15611 20312 15623 20315
rect 16390 20312 16396 20324
rect 15611 20284 16396 20312
rect 15611 20281 15623 20284
rect 15565 20275 15623 20281
rect 16390 20272 16396 20284
rect 16448 20272 16454 20324
rect 17512 20256 17540 20352
rect 18046 20340 18052 20352
rect 18104 20380 18110 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18104 20352 18521 20380
rect 18104 20340 18110 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 20714 20380 20720 20392
rect 20675 20352 20720 20380
rect 18509 20343 18567 20349
rect 20714 20340 20720 20352
rect 20772 20380 20778 20392
rect 21177 20383 21235 20389
rect 21177 20380 21189 20383
rect 20772 20352 21189 20380
rect 20772 20340 20778 20352
rect 21177 20349 21189 20352
rect 21223 20349 21235 20383
rect 24213 20383 24271 20389
rect 24213 20380 24225 20383
rect 21177 20343 21235 20349
rect 24136 20352 24225 20380
rect 19061 20315 19119 20321
rect 19061 20281 19073 20315
rect 19107 20312 19119 20315
rect 19107 20284 19564 20312
rect 19107 20281 19119 20284
rect 19061 20275 19119 20281
rect 19536 20256 19564 20284
rect 24136 20256 24164 20352
rect 24213 20349 24225 20352
rect 24259 20349 24271 20383
rect 24213 20343 24271 20349
rect 25774 20272 25780 20324
rect 25832 20312 25838 20324
rect 25961 20315 26019 20321
rect 25961 20312 25973 20315
rect 25832 20284 25973 20312
rect 25832 20272 25838 20284
rect 25961 20281 25973 20284
rect 26007 20281 26019 20315
rect 25961 20275 26019 20281
rect 9861 20247 9919 20253
rect 9861 20213 9873 20247
rect 9907 20244 9919 20247
rect 9950 20244 9956 20256
rect 9907 20216 9956 20244
rect 9907 20213 9919 20216
rect 9861 20207 9919 20213
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 13998 20244 14004 20256
rect 13959 20216 14004 20244
rect 13998 20204 14004 20216
rect 14056 20204 14062 20256
rect 14918 20244 14924 20256
rect 14879 20216 14924 20244
rect 14918 20204 14924 20216
rect 14976 20204 14982 20256
rect 15102 20244 15108 20256
rect 15063 20216 15108 20244
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 17494 20244 17500 20256
rect 17455 20216 17500 20244
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 19150 20244 19156 20256
rect 19111 20216 19156 20244
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 19518 20244 19524 20256
rect 19479 20216 19524 20244
rect 19518 20204 19524 20216
rect 19576 20204 19582 20256
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 23477 20247 23535 20253
rect 19668 20216 19713 20244
rect 19668 20204 19674 20216
rect 23477 20213 23489 20247
rect 23523 20244 23535 20247
rect 23842 20244 23848 20256
rect 23523 20216 23848 20244
rect 23523 20213 23535 20216
rect 23477 20207 23535 20213
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 24118 20244 24124 20256
rect 24079 20216 24124 20244
rect 24118 20204 24124 20216
rect 24176 20204 24182 20256
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20244 25007 20247
rect 25222 20244 25228 20256
rect 24995 20216 25228 20244
rect 24995 20213 25007 20216
rect 24949 20207 25007 20213
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 25498 20244 25504 20256
rect 25459 20216 25504 20244
rect 25498 20204 25504 20216
rect 25556 20204 25562 20256
rect 25866 20244 25872 20256
rect 25827 20216 25872 20244
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 15102 20000 15108 20052
rect 15160 20040 15166 20052
rect 15470 20040 15476 20052
rect 15160 20012 15476 20040
rect 15160 20000 15166 20012
rect 15470 20000 15476 20012
rect 15528 20040 15534 20052
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 15528 20012 15761 20040
rect 15528 20000 15534 20012
rect 15749 20009 15761 20012
rect 15795 20009 15807 20043
rect 15749 20003 15807 20009
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 17773 20043 17831 20049
rect 17773 20040 17785 20043
rect 17552 20012 17785 20040
rect 17552 20000 17558 20012
rect 17773 20009 17785 20012
rect 17819 20009 17831 20043
rect 17773 20003 17831 20009
rect 24029 19975 24087 19981
rect 24029 19941 24041 19975
rect 24075 19972 24087 19975
rect 25498 19972 25504 19984
rect 24075 19944 25504 19972
rect 24075 19941 24087 19944
rect 24029 19935 24087 19941
rect 25498 19932 25504 19944
rect 25556 19932 25562 19984
rect 11606 19864 11612 19916
rect 11664 19904 11670 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 11664 19876 12357 19904
rect 11664 19864 11670 19876
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 12345 19867 12403 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15657 19907 15715 19913
rect 15657 19904 15669 19907
rect 15252 19876 15669 19904
rect 15252 19864 15258 19876
rect 15657 19873 15669 19876
rect 15703 19904 15715 19907
rect 16482 19904 16488 19916
rect 15703 19876 16488 19904
rect 15703 19873 15715 19876
rect 15657 19867 15715 19873
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 18138 19904 18144 19916
rect 18099 19876 18144 19904
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 24394 19864 24400 19916
rect 24452 19904 24458 19916
rect 25038 19904 25044 19916
rect 24452 19876 25044 19904
rect 24452 19864 24458 19876
rect 25038 19864 25044 19876
rect 25096 19864 25102 19916
rect 25222 19904 25228 19916
rect 25183 19876 25228 19904
rect 25222 19864 25228 19876
rect 25280 19864 25286 19916
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 11808 19808 12449 19836
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 8665 19703 8723 19709
rect 8665 19669 8677 19703
rect 8711 19700 8723 19703
rect 9030 19700 9036 19712
rect 8711 19672 9036 19700
rect 8711 19669 8723 19672
rect 8665 19663 8723 19669
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 10870 19700 10876 19712
rect 10831 19672 10876 19700
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 11422 19660 11428 19712
rect 11480 19700 11486 19712
rect 11808 19709 11836 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 15838 19836 15844 19848
rect 12584 19808 12629 19836
rect 15799 19808 15844 19836
rect 12584 19796 12590 19808
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 18230 19836 18236 19848
rect 18191 19808 18236 19836
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19836 18475 19839
rect 18598 19836 18604 19848
rect 18463 19808 18604 19836
rect 18463 19805 18475 19808
rect 18417 19799 18475 19805
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 25317 19839 25375 19845
rect 25317 19805 25329 19839
rect 25363 19805 25375 19839
rect 25317 19799 25375 19805
rect 24397 19771 24455 19777
rect 24397 19737 24409 19771
rect 24443 19768 24455 19771
rect 24857 19771 24915 19777
rect 24857 19768 24869 19771
rect 24443 19740 24869 19768
rect 24443 19737 24455 19740
rect 24397 19731 24455 19737
rect 24857 19737 24869 19740
rect 24903 19768 24915 19771
rect 25038 19768 25044 19780
rect 24903 19740 25044 19768
rect 24903 19737 24915 19740
rect 24857 19731 24915 19737
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 11793 19703 11851 19709
rect 11793 19700 11805 19703
rect 11480 19672 11805 19700
rect 11480 19660 11486 19672
rect 11793 19669 11805 19672
rect 11839 19669 11851 19703
rect 11974 19700 11980 19712
rect 11935 19672 11980 19700
rect 11793 19663 11851 19669
rect 11974 19660 11980 19672
rect 12032 19660 12038 19712
rect 12802 19660 12808 19712
rect 12860 19700 12866 19712
rect 12989 19703 13047 19709
rect 12989 19700 13001 19703
rect 12860 19672 13001 19700
rect 12860 19660 12866 19672
rect 12989 19669 13001 19672
rect 13035 19669 13047 19703
rect 12989 19663 13047 19669
rect 15013 19703 15071 19709
rect 15013 19669 15025 19703
rect 15059 19700 15071 19703
rect 15286 19700 15292 19712
rect 15059 19672 15292 19700
rect 15059 19669 15071 19672
rect 15013 19663 15071 19669
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 19153 19703 19211 19709
rect 19153 19700 19165 19703
rect 18380 19672 19165 19700
rect 18380 19660 18386 19672
rect 19153 19669 19165 19672
rect 19199 19700 19211 19703
rect 19610 19700 19616 19712
rect 19199 19672 19616 19700
rect 19199 19669 19211 19672
rect 19153 19663 19211 19669
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 24762 19700 24768 19712
rect 24723 19672 24768 19700
rect 24762 19660 24768 19672
rect 24820 19700 24826 19712
rect 25332 19700 25360 19799
rect 25406 19796 25412 19848
rect 25464 19836 25470 19848
rect 25501 19839 25559 19845
rect 25501 19836 25513 19839
rect 25464 19808 25513 19836
rect 25464 19796 25470 19808
rect 25501 19805 25513 19808
rect 25547 19836 25559 19839
rect 26142 19836 26148 19848
rect 25547 19808 26148 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 26510 19836 26516 19848
rect 26471 19808 26516 19836
rect 26510 19796 26516 19808
rect 26568 19796 26574 19848
rect 25866 19700 25872 19712
rect 24820 19672 25360 19700
rect 25827 19672 25872 19700
rect 24820 19660 24826 19672
rect 25866 19660 25872 19672
rect 25924 19660 25930 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 13998 19456 14004 19508
rect 14056 19496 14062 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14056 19468 14933 19496
rect 14056 19456 14062 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 14921 19459 14979 19465
rect 24118 19456 24124 19508
rect 24176 19496 24182 19508
rect 24581 19499 24639 19505
rect 24581 19496 24593 19499
rect 24176 19468 24593 19496
rect 24176 19456 24182 19468
rect 24581 19465 24593 19468
rect 24627 19465 24639 19499
rect 25406 19496 25412 19508
rect 24581 19459 24639 19465
rect 24780 19468 25412 19496
rect 8754 19388 8760 19440
rect 8812 19428 8818 19440
rect 9582 19428 9588 19440
rect 8812 19400 9588 19428
rect 8812 19388 8818 19400
rect 9582 19388 9588 19400
rect 9640 19388 9646 19440
rect 10689 19431 10747 19437
rect 10689 19397 10701 19431
rect 10735 19428 10747 19431
rect 10735 19400 11376 19428
rect 10735 19397 10747 19400
rect 10689 19391 10747 19397
rect 11348 19372 11376 19400
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 8527 19332 9137 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 9125 19329 9137 19332
rect 9171 19360 9183 19363
rect 9490 19360 9496 19372
rect 9171 19332 9496 19360
rect 9171 19329 9183 19332
rect 9125 19323 9183 19329
rect 9490 19320 9496 19332
rect 9548 19320 9554 19372
rect 10870 19320 10876 19372
rect 10928 19360 10934 19372
rect 11330 19360 11336 19372
rect 10928 19332 11008 19360
rect 11243 19332 11336 19360
rect 10928 19320 10934 19332
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 3050 19292 3056 19304
rect 2823 19264 3056 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 3050 19252 3056 19264
rect 3108 19292 3114 19304
rect 3605 19295 3663 19301
rect 3605 19292 3617 19295
rect 3108 19264 3617 19292
rect 3108 19252 3114 19264
rect 3605 19261 3617 19264
rect 3651 19261 3663 19295
rect 10980 19292 11008 19332
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12584 19332 13001 19360
rect 12584 19320 12590 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 15473 19363 15531 19369
rect 15473 19360 15485 19363
rect 12989 19323 13047 19329
rect 15120 19332 15485 19360
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 10980 19264 11253 19292
rect 3605 19255 3663 19261
rect 11241 19261 11253 19264
rect 11287 19292 11299 19295
rect 12342 19292 12348 19304
rect 11287 19264 12348 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 12802 19292 12808 19304
rect 12763 19264 12808 19292
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 14829 19295 14887 19301
rect 14829 19261 14841 19295
rect 14875 19292 14887 19295
rect 15120 19292 15148 19332
rect 15473 19329 15485 19332
rect 15519 19360 15531 19363
rect 16482 19360 16488 19372
rect 15519 19332 16488 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 18230 19360 18236 19372
rect 17880 19332 18236 19360
rect 15286 19292 15292 19304
rect 14875 19264 15148 19292
rect 15247 19264 15292 19292
rect 14875 19261 14887 19264
rect 14829 19255 14887 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 17880 19292 17908 19332
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 17543 19264 17908 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 19024 19264 19073 19292
rect 19024 19252 19030 19264
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 21818 19292 21824 19304
rect 21779 19264 21824 19292
rect 19061 19255 19119 19261
rect 21818 19252 21824 19264
rect 21876 19292 21882 19304
rect 22281 19295 22339 19301
rect 22281 19292 22293 19295
rect 21876 19264 22293 19292
rect 21876 19252 21882 19264
rect 22281 19261 22293 19264
rect 22327 19261 22339 19295
rect 22281 19255 22339 19261
rect 24121 19295 24179 19301
rect 24121 19261 24133 19295
rect 24167 19292 24179 19295
rect 24210 19292 24216 19304
rect 24167 19264 24216 19292
rect 24167 19261 24179 19264
rect 24121 19255 24179 19261
rect 24210 19252 24216 19264
rect 24268 19292 24274 19304
rect 24780 19292 24808 19468
rect 25406 19456 25412 19468
rect 25464 19456 25470 19508
rect 25866 19456 25872 19508
rect 25924 19496 25930 19508
rect 26329 19499 26387 19505
rect 26329 19496 26341 19499
rect 25924 19468 26341 19496
rect 25924 19456 25930 19468
rect 26329 19465 26341 19468
rect 26375 19465 26387 19499
rect 26329 19459 26387 19465
rect 25498 19428 25504 19440
rect 24268 19264 24808 19292
rect 24872 19400 25504 19428
rect 24872 19292 24900 19400
rect 25498 19388 25504 19400
rect 25556 19388 25562 19440
rect 25038 19360 25044 19372
rect 24999 19332 25044 19360
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 25133 19363 25191 19369
rect 25133 19329 25145 19363
rect 25179 19329 25191 19363
rect 25133 19323 25191 19329
rect 26973 19363 27031 19369
rect 26973 19329 26985 19363
rect 27019 19360 27031 19363
rect 27338 19360 27344 19372
rect 27019 19332 27344 19360
rect 27019 19329 27031 19332
rect 26973 19323 27031 19329
rect 24949 19295 25007 19301
rect 24949 19292 24961 19295
rect 24872 19264 24961 19292
rect 24268 19252 24274 19264
rect 24949 19261 24961 19264
rect 24995 19261 25007 19295
rect 24949 19255 25007 19261
rect 1673 19227 1731 19233
rect 1673 19193 1685 19227
rect 1719 19224 1731 19227
rect 2130 19224 2136 19236
rect 1719 19196 2136 19224
rect 1719 19193 1731 19196
rect 1673 19187 1731 19193
rect 2130 19184 2136 19196
rect 2188 19184 2194 19236
rect 8113 19227 8171 19233
rect 8113 19193 8125 19227
rect 8159 19224 8171 19227
rect 8941 19227 8999 19233
rect 8941 19224 8953 19227
rect 8159 19196 8953 19224
rect 8159 19193 8171 19196
rect 8113 19187 8171 19193
rect 8941 19193 8953 19196
rect 8987 19224 8999 19227
rect 9582 19224 9588 19236
rect 8987 19196 9588 19224
rect 8987 19193 8999 19196
rect 8941 19187 8999 19193
rect 9582 19184 9588 19196
rect 9640 19184 9646 19236
rect 10321 19227 10379 19233
rect 10321 19193 10333 19227
rect 10367 19224 10379 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10367 19196 11161 19224
rect 10367 19193 10379 19196
rect 10321 19187 10379 19193
rect 11149 19193 11161 19196
rect 11195 19224 11207 19227
rect 14461 19227 14519 19233
rect 11195 19196 12480 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 1762 19156 1768 19168
rect 1723 19128 1768 19156
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 1946 19116 1952 19168
rect 2004 19156 2010 19168
rect 2225 19159 2283 19165
rect 2225 19156 2237 19159
rect 2004 19128 2237 19156
rect 2004 19116 2010 19128
rect 2225 19125 2237 19128
rect 2271 19125 2283 19159
rect 2958 19156 2964 19168
rect 2919 19128 2964 19156
rect 2225 19119 2283 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3234 19156 3240 19168
rect 3195 19128 3240 19156
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 8570 19156 8576 19168
rect 8531 19128 8576 19156
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 9030 19156 9036 19168
rect 8991 19128 9036 19156
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 10686 19116 10692 19168
rect 10744 19156 10750 19168
rect 10781 19159 10839 19165
rect 10781 19156 10793 19159
rect 10744 19128 10793 19156
rect 10744 19116 10750 19128
rect 10781 19125 10793 19128
rect 10827 19125 10839 19159
rect 10781 19119 10839 19125
rect 11606 19116 11612 19168
rect 11664 19156 11670 19168
rect 12452 19165 12480 19196
rect 14461 19193 14473 19227
rect 14507 19224 14519 19227
rect 15102 19224 15108 19236
rect 14507 19196 15108 19224
rect 14507 19193 14519 19196
rect 14461 19187 14519 19193
rect 15102 19184 15108 19196
rect 15160 19184 15166 19236
rect 17129 19227 17187 19233
rect 17129 19193 17141 19227
rect 17175 19224 17187 19227
rect 18138 19224 18144 19236
rect 17175 19196 18144 19224
rect 17175 19193 17187 19196
rect 17129 19187 17187 19193
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18598 19224 18604 19236
rect 18432 19196 18604 19224
rect 11977 19159 12035 19165
rect 11977 19156 11989 19159
rect 11664 19128 11989 19156
rect 11664 19116 11670 19128
rect 11977 19125 11989 19128
rect 12023 19125 12035 19159
rect 11977 19119 12035 19125
rect 12437 19159 12495 19165
rect 12437 19125 12449 19159
rect 12483 19125 12495 19159
rect 12894 19156 12900 19168
rect 12807 19128 12900 19156
rect 12437 19119 12495 19125
rect 12894 19116 12900 19128
rect 12952 19156 12958 19168
rect 13538 19156 13544 19168
rect 12952 19128 13544 19156
rect 12952 19116 12958 19128
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 13906 19156 13912 19168
rect 13867 19128 13912 19156
rect 13906 19116 13912 19128
rect 13964 19116 13970 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 15252 19128 15393 19156
rect 15252 19116 15258 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 15381 19119 15439 19125
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15896 19128 15945 19156
rect 15896 19116 15902 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19156 17923 19159
rect 18432 19156 18460 19196
rect 18598 19184 18604 19196
rect 18656 19184 18662 19236
rect 19306 19227 19364 19233
rect 19306 19224 19318 19227
rect 18800 19196 19318 19224
rect 17911 19128 18460 19156
rect 18509 19159 18567 19165
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 18800 19156 18828 19196
rect 19306 19193 19318 19196
rect 19352 19224 19364 19227
rect 19702 19224 19708 19236
rect 19352 19196 19708 19224
rect 19352 19193 19364 19196
rect 19306 19187 19364 19193
rect 19702 19184 19708 19196
rect 19760 19224 19766 19236
rect 20254 19224 20260 19236
rect 19760 19196 20260 19224
rect 19760 19184 19766 19196
rect 20254 19184 20260 19196
rect 20312 19184 20318 19236
rect 18966 19156 18972 19168
rect 18555 19128 18828 19156
rect 18927 19128 18972 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 20438 19156 20444 19168
rect 20399 19128 20444 19156
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 22002 19156 22008 19168
rect 21963 19128 22008 19156
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 23750 19116 23756 19168
rect 23808 19156 23814 19168
rect 24397 19159 24455 19165
rect 24397 19156 24409 19159
rect 23808 19128 24409 19156
rect 23808 19116 23814 19128
rect 24397 19125 24409 19128
rect 24443 19156 24455 19159
rect 25148 19156 25176 19323
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 25869 19295 25927 19301
rect 25869 19261 25881 19295
rect 25915 19292 25927 19295
rect 26510 19292 26516 19304
rect 25915 19264 26516 19292
rect 25915 19261 25927 19264
rect 25869 19255 25927 19261
rect 26510 19252 26516 19264
rect 26568 19292 26574 19304
rect 26697 19295 26755 19301
rect 26697 19292 26709 19295
rect 26568 19264 26709 19292
rect 26568 19252 26574 19264
rect 26697 19261 26709 19264
rect 26743 19261 26755 19295
rect 26697 19255 26755 19261
rect 25314 19156 25320 19168
rect 24443 19128 25320 19156
rect 24443 19125 24455 19128
rect 24397 19119 24455 19125
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 25682 19116 25688 19168
rect 25740 19156 25746 19168
rect 26145 19159 26203 19165
rect 26145 19156 26157 19159
rect 25740 19128 26157 19156
rect 25740 19116 25746 19128
rect 26145 19125 26157 19128
rect 26191 19156 26203 19159
rect 26789 19159 26847 19165
rect 26789 19156 26801 19159
rect 26191 19128 26801 19156
rect 26191 19125 26203 19128
rect 26145 19119 26203 19125
rect 26789 19125 26801 19128
rect 26835 19125 26847 19159
rect 27338 19156 27344 19168
rect 27299 19128 27344 19156
rect 26789 19119 26847 19125
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 3234 18952 3240 18964
rect 1627 18924 3240 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 8754 18952 8760 18964
rect 8715 18924 8760 18952
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 10318 18952 10324 18964
rect 10279 18924 10324 18952
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 11330 18952 11336 18964
rect 11291 18924 11336 18952
rect 11330 18912 11336 18924
rect 11388 18912 11394 18964
rect 11793 18955 11851 18961
rect 11793 18921 11805 18955
rect 11839 18952 11851 18955
rect 12526 18952 12532 18964
rect 11839 18924 12532 18952
rect 11839 18921 11851 18924
rect 11793 18915 11851 18921
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 15470 18952 15476 18964
rect 15431 18924 15476 18952
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 19150 18912 19156 18964
rect 19208 18952 19214 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19208 18924 19809 18952
rect 19208 18912 19214 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 21450 18912 21456 18964
rect 21508 18952 21514 18964
rect 22462 18952 22468 18964
rect 21508 18924 22468 18952
rect 21508 18912 21514 18924
rect 22462 18912 22468 18924
rect 22520 18912 22526 18964
rect 25314 18952 25320 18964
rect 25275 18924 25320 18952
rect 25314 18912 25320 18924
rect 25372 18912 25378 18964
rect 25774 18912 25780 18964
rect 25832 18952 25838 18964
rect 26513 18955 26571 18961
rect 26513 18952 26525 18955
rect 25832 18924 26525 18952
rect 25832 18912 25838 18924
rect 26513 18921 26525 18924
rect 26559 18921 26571 18955
rect 26970 18952 26976 18964
rect 26931 18924 26976 18952
rect 26513 18915 26571 18921
rect 26970 18912 26976 18924
rect 27028 18912 27034 18964
rect 11348 18884 11376 18912
rect 12130 18887 12188 18893
rect 12130 18884 12142 18887
rect 11348 18856 12142 18884
rect 12130 18853 12142 18856
rect 12176 18853 12188 18887
rect 12130 18847 12188 18853
rect 16761 18887 16819 18893
rect 16761 18853 16773 18887
rect 16807 18884 16819 18887
rect 16850 18884 16856 18896
rect 16807 18856 16856 18884
rect 16807 18853 16819 18856
rect 16761 18847 16819 18853
rect 16850 18844 16856 18856
rect 16908 18844 16914 18896
rect 24210 18893 24216 18896
rect 23845 18887 23903 18893
rect 23845 18853 23857 18887
rect 23891 18884 23903 18887
rect 24204 18884 24216 18893
rect 23891 18856 24216 18884
rect 23891 18853 23903 18856
rect 23845 18847 23903 18853
rect 24204 18847 24216 18856
rect 24210 18844 24216 18847
rect 24268 18844 24274 18896
rect 1670 18776 1676 18828
rect 1728 18816 1734 18828
rect 1949 18819 2007 18825
rect 1949 18816 1961 18819
rect 1728 18788 1961 18816
rect 1728 18776 1734 18788
rect 1949 18785 1961 18788
rect 1995 18816 2007 18819
rect 2682 18816 2688 18828
rect 1995 18788 2688 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 3418 18816 3424 18828
rect 2832 18788 3424 18816
rect 2832 18776 2838 18788
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 5258 18816 5264 18828
rect 5219 18788 5264 18816
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5353 18819 5411 18825
rect 5353 18785 5365 18819
rect 5399 18816 5411 18819
rect 6454 18816 6460 18828
rect 5399 18788 6460 18816
rect 5399 18785 5411 18788
rect 5353 18779 5411 18785
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 8570 18816 8576 18828
rect 8483 18788 8576 18816
rect 8570 18776 8576 18788
rect 8628 18816 8634 18828
rect 9030 18816 9036 18828
rect 8628 18788 9036 18816
rect 8628 18776 8634 18788
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 10686 18816 10692 18828
rect 9732 18788 10692 18816
rect 9732 18776 9738 18788
rect 10686 18776 10692 18788
rect 10744 18776 10750 18828
rect 16669 18819 16727 18825
rect 16669 18785 16681 18819
rect 16715 18816 16727 18819
rect 17126 18816 17132 18828
rect 16715 18788 17132 18816
rect 16715 18785 16727 18788
rect 16669 18779 16727 18785
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 17773 18819 17831 18825
rect 17773 18785 17785 18819
rect 17819 18816 17831 18819
rect 18132 18819 18190 18825
rect 18132 18816 18144 18819
rect 17819 18788 18144 18816
rect 17819 18785 17831 18788
rect 17773 18779 17831 18785
rect 18132 18785 18144 18788
rect 18178 18816 18190 18819
rect 19426 18816 19432 18828
rect 18178 18788 19432 18816
rect 18178 18785 18190 18788
rect 18132 18779 18190 18785
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 22002 18776 22008 18828
rect 22060 18816 22066 18828
rect 22373 18819 22431 18825
rect 22373 18816 22385 18819
rect 22060 18788 22385 18816
rect 22060 18776 22066 18788
rect 22373 18785 22385 18788
rect 22419 18785 22431 18819
rect 22373 18779 22431 18785
rect 23937 18819 23995 18825
rect 23937 18785 23949 18819
rect 23983 18816 23995 18819
rect 24670 18816 24676 18828
rect 23983 18788 24676 18816
rect 23983 18785 23995 18788
rect 23937 18779 23995 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 26694 18776 26700 18828
rect 26752 18816 26758 18828
rect 26881 18819 26939 18825
rect 26881 18816 26893 18819
rect 26752 18788 26893 18816
rect 26752 18776 26758 18788
rect 26881 18785 26893 18788
rect 26927 18785 26939 18819
rect 26881 18779 26939 18785
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18717 2099 18751
rect 2041 18711 2099 18717
rect 2056 18680 2084 18711
rect 2130 18708 2136 18760
rect 2188 18748 2194 18760
rect 2593 18751 2651 18757
rect 2593 18748 2605 18751
rect 2188 18720 2605 18748
rect 2188 18708 2194 18720
rect 2593 18717 2605 18720
rect 2639 18717 2651 18751
rect 2593 18711 2651 18717
rect 5166 18708 5172 18760
rect 5224 18748 5230 18760
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 5224 18720 5457 18748
rect 5224 18708 5230 18720
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 5445 18711 5503 18717
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18748 10287 18751
rect 10778 18748 10784 18760
rect 10275 18720 10784 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 10778 18708 10784 18720
rect 10836 18708 10842 18760
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18717 11023 18751
rect 11882 18748 11888 18760
rect 11843 18720 11888 18748
rect 10965 18711 11023 18717
rect 2056 18652 3372 18680
rect 3344 18624 3372 18652
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 10980 18680 11008 18711
rect 11882 18708 11888 18720
rect 11940 18708 11946 18760
rect 16942 18748 16948 18760
rect 16903 18720 16948 18748
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17862 18748 17868 18760
rect 17823 18720 17868 18748
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 20898 18748 20904 18760
rect 20859 18720 20904 18748
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 27157 18751 27215 18757
rect 27157 18717 27169 18751
rect 27203 18748 27215 18751
rect 27338 18748 27344 18760
rect 27203 18720 27344 18748
rect 27203 18717 27215 18720
rect 27157 18711 27215 18717
rect 22005 18683 22063 18689
rect 10652 18652 11560 18680
rect 10652 18640 10658 18652
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 3326 18612 3332 18624
rect 3287 18584 3332 18612
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 3697 18615 3755 18621
rect 3697 18612 3709 18615
rect 3568 18584 3709 18612
rect 3568 18572 3574 18584
rect 3697 18581 3709 18584
rect 3743 18581 3755 18615
rect 3697 18575 3755 18581
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4893 18615 4951 18621
rect 4893 18612 4905 18615
rect 4212 18584 4905 18612
rect 4212 18572 4218 18584
rect 4893 18581 4905 18584
rect 4939 18581 4951 18615
rect 11532 18612 11560 18652
rect 22005 18649 22017 18683
rect 22051 18680 22063 18683
rect 22462 18680 22468 18692
rect 22051 18652 22468 18680
rect 22051 18649 22063 18652
rect 22005 18643 22063 18649
rect 22462 18640 22468 18652
rect 22520 18640 22526 18692
rect 12986 18612 12992 18624
rect 11532 18584 12992 18612
rect 4893 18575 4951 18581
rect 12986 18572 12992 18584
rect 13044 18612 13050 18624
rect 13265 18615 13323 18621
rect 13265 18612 13277 18615
rect 13044 18584 13277 18612
rect 13044 18572 13050 18584
rect 13265 18581 13277 18584
rect 13311 18581 13323 18615
rect 13265 18575 13323 18581
rect 15013 18615 15071 18621
rect 15013 18581 15025 18615
rect 15059 18612 15071 18615
rect 15194 18612 15200 18624
rect 15059 18584 15200 18612
rect 15059 18581 15071 18584
rect 15013 18575 15071 18581
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 16298 18612 16304 18624
rect 16259 18584 16304 18612
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 19245 18615 19303 18621
rect 19245 18612 19257 18615
rect 18656 18584 19257 18612
rect 18656 18572 18662 18584
rect 19245 18581 19257 18584
rect 19291 18581 19303 18615
rect 20254 18612 20260 18624
rect 20215 18584 20260 18612
rect 19245 18575 19303 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 21542 18572 21548 18624
rect 21600 18612 21606 18624
rect 21821 18615 21879 18621
rect 21821 18612 21833 18615
rect 21600 18584 21833 18612
rect 21600 18572 21606 18584
rect 21821 18581 21833 18584
rect 21867 18612 21879 18615
rect 22572 18612 22600 18711
rect 27338 18708 27344 18720
rect 27396 18748 27402 18760
rect 28166 18748 28172 18760
rect 27396 18720 28172 18748
rect 27396 18708 27402 18720
rect 28166 18708 28172 18720
rect 28224 18708 28230 18760
rect 23474 18612 23480 18624
rect 21867 18584 22600 18612
rect 23435 18584 23480 18612
rect 21867 18581 21879 18584
rect 21821 18575 21879 18581
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 3050 18408 3056 18420
rect 3011 18380 3056 18408
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 9490 18368 9496 18420
rect 9548 18408 9554 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 9548 18380 9965 18408
rect 9548 18368 9554 18380
rect 9953 18377 9965 18380
rect 9999 18408 10011 18411
rect 10318 18408 10324 18420
rect 9999 18380 10324 18408
rect 9999 18377 10011 18380
rect 9953 18371 10011 18377
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10594 18408 10600 18420
rect 10555 18380 10600 18408
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 11882 18368 11888 18380
rect 11940 18408 11946 18420
rect 12342 18408 12348 18420
rect 11940 18380 12348 18408
rect 11940 18368 11946 18380
rect 12342 18368 12348 18380
rect 12400 18408 12406 18420
rect 12710 18408 12716 18420
rect 12400 18380 12716 18408
rect 12400 18368 12406 18380
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 16482 18408 16488 18420
rect 16443 18380 16488 18408
rect 16482 18368 16488 18380
rect 16540 18368 16546 18420
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 17770 18408 17776 18420
rect 17000 18380 17776 18408
rect 17000 18368 17006 18380
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 18138 18368 18144 18420
rect 18196 18408 18202 18420
rect 18693 18411 18751 18417
rect 18693 18408 18705 18411
rect 18196 18380 18705 18408
rect 18196 18368 18202 18380
rect 18693 18377 18705 18380
rect 18739 18377 18751 18411
rect 18693 18371 18751 18377
rect 19797 18411 19855 18417
rect 19797 18377 19809 18411
rect 19843 18408 19855 18411
rect 20438 18408 20444 18420
rect 19843 18380 20444 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 1489 18343 1547 18349
rect 1489 18309 1501 18343
rect 1535 18340 1547 18343
rect 3510 18340 3516 18352
rect 1535 18312 3516 18340
rect 1535 18309 1547 18312
rect 1489 18303 1547 18309
rect 3510 18300 3516 18312
rect 3568 18300 3574 18352
rect 4890 18300 4896 18352
rect 4948 18340 4954 18352
rect 5350 18340 5356 18352
rect 4948 18312 5356 18340
rect 4948 18300 4954 18312
rect 5350 18300 5356 18312
rect 5408 18300 5414 18352
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1946 18272 1952 18284
rect 1636 18244 1952 18272
rect 1636 18232 1642 18244
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2130 18272 2136 18284
rect 2091 18244 2136 18272
rect 2130 18232 2136 18244
rect 2188 18232 2194 18284
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18272 4215 18275
rect 5074 18272 5080 18284
rect 4203 18244 5080 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 1670 18164 1676 18216
rect 1728 18204 1734 18216
rect 1857 18207 1915 18213
rect 1857 18204 1869 18207
rect 1728 18176 1869 18204
rect 1728 18164 1734 18176
rect 1857 18173 1869 18176
rect 1903 18204 1915 18207
rect 2958 18204 2964 18216
rect 1903 18176 2964 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 2958 18164 2964 18176
rect 3016 18164 3022 18216
rect 3234 18164 3240 18216
rect 3292 18204 3298 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3292 18176 3433 18204
rect 3292 18164 3298 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3620 18204 3648 18235
rect 5074 18232 5080 18244
rect 5132 18272 5138 18284
rect 5537 18275 5595 18281
rect 5537 18272 5549 18275
rect 5132 18244 5549 18272
rect 5132 18232 5138 18244
rect 5537 18241 5549 18244
rect 5583 18241 5595 18275
rect 5537 18235 5595 18241
rect 11241 18275 11299 18281
rect 11241 18241 11253 18275
rect 11287 18272 11299 18275
rect 19150 18272 19156 18284
rect 11287 18244 12572 18272
rect 19111 18244 19156 18272
rect 11287 18241 11299 18244
rect 11241 18235 11299 18241
rect 12544 18216 12572 18244
rect 19150 18232 19156 18244
rect 19208 18232 19214 18284
rect 19337 18275 19395 18281
rect 19337 18241 19349 18275
rect 19383 18272 19395 18275
rect 19426 18272 19432 18284
rect 19383 18244 19432 18272
rect 19383 18241 19395 18244
rect 19337 18235 19395 18241
rect 19426 18232 19432 18244
rect 19484 18272 19490 18284
rect 19812 18272 19840 18371
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 21450 18408 21456 18420
rect 21411 18380 21456 18408
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 23106 18408 23112 18420
rect 23067 18380 23112 18408
rect 23106 18368 23112 18380
rect 23164 18368 23170 18420
rect 26418 18368 26424 18420
rect 26476 18408 26482 18420
rect 26881 18411 26939 18417
rect 26881 18408 26893 18411
rect 26476 18380 26893 18408
rect 26476 18368 26482 18380
rect 26881 18377 26893 18380
rect 26927 18377 26939 18411
rect 26881 18371 26939 18377
rect 26970 18368 26976 18420
rect 27028 18408 27034 18420
rect 27801 18411 27859 18417
rect 27801 18408 27813 18411
rect 27028 18380 27813 18408
rect 27028 18368 27034 18380
rect 27801 18377 27813 18380
rect 27847 18377 27859 18411
rect 27801 18371 27859 18377
rect 24946 18300 24952 18352
rect 25004 18340 25010 18352
rect 25406 18340 25412 18352
rect 25004 18312 25412 18340
rect 25004 18300 25010 18312
rect 25406 18300 25412 18312
rect 25464 18300 25470 18352
rect 19484 18244 19840 18272
rect 19484 18232 19490 18244
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20312 18244 20821 18272
rect 20312 18232 20318 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 21542 18232 21548 18284
rect 21600 18272 21606 18284
rect 22557 18275 22615 18281
rect 22557 18272 22569 18275
rect 21600 18244 22569 18272
rect 21600 18232 21606 18244
rect 22557 18241 22569 18244
rect 22603 18241 22615 18275
rect 22557 18235 22615 18241
rect 23474 18232 23480 18284
rect 23532 18272 23538 18284
rect 24489 18275 24547 18281
rect 24489 18272 24501 18275
rect 23532 18244 24501 18272
rect 23532 18232 23538 18244
rect 24489 18241 24501 18244
rect 24535 18272 24547 18275
rect 24762 18272 24768 18284
rect 24535 18244 24768 18272
rect 24535 18241 24547 18244
rect 24489 18235 24547 18241
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 3421 18167 3479 18173
rect 3528 18176 3648 18204
rect 4525 18207 4583 18213
rect 3528 18136 3556 18176
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4890 18204 4896 18216
rect 4571 18176 4896 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 5166 18164 5172 18216
rect 5224 18204 5230 18216
rect 5997 18207 6055 18213
rect 5997 18204 6009 18207
rect 5224 18176 6009 18204
rect 5224 18164 5230 18176
rect 5997 18173 6009 18176
rect 6043 18173 6055 18207
rect 5997 18167 6055 18173
rect 8478 18164 8484 18216
rect 8536 18204 8542 18216
rect 8573 18207 8631 18213
rect 8573 18204 8585 18207
rect 8536 18176 8585 18204
rect 8536 18164 8542 18176
rect 8573 18173 8585 18176
rect 8619 18173 8631 18207
rect 8573 18167 8631 18173
rect 12342 18164 12348 18216
rect 12400 18204 12406 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12400 18176 12449 18204
rect 12400 18164 12406 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 15010 18204 15016 18216
rect 12584 18176 12677 18204
rect 14971 18176 15016 18204
rect 12584 18164 12590 18176
rect 15010 18164 15016 18176
rect 15068 18204 15074 18216
rect 15105 18207 15163 18213
rect 15105 18204 15117 18207
rect 15068 18176 15117 18204
rect 15068 18164 15074 18176
rect 15105 18173 15117 18176
rect 15151 18173 15163 18207
rect 15105 18167 15163 18173
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18204 20223 18207
rect 20211 18176 20300 18204
rect 20211 18173 20223 18176
rect 20165 18167 20223 18173
rect 5350 18136 5356 18148
rect 2884 18108 3556 18136
rect 4816 18108 5212 18136
rect 5311 18108 5356 18136
rect 2884 18080 2912 18108
rect 1854 18028 1860 18080
rect 1912 18068 1918 18080
rect 2501 18071 2559 18077
rect 2501 18068 2513 18071
rect 1912 18040 2513 18068
rect 1912 18028 1918 18040
rect 2501 18037 2513 18040
rect 2547 18037 2559 18071
rect 2866 18068 2872 18080
rect 2827 18040 2872 18068
rect 2501 18031 2559 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 3510 18068 3516 18080
rect 3471 18040 3516 18068
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4816 18077 4844 18108
rect 4801 18071 4859 18077
rect 4801 18068 4813 18071
rect 4304 18040 4813 18068
rect 4304 18028 4310 18040
rect 4801 18037 4813 18040
rect 4847 18037 4859 18071
rect 4982 18068 4988 18080
rect 4943 18040 4988 18068
rect 4801 18031 4859 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 5184 18068 5212 18108
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 8818 18139 8876 18145
rect 8818 18136 8830 18139
rect 7668 18108 8830 18136
rect 7668 18080 7696 18108
rect 8818 18105 8830 18108
rect 8864 18105 8876 18139
rect 12544 18136 12572 18164
rect 12704 18139 12762 18145
rect 12704 18136 12716 18139
rect 12544 18108 12716 18136
rect 8818 18099 8876 18105
rect 12704 18105 12716 18108
rect 12750 18136 12762 18139
rect 13906 18136 13912 18148
rect 12750 18108 13912 18136
rect 12750 18105 12762 18108
rect 12704 18099 12762 18105
rect 13906 18096 13912 18108
rect 13964 18136 13970 18148
rect 14274 18136 14280 18148
rect 13964 18108 14280 18136
rect 13964 18096 13970 18108
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 14645 18139 14703 18145
rect 14645 18105 14657 18139
rect 14691 18136 14703 18139
rect 15372 18139 15430 18145
rect 15372 18136 15384 18139
rect 14691 18108 15384 18136
rect 14691 18105 14703 18108
rect 14645 18099 14703 18105
rect 15372 18105 15384 18108
rect 15418 18136 15430 18139
rect 15838 18136 15844 18148
rect 15418 18108 15844 18136
rect 15418 18105 15430 18108
rect 15372 18099 15430 18105
rect 15838 18096 15844 18108
rect 15896 18096 15902 18148
rect 19061 18139 19119 18145
rect 19061 18105 19073 18139
rect 19107 18136 19119 18139
rect 20272 18136 20300 18176
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 20404 18176 20637 18204
rect 20404 18164 20410 18176
rect 20625 18173 20637 18176
rect 20671 18204 20683 18207
rect 20898 18204 20904 18216
rect 20671 18176 20904 18204
rect 20671 18173 20683 18176
rect 20625 18167 20683 18173
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 22002 18164 22008 18216
rect 22060 18164 22066 18216
rect 22465 18207 22523 18213
rect 22465 18173 22477 18207
rect 22511 18204 22523 18207
rect 23106 18204 23112 18216
rect 22511 18176 23112 18204
rect 22511 18173 22523 18176
rect 22465 18167 22523 18173
rect 23106 18164 23112 18176
rect 23164 18164 23170 18216
rect 25501 18207 25559 18213
rect 25501 18204 25513 18207
rect 25332 18176 25513 18204
rect 20530 18136 20536 18148
rect 19107 18108 20208 18136
rect 20272 18108 20536 18136
rect 19107 18105 19119 18108
rect 19061 18099 19119 18105
rect 20180 18080 20208 18108
rect 20530 18096 20536 18108
rect 20588 18136 20594 18148
rect 20717 18139 20775 18145
rect 20717 18136 20729 18139
rect 20588 18108 20729 18136
rect 20588 18096 20594 18108
rect 20717 18105 20729 18108
rect 20763 18105 20775 18139
rect 20717 18099 20775 18105
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 21821 18139 21879 18145
rect 21821 18136 21833 18139
rect 20864 18108 21833 18136
rect 20864 18096 20870 18108
rect 21821 18105 21833 18108
rect 21867 18136 21879 18139
rect 22020 18136 22048 18164
rect 22646 18136 22652 18148
rect 21867 18108 22652 18136
rect 21867 18105 21879 18108
rect 21821 18099 21879 18105
rect 22646 18096 22652 18108
rect 22704 18096 22710 18148
rect 22738 18096 22744 18148
rect 22796 18136 22802 18148
rect 23477 18139 23535 18145
rect 23477 18136 23489 18139
rect 22796 18108 23489 18136
rect 22796 18096 22802 18108
rect 23477 18105 23489 18108
rect 23523 18136 23535 18139
rect 24397 18139 24455 18145
rect 24397 18136 24409 18139
rect 23523 18108 24409 18136
rect 23523 18105 23535 18108
rect 23477 18099 23535 18105
rect 24397 18105 24409 18108
rect 24443 18105 24455 18139
rect 24397 18099 24455 18105
rect 5445 18071 5503 18077
rect 5445 18068 5457 18071
rect 5184 18040 5457 18068
rect 5445 18037 5457 18040
rect 5491 18037 5503 18071
rect 6454 18068 6460 18080
rect 6415 18040 6460 18068
rect 5445 18031 5503 18037
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 7650 18068 7656 18080
rect 7611 18040 7656 18068
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 8110 18068 8116 18080
rect 8071 18040 8116 18068
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 8478 18068 8484 18080
rect 8439 18040 8484 18068
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 11333 18071 11391 18077
rect 11333 18037 11345 18071
rect 11379 18068 11391 18071
rect 12802 18068 12808 18080
rect 11379 18040 12808 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 16942 18028 16948 18080
rect 17000 18068 17006 18080
rect 17037 18071 17095 18077
rect 17037 18068 17049 18071
rect 17000 18040 17049 18068
rect 17000 18028 17006 18040
rect 17037 18037 17049 18040
rect 17083 18037 17095 18071
rect 17037 18031 17095 18037
rect 17126 18028 17132 18080
rect 17184 18068 17190 18080
rect 17405 18071 17463 18077
rect 17405 18068 17417 18071
rect 17184 18040 17417 18068
rect 17184 18028 17190 18040
rect 17405 18037 17417 18040
rect 17451 18037 17463 18071
rect 17405 18031 17463 18037
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18325 18071 18383 18077
rect 18325 18068 18337 18071
rect 17920 18040 18337 18068
rect 17920 18028 17926 18040
rect 18325 18037 18337 18040
rect 18371 18068 18383 18071
rect 18966 18068 18972 18080
rect 18371 18040 18972 18068
rect 18371 18037 18383 18040
rect 18325 18031 18383 18037
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20257 18071 20315 18077
rect 20257 18068 20269 18071
rect 20220 18040 20269 18068
rect 20220 18028 20226 18040
rect 20257 18037 20269 18040
rect 20303 18037 20315 18071
rect 20257 18031 20315 18037
rect 21910 18028 21916 18080
rect 21968 18068 21974 18080
rect 22005 18071 22063 18077
rect 22005 18068 22017 18071
rect 21968 18040 22017 18068
rect 21968 18028 21974 18040
rect 22005 18037 22017 18040
rect 22051 18037 22063 18071
rect 22005 18031 22063 18037
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22373 18071 22431 18077
rect 22373 18068 22385 18071
rect 22152 18040 22385 18068
rect 22152 18028 22158 18040
rect 22373 18037 22385 18040
rect 22419 18037 22431 18071
rect 23934 18068 23940 18080
rect 23895 18040 23940 18068
rect 22373 18031 22431 18037
rect 23934 18028 23940 18040
rect 23992 18028 23998 18080
rect 24026 18028 24032 18080
rect 24084 18068 24090 18080
rect 24305 18071 24363 18077
rect 24305 18068 24317 18071
rect 24084 18040 24317 18068
rect 24084 18028 24090 18040
rect 24305 18037 24317 18040
rect 24351 18037 24363 18071
rect 24305 18031 24363 18037
rect 24670 18028 24676 18080
rect 24728 18068 24734 18080
rect 25332 18077 25360 18176
rect 25501 18173 25513 18176
rect 25547 18173 25559 18207
rect 25501 18167 25559 18173
rect 25406 18096 25412 18148
rect 25464 18136 25470 18148
rect 25746 18139 25804 18145
rect 25746 18136 25758 18139
rect 25464 18108 25758 18136
rect 25464 18096 25470 18108
rect 25746 18105 25758 18108
rect 25792 18105 25804 18139
rect 25746 18099 25804 18105
rect 26694 18096 26700 18148
rect 26752 18136 26758 18148
rect 27433 18139 27491 18145
rect 27433 18136 27445 18139
rect 26752 18108 27445 18136
rect 26752 18096 26758 18108
rect 27433 18105 27445 18108
rect 27479 18105 27491 18139
rect 27433 18099 27491 18105
rect 24949 18071 25007 18077
rect 24949 18068 24961 18071
rect 24728 18040 24961 18068
rect 24728 18028 24734 18040
rect 24949 18037 24961 18040
rect 24995 18068 25007 18071
rect 25317 18071 25375 18077
rect 25317 18068 25329 18071
rect 24995 18040 25329 18068
rect 24995 18037 25007 18040
rect 24949 18031 25007 18037
rect 25317 18037 25329 18040
rect 25363 18037 25375 18071
rect 28166 18068 28172 18080
rect 28127 18040 28172 18068
rect 25317 18031 25375 18037
rect 28166 18028 28172 18040
rect 28224 18028 28230 18080
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2866 17824 2872 17836
rect 2924 17864 2930 17876
rect 4249 17867 4307 17873
rect 4249 17864 4261 17867
rect 2924 17836 4261 17864
rect 2924 17824 2930 17836
rect 4249 17833 4261 17836
rect 4295 17864 4307 17867
rect 4338 17864 4344 17876
rect 4295 17836 4344 17864
rect 4295 17833 4307 17836
rect 4249 17827 4307 17833
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 4893 17867 4951 17873
rect 4893 17833 4905 17867
rect 4939 17864 4951 17867
rect 5258 17864 5264 17876
rect 4939 17836 5264 17864
rect 4939 17833 4951 17836
rect 4893 17827 4951 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 9030 17864 9036 17876
rect 8991 17836 9036 17864
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 9493 17867 9551 17873
rect 9493 17833 9505 17867
rect 9539 17864 9551 17867
rect 9674 17864 9680 17876
rect 9539 17836 9680 17864
rect 9539 17833 9551 17836
rect 9493 17827 9551 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 10778 17824 10784 17876
rect 10836 17864 10842 17876
rect 11701 17867 11759 17873
rect 11701 17864 11713 17867
rect 10836 17836 11713 17864
rect 10836 17824 10842 17836
rect 11701 17833 11713 17836
rect 11747 17833 11759 17867
rect 11701 17827 11759 17833
rect 11974 17824 11980 17876
rect 12032 17864 12038 17876
rect 12069 17867 12127 17873
rect 12069 17864 12081 17867
rect 12032 17836 12081 17864
rect 12032 17824 12038 17836
rect 12069 17833 12081 17836
rect 12115 17833 12127 17867
rect 12069 17827 12127 17833
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 12492 17836 13277 17864
rect 12492 17824 12498 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13630 17864 13636 17876
rect 13591 17836 13636 17864
rect 13265 17827 13323 17833
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 14921 17867 14979 17873
rect 14921 17833 14933 17867
rect 14967 17864 14979 17867
rect 15102 17864 15108 17876
rect 14967 17836 15108 17864
rect 14967 17833 14979 17836
rect 14921 17827 14979 17833
rect 15102 17824 15108 17836
rect 15160 17864 15166 17876
rect 15562 17864 15568 17876
rect 15160 17836 15568 17864
rect 15160 17824 15166 17836
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 17770 17864 17776 17876
rect 17731 17836 17776 17864
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18138 17864 18144 17876
rect 18012 17836 18144 17864
rect 18012 17824 18018 17836
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 18230 17824 18236 17876
rect 18288 17864 18294 17876
rect 18877 17867 18935 17873
rect 18877 17864 18889 17867
rect 18288 17836 18889 17864
rect 18288 17824 18294 17836
rect 18877 17833 18889 17836
rect 18923 17833 18935 17867
rect 18877 17827 18935 17833
rect 19981 17867 20039 17873
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20162 17864 20168 17876
rect 20027 17836 20168 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 20346 17864 20352 17876
rect 20307 17836 20352 17864
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 21085 17867 21143 17873
rect 21085 17833 21097 17867
rect 21131 17864 21143 17867
rect 22002 17864 22008 17876
rect 21131 17836 22008 17864
rect 21131 17833 21143 17836
rect 21085 17827 21143 17833
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 1756 17799 1814 17805
rect 1756 17765 1768 17799
rect 1802 17796 1814 17799
rect 2038 17796 2044 17808
rect 1802 17768 2044 17796
rect 1802 17765 1814 17768
rect 1756 17759 1814 17765
rect 2038 17756 2044 17768
rect 2096 17796 2102 17808
rect 2958 17796 2964 17808
rect 2096 17768 2964 17796
rect 2096 17756 2102 17768
rect 2958 17756 2964 17768
rect 3016 17796 3022 17808
rect 3421 17799 3479 17805
rect 3421 17796 3433 17799
rect 3016 17768 3433 17796
rect 3016 17756 3022 17768
rect 3421 17765 3433 17768
rect 3467 17765 3479 17799
rect 3421 17759 3479 17765
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 10686 17796 10692 17808
rect 9456 17768 10692 17796
rect 9456 17756 9462 17768
rect 10686 17756 10692 17768
rect 10744 17756 10750 17808
rect 11330 17756 11336 17808
rect 11388 17796 11394 17808
rect 11517 17799 11575 17805
rect 11517 17796 11529 17799
rect 11388 17768 11529 17796
rect 11388 17756 11394 17768
rect 11517 17765 11529 17768
rect 11563 17796 11575 17799
rect 13814 17796 13820 17808
rect 11563 17768 13820 17796
rect 11563 17765 11575 17768
rect 11517 17759 11575 17765
rect 5074 17688 5080 17740
rect 5132 17728 5138 17740
rect 5241 17731 5299 17737
rect 5241 17728 5253 17731
rect 5132 17700 5253 17728
rect 5132 17688 5138 17700
rect 5241 17697 5253 17700
rect 5287 17697 5299 17731
rect 8386 17728 8392 17740
rect 8347 17700 8392 17728
rect 5241 17691 5299 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 10042 17728 10048 17740
rect 10003 17700 10048 17728
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 1486 17660 1492 17672
rect 1447 17632 1492 17660
rect 1486 17620 1492 17632
rect 1544 17620 1550 17672
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 4985 17663 5043 17669
rect 4985 17660 4997 17663
rect 3936 17632 4997 17660
rect 3936 17620 3942 17632
rect 4985 17629 4997 17632
rect 5031 17629 5043 17663
rect 4985 17623 5043 17629
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 8481 17663 8539 17669
rect 8481 17660 8493 17663
rect 7800 17632 8493 17660
rect 7800 17620 7806 17632
rect 8481 17629 8493 17632
rect 8527 17629 8539 17663
rect 8481 17623 8539 17629
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 8628 17632 8673 17660
rect 8628 17620 8634 17632
rect 9858 17620 9864 17672
rect 9916 17660 9922 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 9916 17632 10149 17660
rect 9916 17620 9922 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10226 17620 10232 17672
rect 10284 17660 10290 17672
rect 12158 17660 12164 17672
rect 10284 17632 10329 17660
rect 12119 17632 12164 17660
rect 10284 17620 10290 17632
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 12360 17669 12388 17768
rect 13814 17756 13820 17768
rect 13872 17756 13878 17808
rect 16574 17756 16580 17808
rect 16632 17805 16638 17808
rect 16632 17799 16696 17805
rect 16632 17765 16650 17799
rect 16684 17765 16696 17799
rect 17788 17796 17816 17824
rect 18601 17799 18659 17805
rect 18601 17796 18613 17799
rect 17788 17768 18613 17796
rect 16632 17759 16696 17765
rect 18601 17765 18613 17768
rect 18647 17796 18659 17799
rect 18782 17796 18788 17808
rect 18647 17768 18788 17796
rect 18647 17765 18659 17768
rect 18601 17759 18659 17765
rect 16632 17756 16638 17759
rect 18782 17756 18788 17768
rect 18840 17756 18846 17808
rect 24765 17799 24823 17805
rect 24765 17765 24777 17799
rect 24811 17796 24823 17799
rect 25225 17799 25283 17805
rect 25225 17796 25237 17799
rect 24811 17768 25237 17796
rect 24811 17765 24823 17768
rect 24765 17759 24823 17765
rect 25225 17765 25237 17768
rect 25271 17796 25283 17799
rect 25682 17796 25688 17808
rect 25271 17768 25688 17796
rect 25271 17765 25283 17768
rect 25225 17759 25283 17765
rect 25682 17756 25688 17768
rect 25740 17756 25746 17808
rect 13725 17731 13783 17737
rect 13725 17697 13737 17731
rect 13771 17728 13783 17731
rect 14366 17728 14372 17740
rect 13771 17700 14372 17728
rect 13771 17697 13783 17700
rect 13725 17691 13783 17697
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 15010 17688 15016 17740
rect 15068 17728 15074 17740
rect 15068 17700 16436 17728
rect 15068 17688 15074 17700
rect 16408 17672 16436 17700
rect 18506 17688 18512 17740
rect 18564 17728 18570 17740
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 18564 17700 19257 17728
rect 18564 17688 18570 17700
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 21358 17688 21364 17740
rect 21416 17728 21422 17740
rect 22370 17737 22376 17740
rect 22364 17728 22376 17737
rect 21416 17700 22376 17728
rect 21416 17688 21422 17700
rect 22364 17691 22376 17700
rect 22370 17688 22376 17691
rect 22428 17688 22434 17740
rect 25317 17731 25375 17737
rect 25317 17697 25329 17731
rect 25363 17728 25375 17731
rect 25774 17728 25780 17740
rect 25363 17700 25780 17728
rect 25363 17697 25375 17700
rect 25317 17691 25375 17697
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 26418 17688 26424 17740
rect 26476 17728 26482 17740
rect 26881 17731 26939 17737
rect 26881 17728 26893 17731
rect 26476 17700 26893 17728
rect 26476 17688 26482 17700
rect 26881 17697 26893 17700
rect 26927 17697 26939 17731
rect 26881 17691 26939 17697
rect 26973 17731 27031 17737
rect 26973 17697 26985 17731
rect 27019 17728 27031 17731
rect 27798 17728 27804 17740
rect 27019 17700 27804 17728
rect 27019 17697 27031 17700
rect 26973 17691 27031 17697
rect 27798 17688 27804 17700
rect 27856 17688 27862 17740
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 13909 17663 13967 17669
rect 13909 17629 13921 17663
rect 13955 17660 13967 17663
rect 14274 17660 14280 17672
rect 13955 17632 14280 17660
rect 13955 17629 13967 17632
rect 13909 17623 13967 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 16298 17660 16304 17672
rect 15335 17632 16304 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 16298 17620 16304 17632
rect 16356 17620 16362 17672
rect 16390 17620 16396 17672
rect 16448 17660 16454 17672
rect 16448 17632 16493 17660
rect 16448 17620 16454 17632
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 19337 17663 19395 17669
rect 19337 17660 19349 17663
rect 18472 17632 19349 17660
rect 18472 17620 18478 17632
rect 19337 17629 19349 17632
rect 19383 17629 19395 17663
rect 19337 17623 19395 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 2740 17564 3801 17592
rect 2740 17552 2746 17564
rect 3789 17561 3801 17564
rect 3835 17561 3847 17595
rect 3789 17555 3847 17561
rect 8021 17595 8079 17601
rect 8021 17561 8033 17595
rect 8067 17592 8079 17595
rect 10962 17592 10968 17604
rect 8067 17564 10968 17592
rect 8067 17561 8079 17564
rect 8021 17555 8079 17561
rect 10962 17552 10968 17564
rect 11020 17592 11026 17604
rect 11057 17595 11115 17601
rect 11057 17592 11069 17595
rect 11020 17564 11069 17592
rect 11020 17552 11026 17564
rect 11057 17561 11069 17564
rect 11103 17561 11115 17595
rect 19352 17592 19380 17623
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 22097 17663 22155 17669
rect 19484 17632 19529 17660
rect 19484 17620 19490 17632
rect 22097 17629 22109 17663
rect 22143 17629 22155 17663
rect 25498 17660 25504 17672
rect 25459 17632 25504 17660
rect 22097 17623 22155 17629
rect 20438 17592 20444 17604
rect 19352 17564 20444 17592
rect 11057 17555 11115 17561
rect 20438 17552 20444 17564
rect 20496 17552 20502 17604
rect 6362 17524 6368 17536
rect 6323 17496 6368 17524
rect 6362 17484 6368 17496
rect 6420 17484 6426 17536
rect 6914 17524 6920 17536
rect 6875 17496 6920 17524
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 7929 17527 7987 17533
rect 7929 17493 7941 17527
rect 7975 17524 7987 17527
rect 8110 17524 8116 17536
rect 7975 17496 8116 17524
rect 7975 17493 7987 17496
rect 7929 17487 7987 17493
rect 8110 17484 8116 17496
rect 8168 17524 8174 17536
rect 8570 17524 8576 17536
rect 8168 17496 8576 17524
rect 8168 17484 8174 17496
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 9677 17527 9735 17533
rect 9677 17493 9689 17527
rect 9723 17524 9735 17527
rect 10410 17524 10416 17536
rect 9723 17496 10416 17524
rect 9723 17493 9735 17496
rect 9677 17487 9735 17493
rect 10410 17484 10416 17496
rect 10468 17484 10474 17536
rect 12802 17524 12808 17536
rect 12763 17496 12808 17524
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 13078 17524 13084 17536
rect 13039 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 21542 17524 21548 17536
rect 21503 17496 21548 17524
rect 21542 17484 21548 17496
rect 21600 17484 21606 17536
rect 22112 17524 22140 17623
rect 25498 17620 25504 17632
rect 25556 17620 25562 17672
rect 27157 17663 27215 17669
rect 27157 17629 27169 17663
rect 27203 17660 27215 17663
rect 27430 17660 27436 17672
rect 27203 17632 27436 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 27430 17620 27436 17632
rect 27488 17620 27494 17672
rect 23477 17595 23535 17601
rect 23477 17561 23489 17595
rect 23523 17592 23535 17595
rect 24118 17592 24124 17604
rect 23523 17564 24124 17592
rect 23523 17561 23535 17564
rect 23477 17555 23535 17561
rect 24118 17552 24124 17564
rect 24176 17552 24182 17604
rect 25590 17552 25596 17604
rect 25648 17592 25654 17604
rect 26513 17595 26571 17601
rect 26513 17592 26525 17595
rect 25648 17564 26525 17592
rect 25648 17552 25654 17564
rect 26513 17561 26525 17564
rect 26559 17561 26571 17595
rect 26513 17555 26571 17561
rect 22278 17524 22284 17536
rect 22112 17496 22284 17524
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 24026 17524 24032 17536
rect 23987 17496 24032 17524
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 24857 17527 24915 17533
rect 24857 17493 24869 17527
rect 24903 17524 24915 17527
rect 25222 17524 25228 17536
rect 24903 17496 25228 17524
rect 24903 17493 24915 17496
rect 24857 17487 24915 17493
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 25406 17484 25412 17536
rect 25464 17524 25470 17536
rect 25869 17527 25927 17533
rect 25869 17524 25881 17527
rect 25464 17496 25881 17524
rect 25464 17484 25470 17496
rect 25869 17493 25881 17496
rect 25915 17493 25927 17527
rect 26326 17524 26332 17536
rect 26287 17496 26332 17524
rect 25869 17487 25927 17493
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 2958 17320 2964 17332
rect 2919 17292 2964 17320
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5132 17292 5457 17320
rect 5132 17280 5138 17292
rect 5445 17289 5457 17292
rect 5491 17320 5503 17323
rect 5534 17320 5540 17332
rect 5491 17292 5540 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 7926 17320 7932 17332
rect 7839 17292 7932 17320
rect 7926 17280 7932 17292
rect 7984 17320 7990 17332
rect 8386 17320 8392 17332
rect 7984 17292 8392 17320
rect 7984 17280 7990 17292
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 9824 17292 10517 17320
rect 9824 17280 9830 17292
rect 10505 17289 10517 17292
rect 10551 17289 10563 17323
rect 10505 17283 10563 17289
rect 13538 17280 13544 17332
rect 13596 17320 13602 17332
rect 13909 17323 13967 17329
rect 13909 17320 13921 17323
rect 13596 17292 13921 17320
rect 13596 17280 13602 17292
rect 13909 17289 13921 17292
rect 13955 17320 13967 17323
rect 14366 17320 14372 17332
rect 13955 17292 14372 17320
rect 13955 17289 13967 17292
rect 13909 17283 13967 17289
rect 14366 17280 14372 17292
rect 14424 17280 14430 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 15010 17320 15016 17332
rect 14783 17292 15016 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 10686 17212 10692 17264
rect 10744 17252 10750 17264
rect 10744 17224 11100 17252
rect 10744 17212 10750 17224
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 1581 17187 1639 17193
rect 1581 17184 1593 17187
rect 1544 17156 1593 17184
rect 1544 17144 1550 17156
rect 1581 17153 1593 17156
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 10962 17184 10968 17196
rect 7055 17156 8156 17184
rect 10923 17156 10968 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 1854 17125 1860 17128
rect 1848 17116 1860 17125
rect 1815 17088 1860 17116
rect 1848 17079 1860 17088
rect 1912 17116 1918 17128
rect 2314 17116 2320 17128
rect 1912 17088 2320 17116
rect 1854 17076 1860 17079
rect 1912 17076 1918 17088
rect 2314 17076 2320 17088
rect 2372 17076 2378 17128
rect 3878 17116 3884 17128
rect 3791 17088 3884 17116
rect 3878 17076 3884 17088
rect 3936 17116 3942 17128
rect 4338 17125 4344 17128
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 3936 17088 4077 17116
rect 3936 17076 3942 17088
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 4332 17116 4344 17125
rect 4299 17088 4344 17116
rect 4065 17079 4123 17085
rect 4332 17079 4344 17088
rect 4338 17076 4344 17079
rect 4396 17076 4402 17128
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7984 17088 8033 17116
rect 7984 17076 7990 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8128 17116 8156 17156
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 11072 17193 11100 17224
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 14844 17252 14872 17292
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16632 17292 17141 17320
rect 16632 17280 16638 17292
rect 17129 17289 17141 17292
rect 17175 17289 17187 17323
rect 20438 17320 20444 17332
rect 20399 17292 20444 17320
rect 17129 17283 17187 17289
rect 20438 17280 20444 17292
rect 20496 17280 20502 17332
rect 21358 17320 21364 17332
rect 21319 17292 21364 17320
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 21818 17320 21824 17332
rect 21779 17292 21824 17320
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 24670 17320 24676 17332
rect 24044 17292 24676 17320
rect 12860 17224 14872 17252
rect 12860 17212 12866 17224
rect 11057 17187 11115 17193
rect 11057 17153 11069 17187
rect 11103 17153 11115 17187
rect 13078 17184 13084 17196
rect 13039 17156 13084 17184
rect 11057 17147 11115 17153
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 13630 17184 13636 17196
rect 13587 17156 13636 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 14844 17193 14872 17224
rect 17865 17255 17923 17261
rect 17865 17221 17877 17255
rect 17911 17252 17923 17255
rect 18506 17252 18512 17264
rect 17911 17224 18512 17252
rect 17911 17221 17923 17224
rect 17865 17215 17923 17221
rect 18506 17212 18512 17224
rect 18564 17212 18570 17264
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 22833 17255 22891 17261
rect 22833 17252 22845 17255
rect 22336 17224 22845 17252
rect 22336 17212 22342 17224
rect 22833 17221 22845 17224
rect 22879 17252 22891 17255
rect 23845 17255 23903 17261
rect 23845 17252 23857 17255
rect 22879 17224 23857 17252
rect 22879 17221 22891 17224
rect 22833 17215 22891 17221
rect 23845 17221 23857 17224
rect 23891 17252 23903 17255
rect 24044 17252 24072 17292
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 25314 17280 25320 17332
rect 25372 17320 25378 17332
rect 25961 17323 26019 17329
rect 25961 17320 25973 17323
rect 25372 17292 25973 17320
rect 25372 17280 25378 17292
rect 25961 17289 25973 17292
rect 26007 17320 26019 17323
rect 26237 17323 26295 17329
rect 26237 17320 26249 17323
rect 26007 17292 26249 17320
rect 26007 17289 26019 17292
rect 25961 17283 26019 17289
rect 26237 17289 26249 17292
rect 26283 17289 26295 17323
rect 26510 17320 26516 17332
rect 26471 17292 26516 17320
rect 26237 17283 26295 17289
rect 26510 17280 26516 17292
rect 26568 17280 26574 17332
rect 23891 17224 24072 17252
rect 23891 17221 23903 17224
rect 23845 17215 23903 17221
rect 24044 17193 24072 17224
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 21729 17187 21787 17193
rect 21729 17153 21741 17187
rect 21775 17184 21787 17187
rect 22465 17187 22523 17193
rect 22465 17184 22477 17187
rect 21775 17156 22477 17184
rect 21775 17153 21787 17156
rect 21729 17147 21787 17153
rect 22465 17153 22477 17156
rect 22511 17153 22523 17187
rect 22465 17147 22523 17153
rect 24029 17187 24087 17193
rect 24029 17153 24041 17187
rect 24075 17153 24087 17187
rect 24029 17147 24087 17153
rect 10042 17116 10048 17128
rect 8128 17088 10048 17116
rect 8021 17079 8079 17085
rect 10042 17076 10048 17088
rect 10100 17116 10106 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 10100 17088 10333 17116
rect 10100 17076 10106 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10321 17079 10379 17085
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 15102 17125 15108 17128
rect 15096 17116 15108 17125
rect 12124 17088 12940 17116
rect 15063 17088 15108 17116
rect 12124 17076 12130 17088
rect 3510 16980 3516 16992
rect 3471 16952 3516 16980
rect 3510 16940 3516 16952
rect 3568 16980 3574 16992
rect 3896 16989 3924 17076
rect 6638 17008 6644 17060
rect 6696 17048 6702 17060
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 6696 17020 7481 17048
rect 6696 17008 6702 17020
rect 7469 17017 7481 17020
rect 7515 17048 7527 17051
rect 7742 17048 7748 17060
rect 7515 17020 7748 17048
rect 7515 17017 7527 17020
rect 7469 17011 7527 17017
rect 7742 17008 7748 17020
rect 7800 17008 7806 17060
rect 8288 17051 8346 17057
rect 8288 17017 8300 17051
rect 8334 17048 8346 17051
rect 8570 17048 8576 17060
rect 8334 17020 8576 17048
rect 8334 17017 8346 17020
rect 8288 17011 8346 17017
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 10410 17008 10416 17060
rect 10468 17048 10474 17060
rect 10873 17051 10931 17057
rect 10873 17048 10885 17051
rect 10468 17020 10885 17048
rect 10468 17008 10474 17020
rect 10873 17017 10885 17020
rect 10919 17017 10931 17051
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 10873 17011 10931 17017
rect 11808 17020 12817 17048
rect 3881 16983 3939 16989
rect 3881 16980 3893 16983
rect 3568 16952 3893 16980
rect 3568 16940 3574 16952
rect 3881 16949 3893 16952
rect 3927 16980 3939 16983
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 3927 16952 6009 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 5997 16949 6009 16952
rect 6043 16949 6055 16983
rect 5997 16943 6055 16949
rect 6549 16983 6607 16989
rect 6549 16949 6561 16983
rect 6595 16980 6607 16983
rect 6822 16980 6828 16992
rect 6595 16952 6828 16980
rect 6595 16949 6607 16952
rect 6549 16943 6607 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 9398 16980 9404 16992
rect 7708 16952 9404 16980
rect 7708 16940 7714 16952
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9916 16952 9965 16980
rect 9916 16940 9922 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 11330 16940 11336 16992
rect 11388 16980 11394 16992
rect 11808 16989 11836 17020
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 12805 17011 12863 17017
rect 12912 16992 12940 17088
rect 15096 17079 15108 17088
rect 15160 17116 15166 17128
rect 15378 17116 15384 17128
rect 15160 17088 15384 17116
rect 15102 17076 15108 17079
rect 15160 17076 15166 17088
rect 15378 17076 15384 17088
rect 15436 17076 15442 17128
rect 18782 17125 18788 17128
rect 18509 17119 18567 17125
rect 18509 17085 18521 17119
rect 18555 17085 18567 17119
rect 18776 17116 18788 17125
rect 18743 17088 18788 17116
rect 18509 17079 18567 17085
rect 18776 17079 18788 17088
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11388 16952 11805 16980
rect 11388 16940 11394 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11793 16943 11851 16949
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 12124 16952 12173 16980
rect 12124 16940 12130 16952
rect 12161 16949 12173 16952
rect 12207 16949 12219 16983
rect 12161 16943 12219 16949
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12526 16980 12532 16992
rect 12483 16952 12532 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 14274 16980 14280 16992
rect 14235 16952 14280 16980
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 15838 16940 15844 16992
rect 15896 16980 15902 16992
rect 16209 16983 16267 16989
rect 16209 16980 16221 16983
rect 15896 16952 16221 16980
rect 15896 16940 15902 16952
rect 16209 16949 16221 16952
rect 16255 16949 16267 16983
rect 16209 16943 16267 16949
rect 16390 16940 16396 16992
rect 16448 16980 16454 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16448 16952 16865 16980
rect 16448 16940 16454 16952
rect 16853 16949 16865 16952
rect 16899 16980 16911 16983
rect 18417 16983 18475 16989
rect 18417 16980 18429 16983
rect 16899 16952 18429 16980
rect 16899 16949 16911 16952
rect 16853 16943 16911 16949
rect 18417 16949 18429 16952
rect 18463 16980 18475 16983
rect 18524 16980 18552 17079
rect 18782 17076 18788 17079
rect 18840 17076 18846 17128
rect 20993 17051 21051 17057
rect 20993 17017 21005 17051
rect 21039 17048 21051 17051
rect 21634 17048 21640 17060
rect 21039 17020 21640 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 21634 17008 21640 17020
rect 21692 17048 21698 17060
rect 22281 17051 22339 17057
rect 22281 17048 22293 17051
rect 21692 17020 22293 17048
rect 21692 17008 21698 17020
rect 22281 17017 22293 17020
rect 22327 17017 22339 17051
rect 22480 17048 22508 17147
rect 25406 17144 25412 17196
rect 25464 17184 25470 17196
rect 27065 17187 27123 17193
rect 27065 17184 27077 17187
rect 25464 17156 27077 17184
rect 25464 17144 25470 17156
rect 27065 17153 27077 17156
rect 27111 17184 27123 17187
rect 27522 17184 27528 17196
rect 27111 17156 27528 17184
rect 27111 17153 27123 17156
rect 27065 17147 27123 17153
rect 27522 17144 27528 17156
rect 27580 17184 27586 17196
rect 27893 17187 27951 17193
rect 27893 17184 27905 17187
rect 27580 17156 27905 17184
rect 27580 17144 27586 17156
rect 27893 17153 27905 17156
rect 27939 17184 27951 17187
rect 28166 17184 28172 17196
rect 27939 17156 28172 17184
rect 27939 17153 27951 17156
rect 27893 17147 27951 17153
rect 28166 17144 28172 17156
rect 28224 17144 28230 17196
rect 26326 17076 26332 17128
rect 26384 17116 26390 17128
rect 26973 17119 27031 17125
rect 26973 17116 26985 17119
rect 26384 17088 26985 17116
rect 26384 17076 26390 17088
rect 26973 17085 26985 17088
rect 27019 17085 27031 17119
rect 26973 17079 27031 17085
rect 24118 17048 24124 17060
rect 22480 17020 24124 17048
rect 22281 17011 22339 17017
rect 24118 17008 24124 17020
rect 24176 17048 24182 17060
rect 24274 17051 24332 17057
rect 24274 17048 24286 17051
rect 24176 17020 24286 17048
rect 24176 17008 24182 17020
rect 24274 17017 24286 17020
rect 24320 17017 24332 17051
rect 24274 17011 24332 17017
rect 26237 17051 26295 17057
rect 26237 17017 26249 17051
rect 26283 17048 26295 17051
rect 26881 17051 26939 17057
rect 26881 17048 26893 17051
rect 26283 17020 26893 17048
rect 26283 17017 26295 17020
rect 26237 17011 26295 17017
rect 26881 17017 26893 17020
rect 26927 17048 26939 17051
rect 27246 17048 27252 17060
rect 26927 17020 27252 17048
rect 26927 17017 26939 17020
rect 26881 17011 26939 17017
rect 27246 17008 27252 17020
rect 27304 17008 27310 17060
rect 27430 17008 27436 17060
rect 27488 17048 27494 17060
rect 28261 17051 28319 17057
rect 28261 17048 28273 17051
rect 27488 17020 28273 17048
rect 27488 17008 27494 17020
rect 28261 17017 28273 17020
rect 28307 17017 28319 17051
rect 28261 17011 28319 17017
rect 18966 16980 18972 16992
rect 18463 16952 18972 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19058 16940 19064 16992
rect 19116 16980 19122 16992
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 19116 16952 19901 16980
rect 19116 16940 19122 16952
rect 19889 16949 19901 16952
rect 19935 16980 19947 16983
rect 20254 16980 20260 16992
rect 19935 16952 20260 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 22186 16980 22192 16992
rect 22147 16952 22192 16980
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 23477 16983 23535 16989
rect 23477 16949 23489 16983
rect 23523 16980 23535 16983
rect 25409 16983 25467 16989
rect 25409 16980 25421 16983
rect 23523 16952 25421 16980
rect 23523 16949 23535 16952
rect 23477 16943 23535 16949
rect 25409 16949 25421 16952
rect 25455 16980 25467 16983
rect 25498 16980 25504 16992
rect 25455 16952 25504 16980
rect 25455 16949 25467 16952
rect 25409 16943 25467 16949
rect 25498 16940 25504 16952
rect 25556 16940 25562 16992
rect 26418 16980 26424 16992
rect 26379 16952 26424 16980
rect 26418 16940 26424 16952
rect 26476 16940 26482 16992
rect 27617 16983 27675 16989
rect 27617 16949 27629 16983
rect 27663 16980 27675 16983
rect 27798 16980 27804 16992
rect 27663 16952 27804 16980
rect 27663 16949 27675 16952
rect 27617 16943 27675 16949
rect 27798 16940 27804 16952
rect 27856 16940 27862 16992
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 2832 16748 4077 16776
rect 2832 16736 2838 16748
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4430 16776 4436 16788
rect 4391 16748 4436 16776
rect 4065 16739 4123 16745
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 5534 16776 5540 16788
rect 5495 16748 5540 16776
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 6457 16779 6515 16785
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 6730 16776 6736 16788
rect 6503 16748 6736 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 6825 16779 6883 16785
rect 6825 16745 6837 16779
rect 6871 16776 6883 16779
rect 6914 16776 6920 16788
rect 6871 16748 6920 16776
rect 6871 16745 6883 16748
rect 6825 16739 6883 16745
rect 6914 16736 6920 16748
rect 6972 16776 6978 16788
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 6972 16748 8033 16776
rect 6972 16736 6978 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 8389 16779 8447 16785
rect 8389 16776 8401 16779
rect 8352 16748 8401 16776
rect 8352 16736 8358 16748
rect 8389 16745 8401 16748
rect 8435 16745 8447 16779
rect 10410 16776 10416 16788
rect 10371 16748 10416 16776
rect 8389 16739 8447 16745
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 13081 16779 13139 16785
rect 13081 16745 13093 16779
rect 13127 16776 13139 16779
rect 13814 16776 13820 16788
rect 13127 16748 13820 16776
rect 13127 16745 13139 16748
rect 13081 16739 13139 16745
rect 13814 16736 13820 16748
rect 13872 16736 13878 16788
rect 14090 16776 14096 16788
rect 14051 16748 14096 16776
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 15286 16776 15292 16788
rect 15247 16748 15292 16776
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 17218 16776 17224 16788
rect 16356 16748 17224 16776
rect 16356 16736 16362 16748
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 17954 16776 17960 16788
rect 17368 16748 17413 16776
rect 17915 16748 17960 16776
rect 17368 16736 17374 16748
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18506 16776 18512 16788
rect 18467 16748 18512 16776
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19521 16779 19579 16785
rect 19521 16776 19533 16779
rect 19484 16748 19533 16776
rect 19484 16736 19490 16748
rect 19521 16745 19533 16748
rect 19567 16745 19579 16779
rect 19521 16739 19579 16745
rect 21818 16736 21824 16788
rect 21876 16776 21882 16788
rect 22186 16776 22192 16788
rect 21876 16748 22192 16776
rect 21876 16736 21882 16748
rect 22186 16736 22192 16748
rect 22244 16736 22250 16788
rect 24118 16776 24124 16788
rect 24079 16748 24124 16776
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25498 16736 25504 16788
rect 25556 16776 25562 16788
rect 26145 16779 26203 16785
rect 26145 16776 26157 16779
rect 25556 16748 26157 16776
rect 25556 16736 25562 16748
rect 26145 16745 26157 16748
rect 26191 16776 26203 16779
rect 26234 16776 26240 16788
rect 26191 16748 26240 16776
rect 26191 16745 26203 16748
rect 26145 16739 26203 16745
rect 26234 16736 26240 16748
rect 26292 16736 26298 16788
rect 26326 16736 26332 16788
rect 26384 16776 26390 16788
rect 26513 16779 26571 16785
rect 26513 16776 26525 16779
rect 26384 16748 26525 16776
rect 26384 16736 26390 16748
rect 26513 16745 26525 16748
rect 26559 16745 26571 16779
rect 26513 16739 26571 16745
rect 2041 16711 2099 16717
rect 2041 16677 2053 16711
rect 2087 16708 2099 16711
rect 2590 16708 2596 16720
rect 2087 16680 2596 16708
rect 2087 16677 2099 16680
rect 2041 16671 2099 16677
rect 2590 16668 2596 16680
rect 2648 16668 2654 16720
rect 7466 16708 7472 16720
rect 7427 16680 7472 16708
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 8481 16711 8539 16717
rect 8481 16708 8493 16711
rect 8312 16680 8493 16708
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2774 16640 2780 16652
rect 2179 16612 2780 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 2774 16600 2780 16612
rect 2832 16640 2838 16652
rect 5261 16643 5319 16649
rect 2832 16612 2877 16640
rect 2832 16600 2838 16612
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 5307 16612 5488 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 2314 16572 2320 16584
rect 2275 16544 2320 16572
rect 2314 16532 2320 16544
rect 2372 16572 2378 16584
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 2372 16544 3433 16572
rect 2372 16532 2378 16544
rect 3421 16541 3433 16544
rect 3467 16572 3479 16575
rect 3694 16572 3700 16584
rect 3467 16544 3700 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 3694 16532 3700 16544
rect 3752 16572 3758 16584
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 3752 16544 3801 16572
rect 3752 16532 3758 16544
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 4522 16572 4528 16584
rect 4483 16544 4528 16572
rect 3789 16535 3847 16541
rect 1486 16464 1492 16516
rect 1544 16504 1550 16516
rect 2774 16504 2780 16516
rect 1544 16476 2780 16504
rect 1544 16464 1550 16476
rect 2774 16464 2780 16476
rect 2832 16504 2838 16516
rect 3053 16507 3111 16513
rect 3053 16504 3065 16507
rect 2832 16476 3065 16504
rect 2832 16464 2838 16476
rect 3053 16473 3065 16476
rect 3099 16504 3111 16507
rect 3510 16504 3516 16516
rect 3099 16476 3516 16504
rect 3099 16473 3111 16476
rect 3053 16467 3111 16473
rect 3510 16464 3516 16476
rect 3568 16464 3574 16516
rect 3804 16504 3832 16535
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 5460 16572 5488 16612
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 5905 16643 5963 16649
rect 5905 16640 5917 16643
rect 5592 16612 5917 16640
rect 5592 16600 5598 16612
rect 5905 16609 5917 16612
rect 5951 16609 5963 16643
rect 8312 16640 8340 16680
rect 8481 16677 8493 16680
rect 8527 16677 8539 16711
rect 8481 16671 8539 16677
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 10842 16711 10900 16717
rect 10842 16708 10854 16711
rect 10376 16680 10854 16708
rect 10376 16668 10382 16680
rect 10842 16677 10854 16680
rect 10888 16708 10900 16711
rect 10962 16708 10968 16720
rect 10888 16680 10968 16708
rect 10888 16677 10900 16680
rect 10842 16671 10900 16677
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 12434 16668 12440 16720
rect 12492 16708 12498 16720
rect 13541 16711 13599 16717
rect 13541 16708 13553 16711
rect 12492 16680 13553 16708
rect 12492 16668 12498 16680
rect 13541 16677 13553 16680
rect 13587 16677 13599 16711
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 13541 16671 13599 16677
rect 15212 16680 15761 16708
rect 13446 16640 13452 16652
rect 5905 16603 5963 16609
rect 8220 16612 8340 16640
rect 13407 16612 13452 16640
rect 5626 16572 5632 16584
rect 5460 16544 5632 16572
rect 4617 16535 4675 16541
rect 4632 16504 4660 16535
rect 5626 16532 5632 16544
rect 5684 16532 5690 16584
rect 6914 16572 6920 16584
rect 6875 16544 6920 16572
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7650 16572 7656 16584
rect 7147 16544 7656 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 3804 16476 4660 16504
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16504 6423 16507
rect 7116 16504 7144 16535
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 8220 16572 8248 16612
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 15212 16640 15240 16680
rect 15749 16677 15761 16680
rect 15795 16677 15807 16711
rect 17972 16708 18000 16736
rect 18969 16711 19027 16717
rect 18969 16708 18981 16711
rect 17972 16680 18981 16708
rect 15749 16671 15807 16677
rect 18969 16677 18981 16680
rect 19015 16677 19027 16711
rect 18969 16671 19027 16677
rect 21545 16711 21603 16717
rect 21545 16677 21557 16711
rect 21591 16708 21603 16711
rect 22002 16708 22008 16720
rect 21591 16680 22008 16708
rect 21591 16677 21603 16680
rect 21545 16671 21603 16677
rect 22002 16668 22008 16680
rect 22060 16708 22066 16720
rect 22094 16708 22100 16720
rect 22060 16680 22100 16708
rect 22060 16668 22066 16680
rect 22094 16668 22100 16680
rect 22152 16668 22158 16720
rect 25222 16708 25228 16720
rect 25135 16680 25228 16708
rect 25222 16668 25228 16680
rect 25280 16708 25286 16720
rect 27617 16711 27675 16717
rect 27617 16708 27629 16711
rect 25280 16680 27629 16708
rect 25280 16668 25286 16680
rect 27617 16677 27629 16680
rect 27663 16677 27675 16711
rect 27617 16671 27675 16677
rect 15654 16640 15660 16652
rect 15120 16612 15240 16640
rect 15615 16612 15660 16640
rect 7800 16544 8248 16572
rect 7800 16532 7806 16544
rect 8570 16532 8576 16584
rect 8628 16572 8634 16584
rect 9858 16572 9864 16584
rect 8628 16544 9864 16572
rect 8628 16532 8634 16544
rect 9858 16532 9864 16544
rect 9916 16572 9922 16584
rect 10226 16572 10232 16584
rect 9916 16544 10232 16572
rect 9916 16532 9922 16544
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 10594 16572 10600 16584
rect 10555 16544 10600 16572
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 13725 16575 13783 16581
rect 13725 16572 13737 16575
rect 13688 16544 13737 16572
rect 13688 16532 13694 16544
rect 13725 16541 13737 16544
rect 13771 16541 13783 16575
rect 13725 16535 13783 16541
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 15120 16572 15148 16612
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 16724 16612 16896 16640
rect 16724 16600 16730 16612
rect 13872 16544 15148 16572
rect 13872 16532 13878 16544
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15804 16544 15853 16572
rect 15804 16532 15810 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 6411 16476 7144 16504
rect 6411 16473 6423 16476
rect 6365 16467 6423 16473
rect 11698 16464 11704 16516
rect 11756 16504 11762 16516
rect 11977 16507 12035 16513
rect 11977 16504 11989 16507
rect 11756 16476 11989 16504
rect 11756 16464 11762 16476
rect 11977 16473 11989 16476
rect 12023 16473 12035 16507
rect 11977 16467 12035 16473
rect 14274 16464 14280 16516
rect 14332 16504 14338 16516
rect 15764 16504 15792 16532
rect 16868 16513 16896 16612
rect 18138 16600 18144 16652
rect 18196 16640 18202 16652
rect 18877 16643 18935 16649
rect 18877 16640 18889 16643
rect 18196 16612 18889 16640
rect 18196 16600 18202 16612
rect 18877 16609 18889 16612
rect 18923 16609 18935 16643
rect 21893 16643 21951 16649
rect 21893 16640 21905 16643
rect 18877 16603 18935 16609
rect 21560 16612 21905 16640
rect 21560 16584 21588 16612
rect 21893 16609 21905 16612
rect 21939 16609 21951 16643
rect 21893 16603 21951 16609
rect 24765 16643 24823 16649
rect 24765 16609 24777 16643
rect 24811 16640 24823 16643
rect 25774 16640 25780 16652
rect 24811 16612 25780 16640
rect 24811 16609 24823 16612
rect 24765 16603 24823 16609
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 26878 16640 26884 16652
rect 26160 16612 26884 16640
rect 17402 16572 17408 16584
rect 17363 16544 17408 16572
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 19058 16572 19064 16584
rect 19019 16544 19064 16572
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 21542 16532 21548 16584
rect 21600 16532 21606 16584
rect 21637 16575 21695 16581
rect 21637 16541 21649 16575
rect 21683 16541 21695 16575
rect 25314 16572 25320 16584
rect 25275 16544 25320 16572
rect 21637 16535 21695 16541
rect 14332 16476 15792 16504
rect 16853 16507 16911 16513
rect 14332 16464 14338 16476
rect 16853 16473 16865 16507
rect 16899 16473 16911 16507
rect 16853 16467 16911 16473
rect 7926 16436 7932 16448
rect 7839 16408 7932 16436
rect 7926 16396 7932 16408
rect 7984 16436 7990 16448
rect 8478 16436 8484 16448
rect 7984 16408 8484 16436
rect 7984 16396 7990 16408
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 8720 16408 9045 16436
rect 8720 16396 8726 16408
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 9033 16399 9091 16405
rect 15105 16439 15163 16445
rect 15105 16405 15117 16439
rect 15151 16436 15163 16439
rect 15562 16436 15568 16448
rect 15151 16408 15568 16436
rect 15151 16405 15163 16408
rect 15105 16399 15163 16405
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 18417 16439 18475 16445
rect 18417 16405 18429 16439
rect 18463 16436 18475 16439
rect 18506 16436 18512 16448
rect 18463 16408 18512 16436
rect 18463 16405 18475 16408
rect 18417 16399 18475 16405
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 21174 16436 21180 16448
rect 21135 16408 21180 16436
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 21652 16436 21680 16535
rect 25314 16532 25320 16544
rect 25372 16532 25378 16584
rect 25406 16532 25412 16584
rect 25464 16572 25470 16584
rect 26160 16572 26188 16612
rect 26878 16600 26884 16612
rect 26936 16600 26942 16652
rect 26973 16643 27031 16649
rect 26973 16609 26985 16643
rect 27019 16609 27031 16643
rect 26973 16603 27031 16609
rect 25464 16544 25509 16572
rect 25792 16544 26188 16572
rect 25464 16532 25470 16544
rect 25498 16464 25504 16516
rect 25556 16504 25562 16516
rect 25792 16504 25820 16544
rect 25556 16476 25820 16504
rect 25556 16464 25562 16476
rect 25866 16464 25872 16516
rect 25924 16504 25930 16516
rect 26988 16504 27016 16603
rect 27065 16575 27123 16581
rect 27065 16541 27077 16575
rect 27111 16541 27123 16575
rect 27065 16535 27123 16541
rect 25924 16476 27016 16504
rect 25924 16464 25930 16476
rect 21910 16436 21916 16448
rect 21652 16408 21916 16436
rect 21910 16396 21916 16408
rect 21968 16436 21974 16448
rect 22278 16436 22284 16448
rect 21968 16408 22284 16436
rect 21968 16396 21974 16408
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 22370 16396 22376 16448
rect 22428 16436 22434 16448
rect 23017 16439 23075 16445
rect 23017 16436 23029 16439
rect 22428 16408 23029 16436
rect 22428 16396 22434 16408
rect 23017 16405 23029 16408
rect 23063 16405 23075 16439
rect 23750 16436 23756 16448
rect 23711 16408 23756 16436
rect 23017 16399 23075 16405
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 26326 16396 26332 16448
rect 26384 16436 26390 16448
rect 27080 16436 27108 16535
rect 26384 16408 27108 16436
rect 26384 16396 26390 16408
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 3145 16235 3203 16241
rect 3145 16201 3157 16235
rect 3191 16232 3203 16235
rect 3326 16232 3332 16244
rect 3191 16204 3332 16232
rect 3191 16201 3203 16204
rect 3145 16195 3203 16201
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 4430 16192 4436 16244
rect 4488 16232 4494 16244
rect 4525 16235 4583 16241
rect 4525 16232 4537 16235
rect 4488 16204 4537 16232
rect 4488 16192 4494 16204
rect 4525 16201 4537 16204
rect 4571 16201 4583 16235
rect 4525 16195 4583 16201
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 5258 16232 5264 16244
rect 5215 16204 5264 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6454 16192 6460 16244
rect 6512 16232 6518 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6512 16204 6837 16232
rect 6512 16192 6518 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 6825 16195 6883 16201
rect 8113 16235 8171 16241
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 8294 16232 8300 16244
rect 8159 16204 8300 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 9858 16232 9864 16244
rect 9819 16204 9864 16232
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 11054 16232 11060 16244
rect 11015 16204 11060 16232
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 11517 16235 11575 16241
rect 11517 16201 11529 16235
rect 11563 16232 11575 16235
rect 12158 16232 12164 16244
rect 11563 16204 12164 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 16301 16235 16359 16241
rect 16301 16201 16313 16235
rect 16347 16232 16359 16235
rect 16390 16232 16396 16244
rect 16347 16204 16396 16232
rect 16347 16201 16359 16204
rect 16301 16195 16359 16201
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 17218 16232 17224 16244
rect 17179 16204 17224 16232
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 18138 16192 18144 16244
rect 18196 16232 18202 16244
rect 18233 16235 18291 16241
rect 18233 16232 18245 16235
rect 18196 16204 18245 16232
rect 18196 16192 18202 16204
rect 18233 16201 18245 16204
rect 18279 16201 18291 16235
rect 18233 16195 18291 16201
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 21818 16232 21824 16244
rect 21232 16204 21824 16232
rect 21232 16192 21238 16204
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 24912 16204 25053 16232
rect 24912 16192 24918 16204
rect 25041 16201 25053 16204
rect 25087 16201 25099 16235
rect 27522 16232 27528 16244
rect 27483 16204 27528 16232
rect 25041 16195 25099 16201
rect 27522 16192 27528 16204
rect 27580 16192 27586 16244
rect 14093 16167 14151 16173
rect 14093 16133 14105 16167
rect 14139 16133 14151 16167
rect 14642 16164 14648 16176
rect 14603 16136 14648 16164
rect 14093 16127 14151 16133
rect 2225 16099 2283 16105
rect 2225 16065 2237 16099
rect 2271 16096 2283 16099
rect 2314 16096 2320 16108
rect 2271 16068 2320 16096
rect 2271 16065 2283 16068
rect 2225 16059 2283 16065
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2590 16096 2596 16108
rect 2551 16068 2596 16096
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 3694 16096 3700 16108
rect 3655 16068 3700 16096
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 5859 16068 5893 16096
rect 6840 16068 7389 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 1762 15988 1768 16040
rect 1820 16028 1826 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1820 16000 2053 16028
rect 1820 15988 1826 16000
rect 2041 15997 2053 16000
rect 2087 16028 2099 16031
rect 2682 16028 2688 16040
rect 2087 16000 2688 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 2682 15988 2688 16000
rect 2740 15988 2746 16040
rect 4706 15988 4712 16040
rect 4764 16028 4770 16040
rect 5828 16028 5856 16059
rect 6840 16040 6868 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 10594 16056 10600 16108
rect 10652 16096 10658 16108
rect 10689 16099 10747 16105
rect 10689 16096 10701 16099
rect 10652 16068 10701 16096
rect 10652 16056 10658 16068
rect 10689 16065 10701 16068
rect 10735 16096 10747 16099
rect 11974 16096 11980 16108
rect 10735 16068 11980 16096
rect 10735 16065 10747 16068
rect 10689 16059 10747 16065
rect 11974 16056 11980 16068
rect 12032 16096 12038 16108
rect 12710 16096 12716 16108
rect 12032 16068 12716 16096
rect 12032 16056 12038 16068
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 14108 16096 14136 16127
rect 14642 16124 14648 16136
rect 14700 16124 14706 16176
rect 16945 16167 17003 16173
rect 16945 16133 16957 16167
rect 16991 16164 17003 16167
rect 17310 16164 17316 16176
rect 16991 16136 17316 16164
rect 16991 16133 17003 16136
rect 16945 16127 17003 16133
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 20993 16167 21051 16173
rect 20993 16133 21005 16167
rect 21039 16164 21051 16167
rect 21358 16164 21364 16176
rect 21039 16136 21364 16164
rect 21039 16133 21051 16136
rect 20993 16127 21051 16133
rect 21358 16124 21364 16136
rect 21416 16124 21422 16176
rect 25498 16124 25504 16176
rect 25556 16164 25562 16176
rect 25593 16167 25651 16173
rect 25593 16164 25605 16167
rect 25556 16136 25605 16164
rect 25556 16124 25562 16136
rect 25593 16133 25605 16136
rect 25639 16133 25651 16167
rect 25593 16127 25651 16133
rect 15562 16096 15568 16108
rect 14108 16068 15568 16096
rect 15562 16056 15568 16068
rect 15620 16096 15626 16108
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15620 16068 15761 16096
rect 15620 16056 15626 16068
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 22370 16096 22376 16108
rect 22331 16068 22376 16096
rect 15749 16059 15807 16065
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 6181 16031 6239 16037
rect 6181 16028 6193 16031
rect 4764 16000 6193 16028
rect 4764 15988 4770 16000
rect 6181 15997 6193 16000
rect 6227 16028 6239 16031
rect 6362 16028 6368 16040
rect 6227 16000 6368 16028
rect 6227 15997 6239 16000
rect 6181 15991 6239 15997
rect 6362 15988 6368 16000
rect 6420 16028 6426 16040
rect 6822 16028 6828 16040
rect 6420 16000 6828 16028
rect 6420 15988 6426 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 16028 7343 16031
rect 7466 16028 7472 16040
rect 7331 16000 7472 16028
rect 7331 15997 7343 16000
rect 7285 15991 7343 15997
rect 7466 15988 7472 16000
rect 7524 15988 7530 16040
rect 8478 16028 8484 16040
rect 8439 16000 8484 16028
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 12986 16037 12992 16040
rect 12980 16028 12992 16037
rect 12820 16000 12992 16028
rect 2866 15920 2872 15972
rect 2924 15960 2930 15972
rect 3605 15963 3663 15969
rect 3605 15960 3617 15963
rect 2924 15932 3617 15960
rect 2924 15920 2930 15932
rect 3605 15929 3617 15932
rect 3651 15929 3663 15963
rect 5074 15960 5080 15972
rect 4987 15932 5080 15960
rect 3605 15923 3663 15929
rect 5074 15920 5080 15932
rect 5132 15960 5138 15972
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 5132 15932 5549 15960
rect 5132 15920 5138 15932
rect 5537 15929 5549 15932
rect 5583 15960 5595 15963
rect 5810 15960 5816 15972
rect 5583 15932 5816 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 8662 15920 8668 15972
rect 8720 15969 8726 15972
rect 8720 15963 8784 15969
rect 8720 15929 8738 15963
rect 8772 15929 8784 15963
rect 8720 15923 8784 15929
rect 11885 15963 11943 15969
rect 11885 15929 11897 15963
rect 11931 15960 11943 15963
rect 12820 15960 12848 16000
rect 12980 15991 12992 16000
rect 12986 15988 12992 15991
rect 13044 15988 13050 16040
rect 14642 15988 14648 16040
rect 14700 16028 14706 16040
rect 15654 16028 15660 16040
rect 14700 16000 15660 16028
rect 14700 15988 14706 16000
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 18417 16031 18475 16037
rect 18417 15997 18429 16031
rect 18463 15997 18475 16031
rect 18417 15991 18475 15997
rect 11931 15932 12848 15960
rect 11931 15929 11943 15932
rect 11885 15923 11943 15929
rect 8720 15920 8726 15923
rect 15470 15920 15476 15972
rect 15528 15960 15534 15972
rect 15565 15963 15623 15969
rect 15565 15960 15577 15963
rect 15528 15932 15577 15960
rect 15528 15920 15534 15932
rect 15565 15929 15577 15932
rect 15611 15960 15623 15963
rect 16390 15960 16396 15972
rect 15611 15932 16396 15960
rect 15611 15929 15623 15932
rect 15565 15923 15623 15929
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 17126 15920 17132 15972
rect 17184 15960 17190 15972
rect 17865 15963 17923 15969
rect 17865 15960 17877 15963
rect 17184 15932 17877 15960
rect 17184 15920 17190 15932
rect 17865 15929 17877 15932
rect 17911 15960 17923 15963
rect 18432 15960 18460 15991
rect 18506 15988 18512 16040
rect 18564 16028 18570 16040
rect 18673 16031 18731 16037
rect 18673 16028 18685 16031
rect 18564 16000 18685 16028
rect 18564 15988 18570 16000
rect 18673 15997 18685 16000
rect 18719 15997 18731 16031
rect 18673 15991 18731 15997
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 22462 16028 22468 16040
rect 22327 16000 22468 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 22462 15988 22468 16000
rect 22520 16028 22526 16040
rect 22833 16031 22891 16037
rect 22833 16028 22845 16031
rect 22520 16000 22845 16028
rect 22520 15988 22526 16000
rect 22833 15997 22845 16000
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 23661 16031 23719 16037
rect 23661 15997 23673 16031
rect 23707 15997 23719 16031
rect 23661 15991 23719 15997
rect 18966 15960 18972 15972
rect 17911 15932 18972 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 18966 15920 18972 15932
rect 19024 15920 19030 15972
rect 23385 15963 23443 15969
rect 23385 15960 23397 15963
rect 21928 15932 23397 15960
rect 21928 15904 21956 15932
rect 23385 15929 23397 15932
rect 23431 15960 23443 15963
rect 23676 15960 23704 15991
rect 23750 15988 23756 16040
rect 23808 16028 23814 16040
rect 23917 16031 23975 16037
rect 23917 16028 23929 16031
rect 23808 16000 23929 16028
rect 23808 15988 23814 16000
rect 23917 15997 23929 16000
rect 23963 15997 23975 16031
rect 26142 16028 26148 16040
rect 26103 16000 26148 16028
rect 23917 15991 23975 15997
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 23431 15932 23704 15960
rect 23431 15929 23443 15932
rect 23385 15923 23443 15929
rect 24946 15920 24952 15972
rect 25004 15960 25010 15972
rect 25866 15960 25872 15972
rect 25004 15932 25872 15960
rect 25004 15920 25010 15932
rect 25866 15920 25872 15932
rect 25924 15960 25930 15972
rect 25961 15963 26019 15969
rect 25961 15960 25973 15963
rect 25924 15932 25973 15960
rect 25924 15920 25930 15932
rect 25961 15929 25973 15932
rect 26007 15929 26019 15963
rect 25961 15923 26019 15929
rect 26326 15920 26332 15972
rect 26384 15969 26390 15972
rect 26384 15963 26448 15969
rect 26384 15929 26402 15963
rect 26436 15960 26448 15963
rect 28077 15963 28135 15969
rect 28077 15960 28089 15963
rect 26436 15932 28089 15960
rect 26436 15929 26448 15932
rect 26384 15923 26448 15929
rect 28077 15929 28089 15932
rect 28123 15929 28135 15963
rect 28077 15923 28135 15929
rect 26384 15920 26390 15923
rect 1578 15852 1584 15904
rect 1636 15892 1642 15904
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1636 15864 1961 15892
rect 1636 15852 1642 15864
rect 1949 15861 1961 15864
rect 1995 15861 2007 15895
rect 1949 15855 2007 15861
rect 3053 15895 3111 15901
rect 3053 15861 3065 15895
rect 3099 15892 3111 15895
rect 3510 15892 3516 15904
rect 3099 15864 3516 15892
rect 3099 15861 3111 15864
rect 3053 15855 3111 15861
rect 3510 15852 3516 15864
rect 3568 15892 3574 15904
rect 3786 15892 3792 15904
rect 3568 15864 3792 15892
rect 3568 15852 3574 15864
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 4522 15892 4528 15904
rect 4295 15864 4528 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 6546 15852 6552 15864
rect 6604 15892 6610 15904
rect 7190 15892 7196 15904
rect 6604 15864 7196 15892
rect 6604 15852 6610 15864
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 11572 15864 12173 15892
rect 11572 15852 11578 15864
rect 12161 15861 12173 15864
rect 12207 15892 12219 15895
rect 12434 15892 12440 15904
rect 12207 15864 12440 15892
rect 12207 15861 12219 15864
rect 12161 15855 12219 15861
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 15010 15892 15016 15904
rect 14971 15864 15016 15892
rect 15010 15852 15016 15864
rect 15068 15852 15074 15904
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 19797 15895 19855 15901
rect 19797 15892 19809 15895
rect 19392 15864 19809 15892
rect 19392 15852 19398 15864
rect 19797 15861 19809 15864
rect 19843 15861 19855 15895
rect 19797 15855 19855 15861
rect 21361 15895 21419 15901
rect 21361 15861 21373 15895
rect 21407 15892 21419 15895
rect 21542 15892 21548 15904
rect 21407 15864 21548 15892
rect 21407 15861 21419 15864
rect 21361 15855 21419 15861
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 21726 15892 21732 15904
rect 21687 15864 21732 15892
rect 21726 15852 21732 15864
rect 21784 15892 21790 15904
rect 21910 15892 21916 15904
rect 21784 15864 21916 15892
rect 21784 15852 21790 15864
rect 21910 15852 21916 15864
rect 21968 15852 21974 15904
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22189 15895 22247 15901
rect 22189 15892 22201 15895
rect 22152 15864 22201 15892
rect 22152 15852 22158 15864
rect 22189 15861 22201 15864
rect 22235 15861 22247 15895
rect 22189 15855 22247 15861
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1762 15688 1768 15700
rect 1723 15660 1768 15688
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 2774 15688 2780 15700
rect 2735 15660 2780 15688
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 3605 15691 3663 15697
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 3694 15688 3700 15700
rect 3651 15660 3700 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 3694 15648 3700 15660
rect 3752 15688 3758 15700
rect 4249 15691 4307 15697
rect 4249 15688 4261 15691
rect 3752 15660 4261 15688
rect 3752 15648 3758 15660
rect 4249 15657 4261 15660
rect 4295 15657 4307 15691
rect 6822 15688 6828 15700
rect 6783 15660 6828 15688
rect 4249 15651 4307 15657
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 6972 15660 8033 15688
rect 6972 15648 6978 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 13173 15691 13231 15697
rect 13173 15657 13185 15691
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 5068 15623 5126 15629
rect 5068 15589 5080 15623
rect 5114 15620 5126 15623
rect 5166 15620 5172 15632
rect 5114 15592 5172 15620
rect 5114 15589 5126 15592
rect 5068 15583 5126 15589
rect 5166 15580 5172 15592
rect 5224 15580 5230 15632
rect 13188 15620 13216 15651
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 13872 15660 14657 15688
rect 13872 15648 13878 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 15105 15691 15163 15697
rect 15105 15657 15117 15691
rect 15151 15688 15163 15691
rect 15746 15688 15752 15700
rect 15151 15660 15752 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 15120 15620 15148 15651
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 18414 15688 18420 15700
rect 18375 15660 18420 15688
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 21358 15648 21364 15700
rect 21416 15688 21422 15700
rect 21729 15691 21787 15697
rect 21729 15688 21741 15691
rect 21416 15660 21741 15688
rect 21416 15648 21422 15660
rect 21729 15657 21741 15660
rect 21775 15657 21787 15691
rect 21729 15651 21787 15657
rect 23293 15691 23351 15697
rect 23293 15657 23305 15691
rect 23339 15657 23351 15691
rect 23293 15651 23351 15657
rect 24857 15691 24915 15697
rect 24857 15657 24869 15691
rect 24903 15688 24915 15691
rect 25314 15688 25320 15700
rect 24903 15660 25320 15688
rect 24903 15657 24915 15660
rect 24857 15651 24915 15657
rect 13188 15592 15148 15620
rect 21542 15580 21548 15632
rect 21600 15620 21606 15632
rect 22830 15620 22836 15632
rect 21600 15592 22836 15620
rect 21600 15580 21606 15592
rect 22830 15580 22836 15592
rect 22888 15620 22894 15632
rect 23308 15620 23336 15651
rect 25314 15648 25320 15660
rect 25372 15688 25378 15700
rect 27617 15691 27675 15697
rect 27617 15688 27629 15691
rect 25372 15660 27629 15688
rect 25372 15648 25378 15660
rect 27617 15657 27629 15660
rect 27663 15657 27675 15691
rect 27617 15651 27675 15657
rect 23845 15623 23903 15629
rect 23845 15620 23857 15623
rect 22888 15592 23857 15620
rect 22888 15580 22894 15592
rect 23845 15589 23857 15592
rect 23891 15620 23903 15623
rect 24210 15620 24216 15632
rect 23891 15592 24216 15620
rect 23891 15589 23903 15592
rect 23845 15583 23903 15589
rect 24210 15580 24216 15592
rect 24268 15580 24274 15632
rect 24765 15623 24823 15629
rect 24765 15589 24777 15623
rect 24811 15620 24823 15623
rect 25406 15620 25412 15632
rect 24811 15592 25412 15620
rect 24811 15589 24823 15592
rect 24765 15583 24823 15589
rect 25406 15580 25412 15592
rect 25464 15580 25470 15632
rect 26418 15580 26424 15632
rect 26476 15620 26482 15632
rect 26970 15620 26976 15632
rect 26476 15592 26976 15620
rect 26476 15580 26482 15592
rect 26970 15580 26976 15592
rect 27028 15580 27034 15632
rect 2130 15552 2136 15564
rect 2091 15524 2136 15552
rect 2130 15512 2136 15524
rect 2188 15512 2194 15564
rect 8386 15552 8392 15564
rect 8347 15524 8392 15552
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 8527 15524 9413 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 9401 15521 9413 15524
rect 9447 15521 9459 15555
rect 9401 15515 9459 15521
rect 2222 15484 2228 15496
rect 2183 15456 2228 15484
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2498 15484 2504 15496
rect 2455 15456 2504 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 3145 15351 3203 15357
rect 3145 15348 3157 15351
rect 2924 15320 3157 15348
rect 2924 15308 2930 15320
rect 3145 15317 3157 15320
rect 3191 15317 3203 15351
rect 4706 15348 4712 15360
rect 4667 15320 4712 15348
rect 3145 15311 3203 15317
rect 4706 15308 4712 15320
rect 4764 15308 4770 15360
rect 4816 15348 4844 15447
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8496 15484 8524 15515
rect 10318 15512 10324 15564
rect 10376 15552 10382 15564
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 10376 15524 10609 15552
rect 10376 15512 10382 15524
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 10597 15515 10655 15521
rect 10689 15555 10747 15561
rect 10689 15521 10701 15555
rect 10735 15552 10747 15555
rect 11606 15552 11612 15564
rect 10735 15524 11612 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 11698 15512 11704 15564
rect 11756 15552 11762 15564
rect 12049 15555 12107 15561
rect 12049 15552 12061 15555
rect 11756 15524 12061 15552
rect 11756 15512 11762 15524
rect 12049 15521 12061 15524
rect 12095 15552 12107 15555
rect 13630 15552 13636 15564
rect 12095 15524 13636 15552
rect 12095 15521 12107 15524
rect 12049 15515 12107 15521
rect 13630 15512 13636 15524
rect 13688 15552 13694 15564
rect 15562 15561 15568 15564
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13688 15524 14105 15552
rect 13688 15512 13694 15524
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 15556 15552 15568 15561
rect 15523 15524 15568 15552
rect 14093 15515 14151 15521
rect 15556 15515 15568 15524
rect 15562 15512 15568 15515
rect 15620 15512 15626 15564
rect 18782 15552 18788 15564
rect 18743 15524 18788 15552
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 21453 15555 21511 15561
rect 21453 15521 21465 15555
rect 21499 15552 21511 15555
rect 22002 15552 22008 15564
rect 21499 15524 22008 15552
rect 21499 15521 21511 15524
rect 21453 15515 21511 15521
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 22180 15555 22238 15561
rect 22180 15521 22192 15555
rect 22226 15552 22238 15555
rect 22554 15552 22560 15564
rect 22226 15524 22560 15552
rect 22226 15521 22238 15524
rect 22180 15515 22238 15521
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 24578 15512 24584 15564
rect 24636 15552 24642 15564
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 24636 15524 25237 15552
rect 24636 15512 24642 15524
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25225 15515 25283 15521
rect 26234 15512 26240 15564
rect 26292 15552 26298 15564
rect 26881 15555 26939 15561
rect 26881 15552 26893 15555
rect 26292 15524 26893 15552
rect 26292 15512 26298 15524
rect 26881 15521 26893 15524
rect 26927 15521 26939 15555
rect 26881 15515 26939 15521
rect 8260 15456 8524 15484
rect 8260 15444 8266 15456
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 10870 15484 10876 15496
rect 8628 15456 8721 15484
rect 10831 15456 10876 15484
rect 8628 15444 8634 15456
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 15289 15447 15347 15453
rect 8588 15416 8616 15444
rect 7484 15388 8616 15416
rect 4982 15348 4988 15360
rect 4816 15320 4988 15348
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 5718 15308 5724 15360
rect 5776 15348 5782 15360
rect 6181 15351 6239 15357
rect 6181 15348 6193 15351
rect 5776 15320 6193 15348
rect 5776 15308 5782 15320
rect 6181 15317 6193 15320
rect 6227 15317 6239 15351
rect 6181 15311 6239 15317
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7484 15357 7512 15388
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 10229 15419 10287 15425
rect 10229 15416 10241 15419
rect 9640 15388 10241 15416
rect 9640 15376 9646 15388
rect 10229 15385 10241 15388
rect 10275 15385 10287 15419
rect 10229 15379 10287 15385
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 6972 15320 7481 15348
rect 6972 15308 6978 15320
rect 7469 15317 7481 15320
rect 7515 15317 7527 15351
rect 7469 15311 7527 15317
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 7837 15351 7895 15357
rect 7837 15348 7849 15351
rect 7800 15320 7849 15348
rect 7800 15308 7806 15320
rect 7837 15317 7849 15320
rect 7883 15317 7895 15351
rect 7837 15311 7895 15317
rect 8110 15308 8116 15360
rect 8168 15348 8174 15360
rect 8478 15348 8484 15360
rect 8168 15320 8484 15348
rect 8168 15308 8174 15320
rect 8478 15308 8484 15320
rect 8536 15348 8542 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8536 15320 9045 15348
rect 8536 15308 8542 15320
rect 9033 15317 9045 15320
rect 9079 15348 9091 15351
rect 9674 15348 9680 15360
rect 9079 15320 9680 15348
rect 9079 15317 9091 15320
rect 9033 15311 9091 15317
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 9858 15348 9864 15360
rect 9819 15320 9864 15348
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 11808 15348 11836 15447
rect 11974 15348 11980 15360
rect 11808 15320 11980 15348
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 13630 15348 13636 15360
rect 13504 15320 13636 15348
rect 13504 15308 13510 15320
rect 13630 15308 13636 15320
rect 13688 15348 13694 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13688 15320 13737 15348
rect 13688 15308 13694 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 15304 15348 15332 15447
rect 17954 15444 17960 15496
rect 18012 15484 18018 15496
rect 18877 15487 18935 15493
rect 18877 15484 18889 15487
rect 18012 15456 18889 15484
rect 18012 15444 18018 15456
rect 18877 15453 18889 15456
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 18969 15487 19027 15493
rect 18969 15453 18981 15487
rect 19015 15484 19027 15487
rect 19058 15484 19064 15496
rect 19015 15456 19064 15484
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 18984 15416 19012 15447
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 21726 15484 21732 15496
rect 21468 15456 21732 15484
rect 18432 15388 19012 15416
rect 18432 15360 18460 15388
rect 21468 15360 21496 15456
rect 21726 15444 21732 15456
rect 21784 15484 21790 15496
rect 21913 15487 21971 15493
rect 21913 15484 21925 15487
rect 21784 15456 21925 15484
rect 21784 15444 21790 15456
rect 21913 15453 21925 15456
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 25317 15487 25375 15493
rect 25317 15453 25329 15487
rect 25363 15453 25375 15487
rect 25498 15484 25504 15496
rect 25411 15456 25504 15484
rect 25317 15447 25375 15453
rect 25332 15416 25360 15447
rect 25498 15444 25504 15456
rect 25556 15484 25562 15496
rect 26326 15484 26332 15496
rect 25556 15456 26332 15484
rect 25556 15444 25562 15456
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15484 27215 15487
rect 27522 15484 27528 15496
rect 27203 15456 27528 15484
rect 27203 15453 27215 15456
rect 27157 15447 27215 15453
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 25406 15416 25412 15428
rect 25332 15388 25412 15416
rect 25406 15376 25412 15388
rect 25464 15376 25470 15428
rect 16298 15348 16304 15360
rect 15304 15320 16304 15348
rect 13725 15311 13783 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 16632 15320 16681 15348
rect 16632 15308 16638 15320
rect 16669 15317 16681 15320
rect 16715 15348 16727 15351
rect 17221 15351 17279 15357
rect 17221 15348 17233 15351
rect 16715 15320 17233 15348
rect 16715 15317 16727 15320
rect 16669 15311 16727 15317
rect 17221 15317 17233 15320
rect 17267 15348 17279 15351
rect 17402 15348 17408 15360
rect 17267 15320 17408 15348
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 18325 15351 18383 15357
rect 18325 15317 18337 15351
rect 18371 15348 18383 15351
rect 18414 15348 18420 15360
rect 18371 15320 18420 15348
rect 18371 15317 18383 15320
rect 18325 15311 18383 15317
rect 18414 15308 18420 15320
rect 18472 15308 18478 15360
rect 21450 15308 21456 15360
rect 21508 15308 21514 15360
rect 24118 15308 24124 15360
rect 24176 15348 24182 15360
rect 24213 15351 24271 15357
rect 24213 15348 24225 15351
rect 24176 15320 24225 15348
rect 24176 15308 24182 15320
rect 24213 15317 24225 15320
rect 24259 15317 24271 15351
rect 24213 15311 24271 15317
rect 26237 15351 26295 15357
rect 26237 15317 26249 15351
rect 26283 15348 26295 15351
rect 26326 15348 26332 15360
rect 26283 15320 26332 15348
rect 26283 15317 26295 15320
rect 26237 15311 26295 15317
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 26513 15351 26571 15357
rect 26513 15317 26525 15351
rect 26559 15348 26571 15351
rect 26970 15348 26976 15360
rect 26559 15320 26976 15348
rect 26559 15317 26571 15320
rect 26513 15311 26571 15317
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 3145 15147 3203 15153
rect 3145 15113 3157 15147
rect 3191 15144 3203 15147
rect 3694 15144 3700 15156
rect 3191 15116 3700 15144
rect 3191 15113 3203 15116
rect 3145 15107 3203 15113
rect 3694 15104 3700 15116
rect 3752 15104 3758 15156
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 6641 15147 6699 15153
rect 3844 15116 5284 15144
rect 3844 15104 3850 15116
rect 2774 15036 2780 15088
rect 2832 15076 2838 15088
rect 3050 15076 3056 15088
rect 2832 15048 3056 15076
rect 2832 15036 2838 15048
rect 3050 15036 3056 15048
rect 3108 15076 3114 15088
rect 4065 15079 4123 15085
rect 4065 15076 4077 15079
rect 3108 15048 4077 15076
rect 3108 15036 3114 15048
rect 4065 15045 4077 15048
rect 4111 15076 4123 15079
rect 5256 15076 5284 15116
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 6822 15144 6828 15156
rect 6687 15116 6828 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 8021 15147 8079 15153
rect 8021 15113 8033 15147
rect 8067 15144 8079 15147
rect 8202 15144 8208 15156
rect 8067 15116 8208 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 11606 15144 11612 15156
rect 11567 15116 11612 15144
rect 11606 15104 11612 15116
rect 11664 15144 11670 15156
rect 11882 15144 11888 15156
rect 11664 15116 11888 15144
rect 11664 15104 11670 15116
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 13170 15144 13176 15156
rect 13131 15116 13176 15144
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 18414 15144 18420 15156
rect 18375 15116 18420 15144
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 21634 15104 21640 15156
rect 21692 15144 21698 15156
rect 21729 15147 21787 15153
rect 21729 15144 21741 15147
rect 21692 15116 21741 15144
rect 21692 15104 21698 15116
rect 21729 15113 21741 15116
rect 21775 15113 21787 15147
rect 21729 15107 21787 15113
rect 25314 15104 25320 15156
rect 25372 15144 25378 15156
rect 25961 15147 26019 15153
rect 25961 15144 25973 15147
rect 25372 15116 25973 15144
rect 25372 15104 25378 15116
rect 25961 15113 25973 15116
rect 26007 15113 26019 15147
rect 26418 15144 26424 15156
rect 25961 15107 26019 15113
rect 26068 15116 26424 15144
rect 9122 15076 9128 15088
rect 4111 15048 4292 15076
rect 5256 15048 9128 15076
rect 4111 15045 4123 15048
rect 4065 15039 4123 15045
rect 1486 14900 1492 14952
rect 1544 14940 1550 14952
rect 1765 14943 1823 14949
rect 1765 14940 1777 14943
rect 1544 14912 1777 14940
rect 1544 14900 1550 14912
rect 1765 14909 1777 14912
rect 1811 14940 1823 14943
rect 2792 14940 2820 15036
rect 4264 15017 4292 15048
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 11974 15076 11980 15088
rect 11935 15048 11980 15076
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 7558 15008 7564 15020
rect 7471 14980 7564 15008
rect 4249 14971 4307 14977
rect 1811 14912 2820 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 4062 14940 4068 14952
rect 3844 14912 4068 14940
rect 3844 14900 3850 14912
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4264 14940 4292 14971
rect 7558 14968 7564 14980
rect 7616 15008 7622 15020
rect 8202 15008 8208 15020
rect 7616 14980 8208 15008
rect 7616 14968 7622 14980
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8662 15008 8668 15020
rect 8623 14980 8668 15008
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 13188 15008 13216 15104
rect 14461 15079 14519 15085
rect 14461 15045 14473 15079
rect 14507 15076 14519 15079
rect 14507 15048 15424 15076
rect 14507 15045 14519 15048
rect 14461 15039 14519 15045
rect 15396 15020 15424 15048
rect 21450 15036 21456 15088
rect 21508 15076 21514 15088
rect 22741 15079 22799 15085
rect 22741 15076 22753 15079
rect 21508 15048 22753 15076
rect 21508 15036 21514 15048
rect 22741 15045 22753 15048
rect 22787 15045 22799 15079
rect 22741 15039 22799 15045
rect 25038 15036 25044 15088
rect 25096 15076 25102 15088
rect 25685 15079 25743 15085
rect 25685 15076 25697 15079
rect 25096 15048 25697 15076
rect 25096 15036 25102 15048
rect 25685 15045 25697 15048
rect 25731 15076 25743 15079
rect 26068 15076 26096 15116
rect 26418 15104 26424 15116
rect 26476 15104 26482 15156
rect 25731 15048 26096 15076
rect 25731 15045 25743 15048
rect 25685 15039 25743 15045
rect 13817 15011 13875 15017
rect 13817 15008 13829 15011
rect 13188 14980 13829 15008
rect 13817 14977 13829 14980
rect 13863 15008 13875 15011
rect 13906 15008 13912 15020
rect 13863 14980 13912 15008
rect 13863 14977 13875 14980
rect 13817 14971 13875 14977
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 14001 15011 14059 15017
rect 14001 14977 14013 15011
rect 14047 15008 14059 15011
rect 14826 15008 14832 15020
rect 14047 14980 14832 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15436 14980 15485 15008
rect 15436 14968 15442 14980
rect 15473 14977 15485 14980
rect 15519 15008 15531 15011
rect 15746 15008 15752 15020
rect 15519 14980 15752 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 15746 14968 15752 14980
rect 15804 15008 15810 15020
rect 16482 15008 16488 15020
rect 15804 14980 16488 15008
rect 15804 14968 15810 14980
rect 16482 14968 16488 14980
rect 16540 14968 16546 15020
rect 18969 15011 19027 15017
rect 18969 14977 18981 15011
rect 19015 15008 19027 15011
rect 19058 15008 19064 15020
rect 19015 14980 19064 15008
rect 19015 14977 19027 14980
rect 18969 14971 19027 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 22370 15008 22376 15020
rect 22331 14980 22376 15008
rect 22370 14968 22376 14980
rect 22428 14968 22434 15020
rect 23474 14968 23480 15020
rect 23532 15008 23538 15020
rect 24118 15008 24124 15020
rect 23532 14980 23796 15008
rect 24079 14980 24124 15008
rect 23532 14968 23538 14980
rect 4982 14940 4988 14952
rect 4264 14912 4988 14940
rect 4982 14900 4988 14912
rect 5040 14900 5046 14952
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 5810 14940 5816 14952
rect 5684 14912 5816 14940
rect 5684 14900 5690 14912
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 9585 14943 9643 14949
rect 9585 14909 9597 14943
rect 9631 14940 9643 14943
rect 9674 14940 9680 14952
rect 9631 14912 9680 14940
rect 9631 14909 9643 14912
rect 9585 14903 9643 14909
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 12912 14912 13737 14940
rect 2032 14875 2090 14881
rect 2032 14841 2044 14875
rect 2078 14872 2090 14875
rect 2498 14872 2504 14884
rect 2078 14844 2504 14872
rect 2078 14841 2090 14844
rect 2032 14835 2090 14841
rect 2498 14832 2504 14844
rect 2556 14832 2562 14884
rect 4516 14875 4574 14881
rect 4516 14841 4528 14875
rect 4562 14872 4574 14875
rect 4706 14872 4712 14884
rect 4562 14844 4712 14872
rect 4562 14841 4574 14844
rect 4516 14835 4574 14841
rect 4706 14832 4712 14844
rect 4764 14872 4770 14884
rect 5074 14872 5080 14884
rect 4764 14844 5080 14872
rect 4764 14832 4770 14844
rect 5074 14832 5080 14844
rect 5132 14832 5138 14884
rect 6546 14832 6552 14884
rect 6604 14872 6610 14884
rect 7837 14875 7895 14881
rect 7837 14872 7849 14875
rect 6604 14844 7849 14872
rect 6604 14832 6610 14844
rect 7837 14841 7849 14844
rect 7883 14872 7895 14875
rect 8481 14875 8539 14881
rect 8481 14872 8493 14875
rect 7883 14844 8493 14872
rect 7883 14841 7895 14844
rect 7837 14835 7895 14841
rect 8481 14841 8493 14844
rect 8527 14872 8539 14875
rect 9306 14872 9312 14884
rect 8527 14844 9312 14872
rect 8527 14841 8539 14844
rect 8481 14835 8539 14841
rect 9306 14832 9312 14844
rect 9364 14832 9370 14884
rect 9858 14881 9864 14884
rect 9852 14872 9864 14881
rect 9819 14844 9864 14872
rect 9852 14835 9864 14844
rect 9858 14832 9864 14835
rect 9916 14832 9922 14884
rect 12912 14816 12940 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14940 21327 14943
rect 21726 14940 21732 14952
rect 21315 14912 21732 14940
rect 21315 14909 21327 14912
rect 21269 14903 21327 14909
rect 21726 14900 21732 14912
rect 21784 14940 21790 14952
rect 21784 14912 21956 14940
rect 21784 14900 21790 14912
rect 19334 14881 19340 14884
rect 15289 14875 15347 14881
rect 15289 14872 15301 14875
rect 13372 14844 15301 14872
rect 1210 14764 1216 14816
rect 1268 14804 1274 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 1268 14776 1593 14804
rect 1268 14764 1274 14776
rect 1581 14773 1593 14776
rect 1627 14804 1639 14807
rect 2222 14804 2228 14816
rect 1627 14776 2228 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 3694 14804 3700 14816
rect 3655 14776 3700 14804
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5224 14776 5641 14804
rect 5224 14764 5230 14776
rect 5629 14773 5641 14776
rect 5675 14804 5687 14807
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 5675 14776 6193 14804
rect 5675 14773 5687 14776
rect 5629 14767 5687 14773
rect 6181 14773 6193 14776
rect 6227 14773 6239 14807
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6181 14767 6239 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 7708 14776 8401 14804
rect 7708 14764 7714 14776
rect 8389 14773 8401 14776
rect 8435 14804 8447 14807
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8435 14776 9045 14804
rect 8435 14773 8447 14776
rect 8389 14767 8447 14773
rect 9033 14773 9045 14776
rect 9079 14773 9091 14807
rect 9398 14804 9404 14816
rect 9359 14776 9404 14804
rect 9033 14767 9091 14773
rect 9398 14764 9404 14776
rect 9456 14804 9462 14816
rect 10318 14804 10324 14816
rect 9456 14776 10324 14804
rect 9456 14764 9462 14776
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10965 14807 11023 14813
rect 10965 14804 10977 14807
rect 10652 14776 10977 14804
rect 10652 14764 10658 14776
rect 10965 14773 10977 14776
rect 11011 14773 11023 14807
rect 12894 14804 12900 14816
rect 12855 14776 12900 14804
rect 10965 14767 11023 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13372 14813 13400 14844
rect 15289 14841 15301 14844
rect 15335 14872 15347 14875
rect 16301 14875 16359 14881
rect 16301 14872 16313 14875
rect 15335 14844 16313 14872
rect 15335 14841 15347 14844
rect 15289 14835 15347 14841
rect 16301 14841 16313 14844
rect 16347 14841 16359 14875
rect 19328 14872 19340 14881
rect 19295 14844 19340 14872
rect 16301 14835 16359 14841
rect 19328 14835 19340 14844
rect 19334 14832 19340 14835
rect 19392 14832 19398 14884
rect 20346 14832 20352 14884
rect 20404 14872 20410 14884
rect 21637 14875 21695 14881
rect 21637 14872 21649 14875
rect 20404 14844 21649 14872
rect 20404 14832 20410 14844
rect 21637 14841 21649 14844
rect 21683 14872 21695 14875
rect 21928 14872 21956 14912
rect 22002 14900 22008 14952
rect 22060 14940 22066 14952
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 22060 14912 22109 14940
rect 22060 14900 22066 14912
rect 22097 14909 22109 14912
rect 22143 14940 22155 14943
rect 23768 14940 23796 14980
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 24268 14980 24313 15008
rect 24268 14968 24274 14980
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 22143 14912 23704 14940
rect 23768 14912 24041 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 22189 14875 22247 14881
rect 22189 14872 22201 14875
rect 21683 14844 21864 14872
rect 21928 14844 22201 14872
rect 21683 14841 21695 14844
rect 21637 14835 21695 14841
rect 13357 14807 13415 14813
rect 13357 14773 13369 14807
rect 13403 14773 13415 14807
rect 14826 14804 14832 14816
rect 14787 14776 14832 14804
rect 13357 14767 13415 14773
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 14921 14807 14979 14813
rect 14921 14773 14933 14807
rect 14967 14804 14979 14807
rect 15102 14804 15108 14816
rect 14967 14776 15108 14804
rect 14967 14773 14979 14776
rect 14921 14767 14979 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 16025 14807 16083 14813
rect 15436 14776 15481 14804
rect 15436 14764 15442 14776
rect 16025 14773 16037 14807
rect 16071 14804 16083 14807
rect 16206 14804 16212 14816
rect 16071 14776 16212 14804
rect 16071 14773 16083 14776
rect 16025 14767 16083 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 17862 14804 17868 14816
rect 17823 14776 17868 14804
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 20438 14804 20444 14816
rect 20399 14776 20444 14804
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 21836 14804 21864 14844
rect 22189 14841 22201 14844
rect 22235 14841 22247 14875
rect 22189 14835 22247 14841
rect 22554 14804 22560 14816
rect 21836 14776 22560 14804
rect 22554 14764 22560 14776
rect 22612 14764 22618 14816
rect 23474 14804 23480 14816
rect 23435 14776 23480 14804
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 23676 14813 23704 14912
rect 24029 14909 24041 14912
rect 24075 14909 24087 14943
rect 26142 14940 26148 14952
rect 26103 14912 26148 14940
rect 24029 14903 24087 14909
rect 26142 14900 26148 14912
rect 26200 14900 26206 14952
rect 24949 14875 25007 14881
rect 24949 14841 24961 14875
rect 24995 14872 25007 14875
rect 25406 14872 25412 14884
rect 24995 14844 25412 14872
rect 24995 14841 25007 14844
rect 24949 14835 25007 14841
rect 25406 14832 25412 14844
rect 25464 14832 25470 14884
rect 26326 14832 26332 14884
rect 26384 14881 26390 14884
rect 26384 14875 26448 14881
rect 26384 14841 26402 14875
rect 26436 14841 26448 14875
rect 26384 14835 26448 14841
rect 26384 14832 26390 14835
rect 23661 14807 23719 14813
rect 23661 14773 23673 14807
rect 23707 14773 23719 14807
rect 23661 14767 23719 14773
rect 24578 14764 24584 14816
rect 24636 14804 24642 14816
rect 25225 14807 25283 14813
rect 25225 14804 25237 14807
rect 24636 14776 25237 14804
rect 24636 14764 24642 14776
rect 25225 14773 25237 14776
rect 25271 14773 25283 14807
rect 27522 14804 27528 14816
rect 27483 14776 27528 14804
rect 25225 14767 25283 14773
rect 27522 14764 27528 14776
rect 27580 14804 27586 14816
rect 28077 14807 28135 14813
rect 28077 14804 28089 14807
rect 27580 14776 28089 14804
rect 27580 14764 27586 14776
rect 28077 14773 28089 14776
rect 28123 14773 28135 14807
rect 28077 14767 28135 14773
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 2498 14560 2504 14612
rect 2556 14600 2562 14612
rect 2869 14603 2927 14609
rect 2869 14600 2881 14603
rect 2556 14572 2881 14600
rect 2556 14560 2562 14572
rect 2869 14569 2881 14572
rect 2915 14600 2927 14603
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 2915 14572 3525 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 3513 14569 3525 14572
rect 3559 14600 3571 14603
rect 3694 14600 3700 14612
rect 3559 14572 3700 14600
rect 3559 14569 3571 14572
rect 3513 14563 3571 14569
rect 3694 14560 3700 14572
rect 3752 14560 3758 14612
rect 4893 14603 4951 14609
rect 4893 14569 4905 14603
rect 4939 14600 4951 14603
rect 4982 14600 4988 14612
rect 4939 14572 4988 14600
rect 4939 14569 4951 14572
rect 4893 14563 4951 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 7190 14600 7196 14612
rect 6880 14572 7196 14600
rect 6880 14560 6886 14572
rect 7190 14560 7196 14572
rect 7248 14600 7254 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 7248 14572 7297 14600
rect 7248 14560 7254 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 7285 14563 7343 14569
rect 8021 14603 8079 14609
rect 8021 14569 8033 14603
rect 8067 14600 8079 14603
rect 10226 14600 10232 14612
rect 8067 14572 10232 14600
rect 8067 14569 8079 14572
rect 8021 14563 8079 14569
rect 10226 14560 10232 14572
rect 10284 14600 10290 14612
rect 10413 14603 10471 14609
rect 10413 14600 10425 14603
rect 10284 14572 10425 14600
rect 10284 14560 10290 14572
rect 10413 14569 10425 14572
rect 10459 14569 10471 14603
rect 11698 14600 11704 14612
rect 11659 14572 11704 14600
rect 10413 14563 10471 14569
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 15378 14560 15384 14612
rect 15436 14600 15442 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 15436 14572 15485 14600
rect 15436 14560 15442 14572
rect 15473 14569 15485 14572
rect 15519 14569 15531 14603
rect 15473 14563 15531 14569
rect 18325 14603 18383 14609
rect 18325 14569 18337 14603
rect 18371 14600 18383 14603
rect 18782 14600 18788 14612
rect 18371 14572 18788 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 20346 14600 20352 14612
rect 20307 14572 20352 14600
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 24029 14603 24087 14609
rect 24029 14569 24041 14603
rect 24075 14600 24087 14603
rect 24118 14600 24124 14612
rect 24075 14572 24124 14600
rect 24075 14569 24087 14572
rect 24029 14563 24087 14569
rect 24118 14560 24124 14572
rect 24176 14560 24182 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 25777 14603 25835 14609
rect 25777 14600 25789 14603
rect 24912 14572 25789 14600
rect 24912 14560 24918 14572
rect 25777 14569 25789 14572
rect 25823 14600 25835 14603
rect 26326 14600 26332 14612
rect 25823 14572 26332 14600
rect 25823 14569 25835 14572
rect 25777 14563 25835 14569
rect 26326 14560 26332 14572
rect 26384 14560 26390 14612
rect 26513 14603 26571 14609
rect 26513 14569 26525 14603
rect 26559 14600 26571 14603
rect 26602 14600 26608 14612
rect 26559 14572 26608 14600
rect 26559 14569 26571 14572
rect 26513 14563 26571 14569
rect 26602 14560 26608 14572
rect 26660 14560 26666 14612
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 1756 14467 1814 14473
rect 1756 14433 1768 14467
rect 1802 14464 1814 14467
rect 2774 14464 2780 14476
rect 1802 14436 2780 14464
rect 1802 14433 1814 14436
rect 1756 14427 1814 14433
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4798 14464 4804 14476
rect 4111 14436 4804 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 5000 14464 5028 14560
rect 5620 14535 5678 14541
rect 5620 14501 5632 14535
rect 5666 14532 5678 14535
rect 5718 14532 5724 14544
rect 5666 14504 5724 14532
rect 5666 14501 5678 14504
rect 5620 14495 5678 14501
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 8481 14535 8539 14541
rect 8481 14501 8493 14535
rect 8527 14532 8539 14535
rect 9214 14532 9220 14544
rect 8527 14504 9220 14532
rect 8527 14501 8539 14504
rect 8481 14495 8539 14501
rect 9214 14492 9220 14504
rect 9272 14532 9278 14544
rect 9582 14532 9588 14544
rect 9272 14504 9588 14532
rect 9272 14492 9278 14504
rect 9582 14492 9588 14504
rect 9640 14492 9646 14544
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 10134 14532 10140 14544
rect 9824 14504 10140 14532
rect 9824 14492 9830 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 16390 14541 16396 14544
rect 16384 14532 16396 14541
rect 16351 14504 16396 14532
rect 16384 14495 16396 14504
rect 16390 14492 16396 14495
rect 16448 14492 16454 14544
rect 19702 14532 19708 14544
rect 19615 14504 19708 14532
rect 19702 14492 19708 14504
rect 19760 14532 19766 14544
rect 20530 14532 20536 14544
rect 19760 14504 20536 14532
rect 19760 14492 19766 14504
rect 20530 14492 20536 14504
rect 20588 14492 20594 14544
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 24397 14535 24455 14541
rect 24397 14532 24409 14535
rect 23716 14504 24409 14532
rect 23716 14492 23722 14504
rect 24397 14501 24409 14504
rect 24443 14532 24455 14535
rect 25130 14532 25136 14544
rect 24443 14504 25136 14532
rect 24443 14501 24455 14504
rect 24397 14495 24455 14501
rect 25130 14492 25136 14504
rect 25188 14492 25194 14544
rect 25498 14532 25504 14544
rect 25459 14504 25504 14532
rect 25498 14492 25504 14504
rect 25556 14492 25562 14544
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 5000 14436 5365 14464
rect 5353 14433 5365 14436
rect 5399 14464 5411 14467
rect 6178 14464 6184 14476
rect 5399 14436 6184 14464
rect 5399 14433 5411 14436
rect 5353 14427 5411 14433
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 9490 14464 9496 14476
rect 8435 14436 9496 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 10686 14464 10692 14476
rect 10551 14436 10692 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10928 14436 11161 14464
rect 10928 14424 10934 14436
rect 11149 14433 11161 14436
rect 11195 14464 11207 14467
rect 11238 14464 11244 14476
rect 11195 14436 11244 14464
rect 11195 14433 11207 14436
rect 11149 14427 11207 14433
rect 11238 14424 11244 14436
rect 11296 14464 11302 14476
rect 12060 14467 12118 14473
rect 12060 14464 12072 14467
rect 11296 14436 12072 14464
rect 11296 14424 11302 14436
rect 12060 14433 12072 14436
rect 12106 14464 12118 14467
rect 13078 14464 13084 14476
rect 12106 14436 13084 14464
rect 12106 14433 12118 14436
rect 12060 14427 12118 14433
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 16206 14464 16212 14476
rect 16163 14436 16212 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 19610 14464 19616 14476
rect 19571 14436 19616 14464
rect 19610 14424 19616 14436
rect 19668 14424 19674 14476
rect 21082 14424 21088 14476
rect 21140 14464 21146 14476
rect 21801 14467 21859 14473
rect 21801 14464 21813 14467
rect 21140 14436 21813 14464
rect 21140 14424 21146 14436
rect 21801 14433 21813 14436
rect 21847 14433 21859 14467
rect 26878 14464 26884 14476
rect 26839 14436 26884 14464
rect 21801 14427 21859 14433
rect 26878 14424 26884 14436
rect 26936 14424 26942 14476
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 8846 14396 8852 14408
rect 8711 14368 8852 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 8846 14356 8852 14368
rect 8904 14396 8910 14408
rect 9858 14396 9864 14408
rect 8904 14368 9864 14396
rect 8904 14356 8910 14368
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10594 14396 10600 14408
rect 10555 14368 10600 14396
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 19886 14396 19892 14408
rect 19847 14368 19892 14396
rect 11793 14359 11851 14365
rect 9030 14328 9036 14340
rect 8991 14300 9036 14328
rect 9030 14288 9036 14300
rect 9088 14288 9094 14340
rect 9950 14288 9956 14340
rect 10008 14328 10014 14340
rect 10045 14331 10103 14337
rect 10045 14328 10057 14331
rect 10008 14300 10057 14328
rect 10008 14288 10014 14300
rect 10045 14297 10057 14300
rect 10091 14297 10103 14331
rect 10045 14291 10103 14297
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4249 14263 4307 14269
rect 4249 14260 4261 14263
rect 4120 14232 4261 14260
rect 4120 14220 4126 14232
rect 4249 14229 4261 14232
rect 4295 14229 4307 14263
rect 4249 14223 4307 14229
rect 5261 14263 5319 14269
rect 5261 14229 5273 14263
rect 5307 14260 5319 14263
rect 5626 14260 5632 14272
rect 5307 14232 5632 14260
rect 5307 14229 5319 14232
rect 5261 14223 5319 14229
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 6730 14260 6736 14272
rect 6691 14232 6736 14260
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 7926 14260 7932 14272
rect 7887 14232 7932 14260
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 9732 14232 9873 14260
rect 9732 14220 9738 14232
rect 9861 14229 9873 14232
rect 9907 14260 9919 14263
rect 11808 14260 11836 14359
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 21545 14399 21603 14405
rect 21545 14396 21557 14399
rect 21508 14368 21557 14396
rect 21508 14356 21514 14368
rect 21545 14365 21557 14368
rect 21591 14365 21603 14399
rect 21545 14359 21603 14365
rect 24026 14356 24032 14408
rect 24084 14396 24090 14408
rect 24489 14399 24547 14405
rect 24489 14396 24501 14399
rect 24084 14368 24501 14396
rect 24084 14356 24090 14368
rect 24489 14365 24501 14368
rect 24535 14365 24547 14399
rect 24489 14359 24547 14365
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14365 24639 14399
rect 26142 14396 26148 14408
rect 24581 14359 24639 14365
rect 25056 14368 26148 14396
rect 19153 14331 19211 14337
rect 19153 14297 19165 14331
rect 19199 14328 19211 14331
rect 19334 14328 19340 14340
rect 19199 14300 19340 14328
rect 19199 14297 19211 14300
rect 19153 14291 19211 14297
rect 19334 14288 19340 14300
rect 19392 14328 19398 14340
rect 24596 14328 24624 14359
rect 19392 14300 19840 14328
rect 19392 14288 19398 14300
rect 19812 14272 19840 14300
rect 23860 14300 24624 14328
rect 11974 14260 11980 14272
rect 9907 14232 11980 14260
rect 9907 14229 9919 14232
rect 9861 14223 9919 14229
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 13817 14263 13875 14269
rect 13817 14229 13829 14263
rect 13863 14260 13875 14263
rect 14826 14260 14832 14272
rect 13863 14232 14832 14260
rect 13863 14229 13875 14232
rect 13817 14223 13875 14229
rect 14826 14220 14832 14232
rect 14884 14260 14890 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14884 14232 15117 14260
rect 14884 14220 14890 14232
rect 15105 14229 15117 14232
rect 15151 14260 15163 14263
rect 15562 14260 15568 14272
rect 15151 14232 15568 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 17494 14260 17500 14272
rect 17455 14232 17500 14260
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 18690 14260 18696 14272
rect 18651 14232 18696 14260
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 19794 14220 19800 14272
rect 19852 14220 19858 14272
rect 21358 14260 21364 14272
rect 21319 14232 21364 14260
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 22554 14220 22560 14272
rect 22612 14260 22618 14272
rect 23860 14269 23888 14300
rect 22925 14263 22983 14269
rect 22925 14260 22937 14263
rect 22612 14232 22937 14260
rect 22612 14220 22618 14232
rect 22925 14229 22937 14232
rect 22971 14260 22983 14263
rect 23845 14263 23903 14269
rect 23845 14260 23857 14263
rect 22971 14232 23857 14260
rect 22971 14229 22983 14232
rect 22925 14223 22983 14229
rect 23845 14229 23857 14232
rect 23891 14229 23903 14263
rect 23845 14223 23903 14229
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 25056 14269 25084 14368
rect 26142 14356 26148 14368
rect 26200 14356 26206 14408
rect 26602 14356 26608 14408
rect 26660 14396 26666 14408
rect 26973 14399 27031 14405
rect 26973 14396 26985 14399
rect 26660 14368 26985 14396
rect 26660 14356 26666 14368
rect 26973 14365 26985 14368
rect 27019 14365 27031 14399
rect 27154 14396 27160 14408
rect 27115 14368 27160 14396
rect 26973 14359 27031 14365
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 25041 14263 25099 14269
rect 25041 14260 25053 14263
rect 24360 14232 25053 14260
rect 24360 14220 24366 14232
rect 25041 14229 25053 14232
rect 25087 14229 25099 14263
rect 25041 14223 25099 14229
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 1857 14059 1915 14065
rect 1857 14025 1869 14059
rect 1903 14056 1915 14059
rect 2130 14056 2136 14068
rect 1903 14028 2136 14056
rect 1903 14025 1915 14028
rect 1857 14019 1915 14025
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 3050 14056 3056 14068
rect 3011 14028 3056 14056
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 3970 14056 3976 14068
rect 3651 14028 3976 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 4798 14056 4804 14068
rect 4755 14028 4804 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 5040 14028 6561 14056
rect 5040 14016 5046 14028
rect 6549 14025 6561 14028
rect 6595 14056 6607 14059
rect 7282 14056 7288 14068
rect 6595 14028 7288 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8662 14056 8668 14068
rect 7984 14028 8668 14056
rect 7984 14016 7990 14028
rect 8662 14016 8668 14028
rect 8720 14056 8726 14068
rect 9769 14059 9827 14065
rect 9769 14056 9781 14059
rect 8720 14028 9781 14056
rect 8720 14016 8726 14028
rect 9769 14025 9781 14028
rect 9815 14025 9827 14059
rect 9769 14019 9827 14025
rect 10413 14059 10471 14065
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 10594 14056 10600 14068
rect 10459 14028 10600 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 2148 13988 2176 14016
rect 3234 13988 3240 14000
rect 2148 13960 3240 13988
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 6822 13988 6828 14000
rect 5592 13960 6828 13988
rect 5592 13948 5598 13960
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2958 13920 2964 13932
rect 2547 13892 2964 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 3936 13892 4261 13920
rect 3936 13880 3942 13892
rect 4249 13889 4261 13892
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4338 13880 4344 13932
rect 4396 13920 4402 13932
rect 4985 13923 5043 13929
rect 4985 13920 4997 13923
rect 4396 13892 4997 13920
rect 4396 13880 4402 13892
rect 4985 13889 4997 13892
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2590 13852 2596 13864
rect 2455 13824 2596 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4154 13852 4160 13864
rect 4111 13824 4160 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 5000 13852 5028 13883
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5132 13892 5825 13920
rect 5132 13880 5138 13892
rect 5813 13889 5825 13892
rect 5859 13920 5871 13923
rect 5994 13920 6000 13932
rect 5859 13892 6000 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 5994 13880 6000 13892
rect 6052 13920 6058 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 6052 13892 7389 13920
rect 6052 13880 6058 13892
rect 7377 13889 7389 13892
rect 7423 13920 7435 13923
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7423 13892 7849 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8297 13923 8355 13929
rect 8297 13920 8309 13923
rect 8168 13892 8309 13920
rect 8168 13880 8174 13892
rect 8297 13889 8309 13892
rect 8343 13920 8355 13923
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 8343 13892 8401 13920
rect 8343 13889 8355 13892
rect 8297 13883 8355 13889
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 6270 13852 6276 13864
rect 5000 13824 5396 13852
rect 6231 13824 6276 13852
rect 5368 13784 5396 13824
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 7190 13852 7196 13864
rect 7151 13824 7196 13852
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7340 13824 7385 13852
rect 7340 13812 7346 13824
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8656 13855 8714 13861
rect 8656 13852 8668 13855
rect 8536 13824 8668 13852
rect 8536 13812 8542 13824
rect 8656 13821 8668 13824
rect 8702 13852 8714 13855
rect 10428 13852 10456 14019
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11238 14056 11244 14068
rect 11199 14028 11244 14056
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 11974 14056 11980 14068
rect 11931 14028 11980 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 14829 14059 14887 14065
rect 14829 14056 14841 14059
rect 14792 14028 14841 14056
rect 14792 14016 14798 14028
rect 14829 14025 14841 14028
rect 14875 14025 14887 14059
rect 14829 14019 14887 14025
rect 15013 14059 15071 14065
rect 15013 14025 15025 14059
rect 15059 14056 15071 14059
rect 15378 14056 15384 14068
rect 15059 14028 15384 14056
rect 15059 14025 15071 14028
rect 15013 14019 15071 14025
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 12492 13960 12537 13988
rect 12492 13948 12498 13960
rect 13078 13920 13084 13932
rect 13039 13892 13084 13920
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 13262 13920 13268 13932
rect 13136 13892 13268 13920
rect 13136 13880 13142 13892
rect 13262 13880 13268 13892
rect 13320 13920 13326 13932
rect 13449 13923 13507 13929
rect 13449 13920 13461 13923
rect 13320 13892 13461 13920
rect 13320 13880 13326 13892
rect 13449 13889 13461 13892
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 10686 13852 10692 13864
rect 8702 13824 10456 13852
rect 10647 13824 10692 13852
rect 8702 13821 8714 13824
rect 8656 13815 8714 13821
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12768 13824 12909 13852
rect 12768 13812 12774 13824
rect 12897 13821 12909 13824
rect 12943 13852 12955 13855
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 12943 13824 13829 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 14844 13852 14872 14019
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 16485 14059 16543 14065
rect 16485 14056 16497 14059
rect 16448 14028 16497 14056
rect 16448 14016 16454 14028
rect 16485 14025 16497 14028
rect 16531 14056 16543 14059
rect 16666 14056 16672 14068
rect 16531 14028 16672 14056
rect 16531 14025 16543 14028
rect 16485 14019 16543 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 17678 14016 17684 14068
rect 17736 14056 17742 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17736 14028 17785 14056
rect 17736 14016 17742 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 17788 13920 17816 14019
rect 18230 14016 18236 14068
rect 18288 14056 18294 14068
rect 18417 14059 18475 14065
rect 18417 14056 18429 14059
rect 18288 14028 18429 14056
rect 18288 14016 18294 14028
rect 18417 14025 18429 14028
rect 18463 14025 18475 14059
rect 18417 14019 18475 14025
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18782 14056 18788 14068
rect 18647 14028 18788 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18432 13988 18460 14019
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19610 14056 19616 14068
rect 19571 14028 19616 14056
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 20165 14059 20223 14065
rect 20165 14025 20177 14059
rect 20211 14056 20223 14059
rect 21358 14056 21364 14068
rect 20211 14028 21364 14056
rect 20211 14025 20223 14028
rect 20165 14019 20223 14025
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 21508 14028 21557 14056
rect 21508 14016 21514 14028
rect 21545 14025 21557 14028
rect 21591 14025 21603 14059
rect 21726 14056 21732 14068
rect 21687 14028 21732 14056
rect 21545 14019 21603 14025
rect 21726 14016 21732 14028
rect 21784 14016 21790 14068
rect 22830 14056 22836 14068
rect 22791 14028 22836 14056
rect 22830 14016 22836 14028
rect 22888 14016 22894 14068
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 23658 14056 23664 14068
rect 23523 14028 23664 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 24026 14056 24032 14068
rect 23987 14028 24032 14056
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 25866 14016 25872 14068
rect 25924 14056 25930 14068
rect 27154 14056 27160 14068
rect 25924 14028 27160 14056
rect 25924 14016 25930 14028
rect 27154 14016 27160 14028
rect 27212 14056 27218 14068
rect 27893 14059 27951 14065
rect 27893 14056 27905 14059
rect 27212 14028 27905 14056
rect 27212 14016 27218 14028
rect 27893 14025 27905 14028
rect 27939 14025 27951 14059
rect 27893 14019 27951 14025
rect 18874 13988 18880 14000
rect 18432 13960 18880 13988
rect 18874 13948 18880 13960
rect 18932 13948 18938 14000
rect 19628 13988 19656 14016
rect 20806 13988 20812 14000
rect 19628 13960 20812 13988
rect 20806 13948 20812 13960
rect 20864 13948 20870 14000
rect 19150 13920 19156 13932
rect 17788 13892 19156 13920
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 20717 13923 20775 13929
rect 20717 13920 20729 13923
rect 20404 13892 20729 13920
rect 20404 13880 20410 13892
rect 20717 13889 20729 13892
rect 20763 13889 20775 13923
rect 21376 13920 21404 14016
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21376 13892 22201 13920
rect 20717 13883 20775 13889
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 22373 13923 22431 13929
rect 22373 13889 22385 13923
rect 22419 13920 22431 13923
rect 22848 13920 22876 14016
rect 26602 13948 26608 14000
rect 26660 13988 26666 14000
rect 28261 13991 28319 13997
rect 28261 13988 28273 13991
rect 26660 13960 28273 13988
rect 26660 13948 26666 13960
rect 28261 13957 28273 13960
rect 28307 13957 28319 13991
rect 28261 13951 28319 13957
rect 26786 13920 26792 13932
rect 22419 13892 22876 13920
rect 26747 13892 26792 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 26786 13880 26792 13892
rect 26844 13920 26850 13932
rect 27341 13923 27399 13929
rect 27341 13920 27353 13923
rect 26844 13892 27353 13920
rect 26844 13880 26850 13892
rect 27341 13889 27353 13892
rect 27387 13889 27399 13923
rect 27522 13920 27528 13932
rect 27483 13892 27528 13920
rect 27341 13883 27399 13889
rect 27522 13880 27528 13892
rect 27580 13920 27586 13932
rect 27706 13920 27712 13932
rect 27580 13892 27712 13920
rect 27580 13880 27586 13892
rect 27706 13880 27712 13892
rect 27764 13880 27770 13932
rect 15470 13852 15476 13864
rect 14844 13824 15476 13852
rect 13817 13815 13875 13821
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13852 16267 13855
rect 16298 13852 16304 13864
rect 16255 13824 16304 13852
rect 16255 13821 16267 13824
rect 16209 13815 16267 13821
rect 16298 13812 16304 13824
rect 16356 13852 16362 13864
rect 16356 13824 16620 13852
rect 16356 13812 16362 13824
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5368 13756 5549 13784
rect 5537 13753 5549 13756
rect 5583 13753 5595 13787
rect 11330 13784 11336 13796
rect 11291 13756 11336 13784
rect 5537 13747 5595 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 16592 13784 16620 13824
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18840 13824 19073 13852
rect 18840 13812 18846 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19610 13812 19616 13864
rect 19668 13852 19674 13864
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19668 13824 20085 13852
rect 19668 13812 19674 13824
rect 20073 13821 20085 13824
rect 20119 13852 20131 13855
rect 20254 13852 20260 13864
rect 20119 13824 20260 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20254 13812 20260 13824
rect 20312 13852 20318 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20312 13824 20637 13852
rect 20312 13812 20318 13824
rect 20625 13821 20637 13824
rect 20671 13852 20683 13855
rect 22738 13852 22744 13864
rect 20671 13824 22744 13852
rect 20671 13821 20683 13824
rect 20625 13815 20683 13821
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 24302 13812 24308 13864
rect 24360 13852 24366 13864
rect 24397 13855 24455 13861
rect 24397 13852 24409 13855
rect 24360 13824 24409 13852
rect 24360 13812 24366 13824
rect 24397 13821 24409 13824
rect 24443 13821 24455 13855
rect 24397 13815 24455 13821
rect 17034 13784 17040 13796
rect 16592 13756 17040 13784
rect 17034 13744 17040 13756
rect 17092 13744 17098 13796
rect 20438 13744 20444 13796
rect 20496 13784 20502 13796
rect 21082 13784 21088 13796
rect 20496 13756 21088 13784
rect 20496 13744 20502 13756
rect 21082 13744 21088 13756
rect 21140 13784 21146 13796
rect 21177 13787 21235 13793
rect 21177 13784 21189 13787
rect 21140 13756 21189 13784
rect 21140 13744 21146 13756
rect 21177 13753 21189 13756
rect 21223 13753 21235 13787
rect 21177 13747 21235 13753
rect 23934 13744 23940 13796
rect 23992 13784 23998 13796
rect 24642 13787 24700 13793
rect 24642 13784 24654 13787
rect 23992 13756 24654 13784
rect 23992 13744 23998 13756
rect 24642 13753 24654 13756
rect 24688 13753 24700 13787
rect 24642 13747 24700 13753
rect 26421 13787 26479 13793
rect 26421 13753 26433 13787
rect 26467 13784 26479 13787
rect 27249 13787 27307 13793
rect 27249 13784 27261 13787
rect 26467 13756 27261 13784
rect 26467 13753 26479 13756
rect 26421 13747 26479 13753
rect 27249 13753 27261 13756
rect 27295 13784 27307 13787
rect 27614 13784 27620 13796
rect 27295 13756 27620 13784
rect 27295 13753 27307 13756
rect 27249 13747 27307 13753
rect 27614 13744 27620 13756
rect 27672 13744 27678 13796
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 2314 13716 2320 13728
rect 2275 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 3329 13719 3387 13725
rect 3329 13716 3341 13719
rect 2832 13688 3341 13716
rect 2832 13676 2838 13688
rect 3329 13685 3341 13688
rect 3375 13685 3387 13719
rect 3970 13716 3976 13728
rect 3931 13688 3976 13716
rect 3329 13679 3387 13685
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 5169 13719 5227 13725
rect 5169 13685 5181 13719
rect 5215 13716 5227 13719
rect 5258 13716 5264 13728
rect 5215 13688 5264 13716
rect 5215 13685 5227 13688
rect 5169 13679 5227 13685
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 12250 13716 12256 13728
rect 5684 13688 5729 13716
rect 12163 13688 12256 13716
rect 5684 13676 5690 13688
rect 12250 13676 12256 13688
rect 12308 13716 12314 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 12308 13688 12817 13716
rect 12308 13676 12314 13688
rect 12805 13685 12817 13688
rect 12851 13716 12863 13719
rect 12986 13716 12992 13728
rect 12851 13688 12992 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 14918 13676 14924 13728
rect 14976 13716 14982 13728
rect 15381 13719 15439 13725
rect 15381 13716 15393 13719
rect 14976 13688 15393 13716
rect 14976 13676 14982 13688
rect 15381 13685 15393 13688
rect 15427 13685 15439 13719
rect 15381 13679 15439 13685
rect 16945 13719 17003 13725
rect 16945 13685 16957 13719
rect 16991 13716 17003 13719
rect 17678 13716 17684 13728
rect 16991 13688 17684 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 17678 13676 17684 13688
rect 17736 13676 17742 13728
rect 18690 13676 18696 13728
rect 18748 13716 18754 13728
rect 18969 13719 19027 13725
rect 18969 13716 18981 13719
rect 18748 13688 18981 13716
rect 18748 13676 18754 13688
rect 18969 13685 18981 13688
rect 19015 13716 19027 13719
rect 19242 13716 19248 13728
rect 19015 13688 19248 13716
rect 19015 13685 19027 13688
rect 18969 13679 19027 13685
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 20530 13716 20536 13728
rect 20491 13688 20536 13716
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 25777 13719 25835 13725
rect 22152 13688 22197 13716
rect 22152 13676 22158 13688
rect 25777 13685 25789 13719
rect 25823 13716 25835 13719
rect 25958 13716 25964 13728
rect 25823 13688 25964 13716
rect 25823 13685 25835 13688
rect 25777 13679 25835 13685
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 26786 13676 26792 13728
rect 26844 13716 26850 13728
rect 26881 13719 26939 13725
rect 26881 13716 26893 13719
rect 26844 13688 26893 13716
rect 26844 13676 26850 13688
rect 26881 13685 26893 13688
rect 26927 13685 26939 13719
rect 26881 13679 26939 13685
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4028 13484 4813 13512
rect 4028 13472 4034 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 4801 13475 4859 13481
rect 5169 13515 5227 13521
rect 5169 13481 5181 13515
rect 5215 13512 5227 13515
rect 5442 13512 5448 13524
rect 5215 13484 5448 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 1664 13447 1722 13453
rect 1664 13413 1676 13447
rect 1710 13444 1722 13447
rect 1854 13444 1860 13456
rect 1710 13416 1860 13444
rect 1710 13413 1722 13416
rect 1664 13407 1722 13413
rect 1854 13404 1860 13416
rect 1912 13444 1918 13456
rect 3694 13444 3700 13456
rect 1912 13416 3700 13444
rect 1912 13404 1918 13416
rect 3694 13404 3700 13416
rect 3752 13404 3758 13456
rect 4816 13444 4844 13475
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5776 13484 5825 13512
rect 5776 13472 5782 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 6178 13512 6184 13524
rect 6139 13484 6184 13512
rect 5813 13475 5871 13481
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 8478 13512 8484 13524
rect 8439 13484 8484 13512
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 8846 13512 8852 13524
rect 8807 13484 8852 13512
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 9214 13512 9220 13524
rect 9175 13484 9220 13512
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 10226 13512 10232 13524
rect 10187 13484 10232 13512
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 12710 13512 12716 13524
rect 12671 13484 12716 13512
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 13078 13512 13084 13524
rect 12991 13484 13084 13512
rect 13078 13472 13084 13484
rect 13136 13512 13142 13524
rect 13722 13512 13728 13524
rect 13136 13484 13728 13512
rect 13136 13472 13142 13484
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14918 13472 14924 13524
rect 14976 13512 14982 13524
rect 15013 13515 15071 13521
rect 15013 13512 15025 13515
rect 14976 13484 15025 13512
rect 14976 13472 14982 13484
rect 15013 13481 15025 13484
rect 15059 13481 15071 13515
rect 15013 13475 15071 13481
rect 15102 13472 15108 13524
rect 15160 13512 15166 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 15160 13484 15761 13512
rect 15160 13472 15166 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19886 13512 19892 13524
rect 19383 13484 19892 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 20346 13512 20352 13524
rect 20259 13484 20352 13512
rect 20346 13472 20352 13484
rect 20404 13512 20410 13524
rect 20530 13512 20536 13524
rect 20404 13484 20536 13512
rect 20404 13472 20410 13484
rect 20530 13472 20536 13484
rect 20588 13512 20594 13524
rect 21726 13512 21732 13524
rect 20588 13484 21732 13512
rect 20588 13472 20594 13484
rect 21726 13472 21732 13484
rect 21784 13472 21790 13524
rect 22094 13472 22100 13524
rect 22152 13512 22158 13524
rect 23201 13515 23259 13521
rect 23201 13512 23213 13515
rect 22152 13484 23213 13512
rect 22152 13472 22158 13484
rect 23201 13481 23213 13484
rect 23247 13481 23259 13515
rect 23201 13475 23259 13481
rect 23845 13515 23903 13521
rect 23845 13481 23857 13515
rect 23891 13512 23903 13515
rect 23934 13512 23940 13524
rect 23891 13484 23940 13512
rect 23891 13481 23903 13484
rect 23845 13475 23903 13481
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 25317 13515 25375 13521
rect 25317 13481 25329 13515
rect 25363 13512 25375 13515
rect 25406 13512 25412 13524
rect 25363 13484 25412 13512
rect 25363 13481 25375 13484
rect 25317 13475 25375 13481
rect 25406 13472 25412 13484
rect 25464 13512 25470 13524
rect 25866 13512 25872 13524
rect 25464 13484 25872 13512
rect 25464 13472 25470 13484
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 26329 13515 26387 13521
rect 26329 13481 26341 13515
rect 26375 13512 26387 13515
rect 26513 13515 26571 13521
rect 26513 13512 26525 13515
rect 26375 13484 26525 13512
rect 26375 13481 26387 13484
rect 26329 13475 26387 13481
rect 26513 13481 26525 13484
rect 26559 13512 26571 13515
rect 26878 13512 26884 13524
rect 26559 13484 26884 13512
rect 26559 13481 26571 13484
rect 26513 13475 26571 13481
rect 26878 13472 26884 13484
rect 26936 13472 26942 13524
rect 26970 13472 26976 13524
rect 27028 13512 27034 13524
rect 27617 13515 27675 13521
rect 27028 13484 27073 13512
rect 27028 13472 27034 13484
rect 27617 13481 27629 13515
rect 27663 13512 27675 13515
rect 27706 13512 27712 13524
rect 27663 13484 27712 13512
rect 27663 13481 27675 13484
rect 27617 13475 27675 13481
rect 27706 13472 27712 13484
rect 27764 13472 27770 13524
rect 5350 13444 5356 13456
rect 4816 13416 5356 13444
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 6454 13404 6460 13456
rect 6512 13444 6518 13456
rect 6632 13447 6690 13453
rect 6632 13444 6644 13447
rect 6512 13416 6644 13444
rect 6512 13404 6518 13416
rect 6632 13413 6644 13416
rect 6678 13444 6690 13447
rect 6730 13444 6736 13456
rect 6678 13416 6736 13444
rect 6678 13413 6690 13416
rect 6632 13407 6690 13413
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 11517 13447 11575 13453
rect 11517 13413 11529 13447
rect 11563 13444 11575 13447
rect 11698 13444 11704 13456
rect 11563 13416 11704 13444
rect 11563 13413 11575 13416
rect 11517 13407 11575 13413
rect 11698 13404 11704 13416
rect 11756 13444 11762 13456
rect 13630 13444 13636 13456
rect 11756 13416 13636 13444
rect 11756 13404 11762 13416
rect 13630 13404 13636 13416
rect 13688 13444 13694 13456
rect 15470 13444 15476 13456
rect 13688 13416 15476 13444
rect 13688 13404 13694 13416
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 17304 13447 17362 13453
rect 17304 13413 17316 13447
rect 17350 13444 17362 13447
rect 17494 13444 17500 13456
rect 17350 13416 17500 13444
rect 17350 13413 17362 13416
rect 17304 13407 17362 13413
rect 17494 13404 17500 13416
rect 17552 13404 17558 13456
rect 19702 13444 19708 13456
rect 19663 13416 19708 13444
rect 19702 13404 19708 13416
rect 19760 13404 19766 13456
rect 21450 13444 21456 13456
rect 21100 13416 21456 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1486 13376 1492 13388
rect 1443 13348 1492 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1486 13336 1492 13348
rect 1544 13376 1550 13388
rect 2498 13376 2504 13388
rect 1544 13348 2504 13376
rect 1544 13336 1550 13348
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 6472 13376 6500 13404
rect 4387 13348 6500 13376
rect 14737 13379 14795 13385
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 15010 13376 15016 13388
rect 14783 13348 15016 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 15010 13336 15016 13348
rect 15068 13376 15074 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15068 13348 15669 13376
rect 15068 13336 15074 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 17034 13376 17040 13388
rect 16995 13348 17040 13376
rect 15657 13339 15715 13345
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 4522 13268 4528 13320
rect 4580 13308 4586 13320
rect 4890 13308 4896 13320
rect 4580 13280 4896 13308
rect 4580 13268 4586 13280
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 5258 13308 5264 13320
rect 5219 13280 5264 13308
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5442 13308 5448 13320
rect 5403 13280 5448 13308
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5902 13308 5908 13320
rect 5776 13280 5908 13308
rect 5776 13268 5782 13280
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 6328 13280 6377 13308
rect 6328 13268 6334 13280
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 6365 13271 6423 13277
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 13170 13308 13176 13320
rect 13131 13280 13176 13308
rect 11701 13271 11759 13277
rect 4709 13243 4767 13249
rect 4709 13209 4721 13243
rect 4755 13240 4767 13243
rect 5994 13240 6000 13252
rect 4755 13212 6000 13240
rect 4755 13209 4767 13212
rect 4709 13203 4767 13209
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 11716 13240 11744 13271
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 13354 13308 13360 13320
rect 13315 13280 13360 13308
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 20346 13308 20352 13320
rect 19843 13280 20352 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 20346 13268 20352 13280
rect 20404 13268 20410 13320
rect 21100 13308 21128 13416
rect 21450 13404 21456 13416
rect 21508 13444 21514 13456
rect 23014 13444 23020 13456
rect 21508 13416 23020 13444
rect 21508 13404 21514 13416
rect 23014 13404 23020 13416
rect 23072 13444 23078 13456
rect 24302 13444 24308 13456
rect 23072 13416 24308 13444
rect 23072 13404 23078 13416
rect 21177 13379 21235 13385
rect 21177 13345 21189 13379
rect 21223 13376 21235 13379
rect 21536 13379 21594 13385
rect 21536 13376 21548 13379
rect 21223 13348 21548 13376
rect 21223 13345 21235 13348
rect 21177 13339 21235 13345
rect 21536 13345 21548 13348
rect 21582 13376 21594 13379
rect 21910 13376 21916 13388
rect 21582 13348 21916 13376
rect 21582 13345 21594 13348
rect 21536 13339 21594 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 23952 13385 23980 13416
rect 24302 13404 24308 13416
rect 24360 13404 24366 13456
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13345 23995 13379
rect 24204 13379 24262 13385
rect 24204 13376 24216 13379
rect 23937 13339 23995 13345
rect 24044 13348 24216 13376
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 21100 13280 21281 13308
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 21269 13271 21327 13277
rect 23750 13268 23756 13320
rect 23808 13308 23814 13320
rect 24044 13308 24072 13348
rect 24204 13345 24216 13348
rect 24250 13376 24262 13379
rect 26878 13376 26884 13388
rect 24250 13348 26004 13376
rect 26839 13348 26884 13376
rect 24250 13345 24262 13348
rect 24204 13339 24262 13345
rect 25976 13320 26004 13348
rect 26878 13336 26884 13348
rect 26936 13336 26942 13388
rect 23808 13280 24072 13308
rect 23808 13268 23814 13280
rect 25958 13268 25964 13320
rect 26016 13308 26022 13320
rect 27062 13308 27068 13320
rect 26016 13280 27068 13308
rect 26016 13268 26022 13280
rect 27062 13268 27068 13280
rect 27120 13268 27126 13320
rect 15286 13240 15292 13252
rect 11072 13212 11744 13240
rect 15247 13212 15292 13240
rect 11072 13184 11100 13212
rect 15286 13200 15292 13212
rect 15344 13200 15350 13252
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 2832 13144 2877 13172
rect 2832 13132 2838 13144
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 3329 13175 3387 13181
rect 3329 13172 3341 13175
rect 3016 13144 3341 13172
rect 3016 13132 3022 13144
rect 3329 13141 3341 13144
rect 3375 13141 3387 13175
rect 3329 13135 3387 13141
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 5258 13172 5264 13184
rect 4672 13144 5264 13172
rect 4672 13132 4678 13144
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 7282 13132 7288 13184
rect 7340 13172 7346 13184
rect 7745 13175 7803 13181
rect 7745 13172 7757 13175
rect 7340 13144 7757 13172
rect 7340 13132 7346 13144
rect 7745 13141 7757 13144
rect 7791 13141 7803 13175
rect 9950 13172 9956 13184
rect 9911 13144 9956 13172
rect 7745 13135 7803 13141
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 11054 13172 11060 13184
rect 11015 13144 11060 13172
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11149 13175 11207 13181
rect 11149 13141 11161 13175
rect 11195 13172 11207 13175
rect 11422 13172 11428 13184
rect 11195 13144 11428 13172
rect 11195 13141 11207 13144
rect 11149 13135 11207 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12802 13172 12808 13184
rect 12575 13144 12808 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 16942 13172 16948 13184
rect 13044 13144 16948 13172
rect 13044 13132 13050 13144
rect 16942 13132 16948 13144
rect 17000 13172 17006 13184
rect 17310 13172 17316 13184
rect 17000 13144 17316 13172
rect 17000 13132 17006 13144
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 18414 13172 18420 13184
rect 18375 13144 18420 13172
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 20990 13132 20996 13184
rect 21048 13172 21054 13184
rect 22649 13175 22707 13181
rect 22649 13172 22661 13175
rect 21048 13144 22661 13172
rect 21048 13132 21054 13144
rect 22649 13141 22661 13144
rect 22695 13141 22707 13175
rect 22649 13135 22707 13141
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 2041 12971 2099 12977
rect 2041 12937 2053 12971
rect 2087 12968 2099 12971
rect 2866 12968 2872 12980
rect 2087 12940 2872 12968
rect 2087 12937 2099 12940
rect 2041 12931 2099 12937
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2056 12764 2084 12931
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 3694 12928 3700 12980
rect 3752 12968 3758 12980
rect 4065 12971 4123 12977
rect 4065 12968 4077 12971
rect 3752 12940 4077 12968
rect 3752 12928 3758 12940
rect 4065 12937 4077 12940
rect 4111 12937 4123 12971
rect 4065 12931 4123 12937
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5166 12968 5172 12980
rect 4755 12940 5172 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5166 12928 5172 12940
rect 5224 12968 5230 12980
rect 5442 12968 5448 12980
rect 5224 12940 5448 12968
rect 5224 12928 5230 12940
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 6328 12940 6377 12968
rect 6328 12928 6334 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 8294 12968 8300 12980
rect 8255 12940 8300 12968
rect 6365 12931 6423 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 9674 12968 9680 12980
rect 9635 12940 9680 12968
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 11112 12940 11253 12968
rect 11112 12928 11118 12940
rect 11241 12937 11253 12940
rect 11287 12968 11299 12971
rect 11514 12968 11520 12980
rect 11287 12940 11520 12968
rect 11287 12937 11299 12940
rect 11241 12931 11299 12937
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13446 12968 13452 12980
rect 13228 12940 13452 12968
rect 13228 12928 13234 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 14608 12940 14841 12968
rect 14608 12928 14614 12940
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 15010 12968 15016 12980
rect 14971 12940 15016 12968
rect 14829 12931 14887 12937
rect 2498 12900 2504 12912
rect 2459 12872 2504 12900
rect 2498 12860 2504 12872
rect 2556 12900 2562 12912
rect 2556 12872 2728 12900
rect 2556 12860 2562 12872
rect 2700 12841 2728 12872
rect 8478 12860 8484 12912
rect 8536 12900 8542 12912
rect 9692 12900 9720 12928
rect 8536 12872 9720 12900
rect 8536 12860 8542 12872
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6454 12832 6460 12844
rect 5859 12804 6460 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7561 12835 7619 12841
rect 7561 12832 7573 12835
rect 7432 12804 7573 12832
rect 7432 12792 7438 12804
rect 7561 12801 7573 12804
rect 7607 12832 7619 12835
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 7607 12804 7941 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 7929 12801 7941 12804
rect 7975 12801 7987 12835
rect 9692 12832 9720 12872
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9692 12804 9873 12832
rect 7929 12795 7987 12801
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 2958 12773 2964 12776
rect 2952 12764 2964 12773
rect 1443 12736 2084 12764
rect 2919 12736 2964 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2952 12727 2964 12736
rect 2958 12724 2964 12727
rect 3016 12724 3022 12776
rect 7650 12764 7656 12776
rect 6748 12736 7656 12764
rect 1210 12656 1216 12708
rect 1268 12696 1274 12708
rect 5629 12699 5687 12705
rect 5629 12696 5641 12699
rect 1268 12668 2636 12696
rect 1268 12656 1274 12668
rect 1486 12588 1492 12640
rect 1544 12628 1550 12640
rect 1581 12631 1639 12637
rect 1581 12628 1593 12631
rect 1544 12600 1593 12628
rect 1544 12588 1550 12600
rect 1581 12597 1593 12600
rect 1627 12597 1639 12631
rect 2608 12628 2636 12668
rect 5000 12668 5641 12696
rect 5000 12637 5028 12668
rect 5629 12665 5641 12668
rect 5675 12696 5687 12699
rect 6546 12696 6552 12708
rect 5675 12668 6552 12696
rect 5675 12665 5687 12668
rect 5629 12659 5687 12665
rect 6546 12656 6552 12668
rect 6604 12656 6610 12708
rect 4985 12631 5043 12637
rect 4985 12628 4997 12631
rect 2608 12600 4997 12628
rect 1581 12591 1639 12597
rect 4985 12597 4997 12600
rect 5031 12597 5043 12631
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 4985 12591 5043 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 5442 12588 5448 12640
rect 5500 12628 5506 12640
rect 5537 12631 5595 12637
rect 5537 12628 5549 12631
rect 5500 12600 5549 12628
rect 5500 12588 5506 12600
rect 5537 12597 5549 12600
rect 5583 12628 5595 12631
rect 6748 12628 6776 12736
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 7791 12736 8953 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 7285 12699 7343 12705
rect 6880 12668 7052 12696
rect 6880 12656 6886 12668
rect 6914 12628 6920 12640
rect 5583 12600 6776 12628
rect 6875 12600 6920 12628
rect 5583 12597 5595 12600
rect 5537 12591 5595 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7024 12628 7052 12668
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 8662 12696 8668 12708
rect 7331 12668 8668 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 8662 12656 8668 12668
rect 8720 12696 8726 12708
rect 9309 12699 9367 12705
rect 9309 12696 9321 12699
rect 8720 12668 9321 12696
rect 8720 12656 8726 12668
rect 9309 12665 9321 12668
rect 9355 12665 9367 12699
rect 9876 12696 9904 12795
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 11572 12804 13093 12832
rect 11572 12792 11578 12804
rect 13081 12801 13093 12804
rect 13127 12832 13139 12835
rect 13354 12832 13360 12844
rect 13127 12804 13360 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13354 12792 13360 12804
rect 13412 12832 13418 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13412 12804 13921 12832
rect 13412 12792 13418 12804
rect 13909 12801 13921 12804
rect 13955 12832 13967 12835
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13955 12804 14197 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10117 12767 10175 12773
rect 10117 12764 10129 12767
rect 10008 12736 10129 12764
rect 10008 12724 10014 12736
rect 10117 12733 10129 12736
rect 10163 12733 10175 12767
rect 10117 12727 10175 12733
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12618 12764 12624 12776
rect 12299 12736 12624 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12618 12724 12624 12736
rect 12676 12724 12682 12776
rect 12802 12764 12808 12776
rect 12763 12736 12808 12764
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 10870 12696 10876 12708
rect 9876 12668 10876 12696
rect 9309 12659 9367 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 12636 12696 12664 12724
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 12636 12668 12909 12696
rect 12897 12665 12909 12668
rect 12943 12665 12955 12699
rect 14844 12696 14872 12931
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15896 12940 16037 12968
rect 15896 12928 15902 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 17126 12968 17132 12980
rect 17087 12940 17132 12968
rect 16025 12931 16083 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 17494 12968 17500 12980
rect 17455 12940 17500 12968
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18601 12971 18659 12977
rect 18601 12968 18613 12971
rect 18012 12940 18613 12968
rect 18012 12928 18018 12940
rect 18601 12937 18613 12940
rect 18647 12937 18659 12971
rect 18601 12931 18659 12937
rect 20441 12971 20499 12977
rect 20441 12937 20453 12971
rect 20487 12968 20499 12971
rect 20622 12968 20628 12980
rect 20487 12940 20628 12968
rect 20487 12937 20499 12940
rect 20441 12931 20499 12937
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 21729 12971 21787 12977
rect 21729 12968 21741 12971
rect 20864 12940 21741 12968
rect 20864 12928 20870 12940
rect 21729 12937 21741 12940
rect 21775 12968 21787 12971
rect 21821 12971 21879 12977
rect 21821 12968 21833 12971
rect 21775 12940 21833 12968
rect 21775 12937 21787 12940
rect 21729 12931 21787 12937
rect 21821 12937 21833 12940
rect 21867 12937 21879 12971
rect 21821 12931 21879 12937
rect 22005 12971 22063 12977
rect 22005 12937 22017 12971
rect 22051 12968 22063 12971
rect 22094 12968 22100 12980
rect 22051 12940 22100 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 23014 12968 23020 12980
rect 22975 12940 23020 12968
rect 23014 12928 23020 12940
rect 23072 12968 23078 12980
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23072 12940 23857 12968
rect 23072 12928 23078 12940
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 24213 12971 24271 12977
rect 24213 12937 24225 12971
rect 24259 12968 24271 12971
rect 25314 12968 25320 12980
rect 24259 12940 25320 12968
rect 24259 12937 24271 12940
rect 24213 12931 24271 12937
rect 23477 12903 23535 12909
rect 23477 12869 23489 12903
rect 23523 12900 23535 12903
rect 23750 12900 23756 12912
rect 23523 12872 23756 12900
rect 23523 12869 23535 12872
rect 23477 12863 23535 12869
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 15252 12804 15485 12832
rect 15252 12792 15258 12804
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 15657 12835 15715 12841
rect 15657 12801 15669 12835
rect 15703 12832 15715 12835
rect 15746 12832 15752 12844
rect 15703 12804 15752 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 15672 12764 15700 12795
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 17034 12792 17040 12844
rect 17092 12832 17098 12844
rect 17773 12835 17831 12841
rect 17773 12832 17785 12835
rect 17092 12804 17785 12832
rect 17092 12792 17098 12804
rect 17773 12801 17785 12804
rect 17819 12832 17831 12835
rect 19150 12832 19156 12844
rect 17819 12804 19012 12832
rect 19111 12804 19156 12832
rect 17819 12801 17831 12804
rect 17773 12795 17831 12801
rect 15068 12736 15700 12764
rect 15068 12724 15074 12736
rect 16482 12724 16488 12776
rect 16540 12724 16546 12776
rect 18984 12773 19012 12804
rect 19150 12792 19156 12804
rect 19208 12832 19214 12844
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19208 12804 19625 12832
rect 19208 12792 19214 12804
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12832 20407 12835
rect 20438 12832 20444 12844
rect 20395 12804 20444 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 20438 12792 20444 12804
rect 20496 12832 20502 12844
rect 20990 12832 20996 12844
rect 20496 12804 20996 12832
rect 20496 12792 20502 12804
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 22554 12832 22560 12844
rect 22515 12804 22560 12832
rect 22554 12792 22560 12804
rect 22612 12792 22618 12844
rect 18969 12767 19027 12773
rect 18969 12733 18981 12767
rect 19015 12764 19027 12767
rect 19015 12736 20760 12764
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 15381 12699 15439 12705
rect 15381 12696 15393 12699
rect 14844 12668 15393 12696
rect 12897 12659 12955 12665
rect 15381 12665 15393 12668
rect 15427 12696 15439 12699
rect 16500 12696 16528 12724
rect 15427 12668 16528 12696
rect 15427 12665 15439 12668
rect 15381 12659 15439 12665
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 17828 12668 18521 12696
rect 17828 12656 17834 12668
rect 18509 12665 18521 12668
rect 18555 12696 18567 12699
rect 19058 12696 19064 12708
rect 18555 12668 19064 12696
rect 18555 12665 18567 12668
rect 18509 12659 18567 12665
rect 19058 12656 19064 12668
rect 19116 12656 19122 12708
rect 20732 12696 20760 12736
rect 20806 12724 20812 12776
rect 20864 12764 20870 12776
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 20864 12736 20913 12764
rect 20864 12724 20870 12736
rect 20901 12733 20913 12736
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 21545 12767 21603 12773
rect 21545 12733 21557 12767
rect 21591 12764 21603 12767
rect 22186 12764 22192 12776
rect 21591 12736 22192 12764
rect 21591 12733 21603 12736
rect 21545 12727 21603 12733
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 21634 12696 21640 12708
rect 20732 12668 21640 12696
rect 21634 12656 21640 12668
rect 21692 12656 21698 12708
rect 21729 12699 21787 12705
rect 21729 12665 21741 12699
rect 21775 12696 21787 12699
rect 21775 12668 22508 12696
rect 21775 12665 21787 12668
rect 21729 12659 21787 12665
rect 22480 12640 22508 12668
rect 23658 12656 23664 12708
rect 23716 12696 23722 12708
rect 23860 12696 23888 12931
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 26878 12928 26884 12980
rect 26936 12968 26942 12980
rect 28077 12971 28135 12977
rect 28077 12968 28089 12971
rect 26936 12940 28089 12968
rect 26936 12928 26942 12940
rect 28077 12937 28089 12940
rect 28123 12937 28135 12971
rect 28077 12931 28135 12937
rect 24026 12860 24032 12912
rect 24084 12900 24090 12912
rect 24581 12903 24639 12909
rect 24581 12900 24593 12903
rect 24084 12872 24593 12900
rect 24084 12860 24090 12872
rect 24581 12869 24593 12872
rect 24627 12869 24639 12903
rect 24581 12863 24639 12869
rect 26970 12860 26976 12912
rect 27028 12900 27034 12912
rect 27433 12903 27491 12909
rect 27433 12900 27445 12903
rect 27028 12872 27445 12900
rect 27028 12860 27034 12872
rect 27433 12869 27445 12872
rect 27479 12869 27491 12903
rect 27433 12863 27491 12869
rect 24044 12773 24072 12860
rect 27062 12832 27068 12844
rect 27023 12804 27068 12832
rect 27062 12792 27068 12804
rect 27120 12792 27126 12844
rect 27614 12832 27620 12844
rect 27575 12804 27620 12832
rect 27614 12792 27620 12804
rect 27672 12792 27678 12844
rect 25406 12773 25412 12776
rect 24029 12767 24087 12773
rect 24029 12733 24041 12767
rect 24075 12733 24087 12767
rect 24029 12727 24087 12733
rect 25133 12767 25191 12773
rect 25133 12733 25145 12767
rect 25179 12733 25191 12767
rect 25400 12764 25412 12773
rect 25367 12736 25412 12764
rect 25133 12727 25191 12733
rect 25400 12727 25412 12736
rect 24949 12699 25007 12705
rect 24949 12696 24961 12699
rect 23716 12668 24961 12696
rect 23716 12656 23722 12668
rect 24949 12665 24961 12668
rect 24995 12696 25007 12699
rect 25148 12696 25176 12727
rect 25406 12724 25412 12727
rect 25464 12724 25470 12776
rect 25682 12696 25688 12708
rect 24995 12668 25688 12696
rect 24995 12665 25007 12668
rect 24949 12659 25007 12665
rect 25682 12656 25688 12668
rect 25740 12656 25746 12708
rect 7377 12631 7435 12637
rect 7377 12628 7389 12631
rect 7024 12600 7389 12628
rect 7377 12597 7389 12600
rect 7423 12628 7435 12631
rect 7745 12631 7803 12637
rect 7745 12628 7757 12631
rect 7423 12600 7757 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7745 12597 7757 12600
rect 7791 12597 7803 12631
rect 7745 12591 7803 12597
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 8481 12631 8539 12637
rect 8481 12628 8493 12631
rect 8352 12600 8493 12628
rect 8352 12588 8358 12600
rect 8481 12597 8493 12600
rect 8527 12597 8539 12631
rect 8481 12591 8539 12597
rect 10778 12588 10784 12640
rect 10836 12628 10842 12640
rect 11606 12628 11612 12640
rect 10836 12600 11612 12628
rect 10836 12588 10842 12600
rect 11606 12588 11612 12600
rect 11664 12628 11670 12640
rect 11793 12631 11851 12637
rect 11793 12628 11805 12631
rect 11664 12600 11805 12628
rect 11664 12588 11670 12600
rect 11793 12597 11805 12600
rect 11839 12597 11851 12631
rect 12434 12628 12440 12640
rect 12395 12600 12440 12628
rect 11793 12591 11851 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 16482 12628 16488 12640
rect 16443 12600 16488 12628
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 20809 12631 20867 12637
rect 20809 12628 20821 12631
rect 20772 12600 20821 12628
rect 20772 12588 20778 12600
rect 20809 12597 20821 12600
rect 20855 12628 20867 12631
rect 21266 12628 21272 12640
rect 20855 12600 21272 12628
rect 20855 12597 20867 12600
rect 20809 12591 20867 12597
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 22186 12588 22192 12640
rect 22244 12628 22250 12640
rect 22373 12631 22431 12637
rect 22373 12628 22385 12631
rect 22244 12600 22385 12628
rect 22244 12588 22250 12600
rect 22373 12597 22385 12600
rect 22419 12597 22431 12631
rect 22373 12591 22431 12597
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22520 12600 22565 12628
rect 22520 12588 22526 12600
rect 26418 12588 26424 12640
rect 26476 12628 26482 12640
rect 26513 12631 26571 12637
rect 26513 12628 26525 12631
rect 26476 12600 26525 12628
rect 26476 12588 26482 12600
rect 26513 12597 26525 12600
rect 26559 12597 26571 12631
rect 26513 12591 26571 12597
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 2498 12424 2504 12436
rect 1719 12396 2504 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 2498 12384 2504 12396
rect 2556 12384 2562 12436
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 3697 12427 3755 12433
rect 3697 12424 3709 12427
rect 3016 12396 3709 12424
rect 3016 12384 3022 12396
rect 3697 12393 3709 12396
rect 3743 12424 3755 12427
rect 4798 12424 4804 12436
rect 3743 12396 4804 12424
rect 3743 12393 3755 12396
rect 3697 12387 3755 12393
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 6362 12424 6368 12436
rect 5920 12396 6368 12424
rect 2222 12316 2228 12368
rect 2280 12356 2286 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2280 12328 2789 12356
rect 2280 12316 2286 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 2777 12319 2835 12325
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 5074 12356 5080 12368
rect 3292 12328 5080 12356
rect 3292 12316 3298 12328
rect 5074 12316 5080 12328
rect 5132 12356 5138 12368
rect 5169 12359 5227 12365
rect 5169 12356 5181 12359
rect 5132 12328 5181 12356
rect 5132 12316 5138 12328
rect 5169 12325 5181 12328
rect 5215 12356 5227 12359
rect 5442 12356 5448 12368
rect 5215 12328 5448 12356
rect 5215 12325 5227 12328
rect 5169 12319 5227 12325
rect 5442 12316 5448 12328
rect 5500 12316 5506 12368
rect 5920 12300 5948 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 7101 12427 7159 12433
rect 7101 12393 7113 12427
rect 7147 12424 7159 12427
rect 7834 12424 7840 12436
rect 7147 12396 7840 12424
rect 7147 12393 7159 12396
rect 7101 12387 7159 12393
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12424 9827 12427
rect 10686 12424 10692 12436
rect 9815 12396 10692 12424
rect 9815 12393 9827 12396
rect 9769 12387 9827 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 12710 12424 12716 12436
rect 12623 12396 12716 12424
rect 12710 12384 12716 12396
rect 12768 12424 12774 12436
rect 13262 12424 13268 12436
rect 12768 12396 13268 12424
rect 12768 12384 12774 12396
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 15010 12424 15016 12436
rect 14971 12396 15016 12424
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15473 12427 15531 12433
rect 15473 12424 15485 12427
rect 15252 12396 15485 12424
rect 15252 12384 15258 12396
rect 15473 12393 15485 12396
rect 15519 12393 15531 12427
rect 15473 12387 15531 12393
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 16298 12424 16304 12436
rect 15620 12396 16304 12424
rect 15620 12384 15626 12396
rect 16298 12384 16304 12396
rect 16356 12424 16362 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 16356 12396 16773 12424
rect 16356 12384 16362 12396
rect 16761 12393 16773 12396
rect 16807 12424 16819 12427
rect 17770 12424 17776 12436
rect 16807 12396 17776 12424
rect 16807 12393 16819 12396
rect 16761 12387 16819 12393
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 21910 12384 21916 12436
rect 21968 12424 21974 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 21968 12396 22293 12424
rect 21968 12384 21974 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 22281 12387 22339 12393
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 22612 12396 22845 12424
rect 22612 12384 22618 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 24670 12424 24676 12436
rect 24631 12396 24676 12424
rect 22833 12387 22891 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 25406 12384 25412 12436
rect 25464 12424 25470 12436
rect 25685 12427 25743 12433
rect 25685 12424 25697 12427
rect 25464 12396 25697 12424
rect 25464 12384 25470 12396
rect 25685 12393 25697 12396
rect 25731 12393 25743 12427
rect 25685 12387 25743 12393
rect 7006 12316 7012 12368
rect 7064 12356 7070 12368
rect 8113 12359 8171 12365
rect 8113 12356 8125 12359
rect 7064 12328 8125 12356
rect 7064 12316 7070 12328
rect 8113 12325 8125 12328
rect 8159 12325 8171 12359
rect 8113 12319 8171 12325
rect 11514 12316 11520 12368
rect 11572 12365 11578 12368
rect 11572 12359 11636 12365
rect 11572 12325 11590 12359
rect 11624 12325 11636 12359
rect 11572 12319 11636 12325
rect 14737 12359 14795 12365
rect 14737 12325 14749 12359
rect 14783 12356 14795 12359
rect 15102 12356 15108 12368
rect 14783 12328 15108 12356
rect 14783 12325 14795 12328
rect 14737 12319 14795 12325
rect 11572 12316 11578 12319
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 18132 12359 18190 12365
rect 18132 12325 18144 12359
rect 18178 12356 18190 12359
rect 18414 12356 18420 12368
rect 18178 12328 18420 12356
rect 18178 12325 18190 12328
rect 18132 12319 18190 12325
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 21450 12356 21456 12368
rect 20916 12328 21456 12356
rect 20916 12300 20944 12328
rect 21450 12316 21456 12328
rect 21508 12316 21514 12368
rect 25041 12359 25099 12365
rect 25041 12325 25053 12359
rect 25087 12356 25099 12359
rect 25590 12356 25596 12368
rect 25087 12328 25596 12356
rect 25087 12325 25099 12328
rect 25041 12319 25099 12325
rect 25590 12316 25596 12328
rect 25648 12316 25654 12368
rect 26694 12316 26700 12368
rect 26752 12356 26758 12368
rect 27430 12356 27436 12368
rect 26752 12328 27436 12356
rect 26752 12316 26758 12328
rect 27430 12316 27436 12328
rect 27488 12316 27494 12368
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2685 12291 2743 12297
rect 2685 12288 2697 12291
rect 2179 12260 2697 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2685 12257 2697 12260
rect 2731 12288 2743 12291
rect 2866 12288 2872 12300
rect 2731 12260 2872 12288
rect 2731 12257 2743 12260
rect 2685 12251 2743 12257
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3660 12260 4077 12288
rect 3660 12248 3666 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 5902 12288 5908 12300
rect 5863 12260 5908 12288
rect 4065 12251 4123 12257
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 6638 12288 6644 12300
rect 6420 12260 6644 12288
rect 6420 12248 6426 12260
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7156 12260 7481 12288
rect 7156 12248 7162 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12288 7619 12291
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 7607 12260 9413 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 10134 12288 10140 12300
rect 10047 12260 10140 12288
rect 9401 12251 9459 12257
rect 2958 12220 2964 12232
rect 2871 12192 2964 12220
rect 2958 12180 2964 12192
rect 3016 12220 3022 12232
rect 3016 12192 3464 12220
rect 3016 12180 3022 12192
rect 3436 12161 3464 12192
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5810 12220 5816 12232
rect 5684 12192 5816 12220
rect 5684 12180 5690 12192
rect 5810 12180 5816 12192
rect 5868 12220 5874 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5868 12192 6009 12220
rect 5868 12180 5874 12192
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6454 12220 6460 12232
rect 6227 12192 6460 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7576 12220 7604 12251
rect 10134 12248 10140 12260
rect 10192 12288 10198 12300
rect 10502 12288 10508 12300
rect 10192 12260 10508 12288
rect 10192 12248 10198 12260
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 11330 12288 11336 12300
rect 10928 12260 11336 12288
rect 10928 12248 10934 12260
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 16669 12291 16727 12297
rect 16669 12288 16681 12291
rect 15528 12260 16681 12288
rect 15528 12248 15534 12260
rect 16669 12257 16681 12260
rect 16715 12288 16727 12291
rect 17034 12288 17040 12300
rect 16715 12260 17040 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17184 12260 17877 12288
rect 17184 12248 17190 12260
rect 17865 12257 17877 12260
rect 17911 12288 17923 12291
rect 17954 12288 17960 12300
rect 17911 12260 17960 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 20898 12288 20904 12300
rect 20811 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 21174 12297 21180 12300
rect 21168 12288 21180 12297
rect 21135 12260 21180 12288
rect 21168 12251 21180 12260
rect 21174 12248 21180 12251
rect 21232 12248 21238 12300
rect 23566 12288 23572 12300
rect 23527 12260 23572 12288
rect 23566 12248 23572 12260
rect 23624 12248 23630 12300
rect 24118 12288 24124 12300
rect 24079 12260 24124 12288
rect 24118 12248 24124 12260
rect 24176 12248 24182 12300
rect 25866 12288 25872 12300
rect 25332 12260 25872 12288
rect 7742 12220 7748 12232
rect 6972 12192 7604 12220
rect 7703 12192 7748 12220
rect 6972 12180 6978 12192
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12189 10379 12223
rect 16942 12220 16948 12232
rect 16903 12192 16948 12220
rect 10321 12183 10379 12189
rect 3421 12155 3479 12161
rect 3421 12121 3433 12155
rect 3467 12152 3479 12155
rect 5537 12155 5595 12161
rect 3467 12124 4752 12152
rect 3467 12121 3479 12124
rect 3421 12115 3479 12121
rect 4724 12096 4752 12124
rect 5537 12121 5549 12155
rect 5583 12152 5595 12155
rect 6730 12152 6736 12164
rect 5583 12124 6736 12152
rect 5583 12121 5595 12124
rect 5537 12115 5595 12121
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10336 12152 10364 12183
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 24946 12180 24952 12232
rect 25004 12220 25010 12232
rect 25130 12220 25136 12232
rect 25004 12192 25136 12220
rect 25004 12180 25010 12192
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 25332 12229 25360 12260
rect 25866 12248 25872 12260
rect 25924 12248 25930 12300
rect 26878 12288 26884 12300
rect 26839 12260 26884 12288
rect 26878 12248 26884 12260
rect 26936 12248 26942 12300
rect 25317 12223 25375 12229
rect 25317 12189 25329 12223
rect 25363 12189 25375 12223
rect 25317 12183 25375 12189
rect 25498 12180 25504 12232
rect 25556 12220 25562 12232
rect 26602 12220 26608 12232
rect 25556 12192 26608 12220
rect 25556 12180 25562 12192
rect 26602 12180 26608 12192
rect 26660 12220 26666 12232
rect 26973 12223 27031 12229
rect 26973 12220 26985 12223
rect 26660 12192 26985 12220
rect 26660 12180 26666 12192
rect 26973 12189 26985 12192
rect 27019 12189 27031 12223
rect 27154 12220 27160 12232
rect 27115 12192 27160 12220
rect 26973 12183 27031 12189
rect 27154 12180 27160 12192
rect 27212 12180 27218 12232
rect 10594 12152 10600 12164
rect 9916 12124 10600 12152
rect 9916 12112 9922 12124
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 15746 12112 15752 12164
rect 15804 12152 15810 12164
rect 16301 12155 16359 12161
rect 16301 12152 16313 12155
rect 15804 12124 16313 12152
rect 15804 12112 15810 12124
rect 16301 12121 16313 12124
rect 16347 12121 16359 12155
rect 16301 12115 16359 12121
rect 26237 12155 26295 12161
rect 26237 12121 26249 12155
rect 26283 12152 26295 12155
rect 26418 12152 26424 12164
rect 26283 12124 26424 12152
rect 26283 12121 26295 12124
rect 26237 12115 26295 12121
rect 26418 12112 26424 12124
rect 26476 12152 26482 12164
rect 27172 12152 27200 12180
rect 26476 12124 27200 12152
rect 26476 12112 26482 12124
rect 2314 12084 2320 12096
rect 2275 12056 2320 12084
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 4246 12084 4252 12096
rect 4207 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4706 12084 4712 12096
rect 4667 12056 4712 12084
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 6638 12084 6644 12096
rect 6512 12056 6644 12084
rect 6512 12044 6518 12056
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 7009 12087 7067 12093
rect 7009 12053 7021 12087
rect 7055 12084 7067 12087
rect 7374 12084 7380 12096
rect 7055 12056 7380 12084
rect 7055 12053 7067 12056
rect 7009 12047 7067 12053
rect 7374 12044 7380 12056
rect 7432 12084 7438 12096
rect 7650 12084 7656 12096
rect 7432 12056 7656 12084
rect 7432 12044 7438 12056
rect 7650 12044 7656 12056
rect 7708 12084 7714 12096
rect 8665 12087 8723 12093
rect 8665 12084 8677 12087
rect 7708 12056 8677 12084
rect 7708 12044 7714 12056
rect 8665 12053 8677 12056
rect 8711 12084 8723 12087
rect 8754 12084 8760 12096
rect 8711 12056 8760 12084
rect 8711 12053 8723 12056
rect 8665 12047 8723 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 9030 12084 9036 12096
rect 8991 12056 9036 12084
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10686 12084 10692 12096
rect 10376 12056 10692 12084
rect 10376 12044 10382 12056
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10836 12056 11161 12084
rect 10836 12044 10842 12056
rect 11149 12053 11161 12056
rect 11195 12084 11207 12087
rect 11698 12084 11704 12096
rect 11195 12056 11704 12084
rect 11195 12053 11207 12056
rect 11149 12047 11207 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13136 12056 13277 12084
rect 13136 12044 13142 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 15838 12044 15844 12096
rect 15896 12084 15902 12096
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 15896 12056 16129 12084
rect 15896 12044 15902 12056
rect 16117 12053 16129 12056
rect 16163 12053 16175 12087
rect 16117 12047 16175 12053
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 19245 12087 19303 12093
rect 19245 12084 19257 12087
rect 19208 12056 19257 12084
rect 19208 12044 19214 12056
rect 19245 12053 19257 12056
rect 19291 12053 19303 12087
rect 20530 12084 20536 12096
rect 20491 12056 20536 12084
rect 19245 12047 19303 12053
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 23750 12084 23756 12096
rect 23711 12056 23756 12084
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 24302 12044 24308 12096
rect 24360 12084 24366 12096
rect 24489 12087 24547 12093
rect 24489 12084 24501 12087
rect 24360 12056 24501 12084
rect 24360 12044 24366 12056
rect 24489 12053 24501 12056
rect 24535 12053 24547 12087
rect 26510 12084 26516 12096
rect 26471 12056 26516 12084
rect 24489 12047 24547 12053
rect 26510 12044 26516 12056
rect 26568 12044 26574 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11880 1915 11883
rect 2222 11880 2228 11892
rect 1903 11852 2228 11880
rect 1903 11849 1915 11852
rect 1857 11843 1915 11849
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 2590 11880 2596 11892
rect 2363 11852 2596 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 3881 11883 3939 11889
rect 3881 11880 3893 11883
rect 3660 11852 3893 11880
rect 3660 11840 3666 11852
rect 3881 11849 3893 11852
rect 3927 11849 3939 11883
rect 3881 11843 3939 11849
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 4856 11852 5457 11880
rect 4856 11840 4862 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7800 11852 8217 11880
rect 7800 11840 7806 11852
rect 8205 11849 8217 11852
rect 8251 11880 8263 11883
rect 9950 11880 9956 11892
rect 8251 11852 9956 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 9950 11840 9956 11852
rect 10008 11880 10014 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 10008 11852 10057 11880
rect 10008 11840 10014 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 10870 11880 10876 11892
rect 10284 11852 10876 11880
rect 10284 11840 10290 11852
rect 10870 11840 10876 11852
rect 10928 11880 10934 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10928 11852 10977 11880
rect 10928 11840 10934 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 11330 11880 11336 11892
rect 11291 11852 11336 11880
rect 10965 11843 11023 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11701 11883 11759 11889
rect 11701 11880 11713 11883
rect 11572 11852 11713 11880
rect 11572 11840 11578 11852
rect 11701 11849 11713 11852
rect 11747 11849 11759 11883
rect 11701 11843 11759 11849
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 13964 11852 14657 11880
rect 13964 11840 13970 11852
rect 14645 11849 14657 11852
rect 14691 11880 14703 11883
rect 14691 11852 15240 11880
rect 14691 11849 14703 11852
rect 14645 11843 14703 11849
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 3418 11812 3424 11824
rect 2556 11784 3424 11812
rect 2556 11772 2562 11784
rect 3418 11772 3424 11784
rect 3476 11812 3482 11824
rect 10594 11812 10600 11824
rect 3476 11784 4108 11812
rect 10555 11784 10600 11812
rect 3476 11772 3482 11784
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 2130 11704 2136 11716
rect 2188 11744 2194 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2188 11716 2789 11744
rect 2188 11704 2194 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 2958 11744 2964 11756
rect 2919 11716 2964 11744
rect 2777 11707 2835 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 4080 11753 4108 11784
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 7650 11744 7656 11756
rect 7611 11716 7656 11744
rect 4065 11707 4123 11713
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 2731 11648 3341 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 3344 11540 3372 11639
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8536 11648 8677 11676
rect 8536 11636 8542 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 15212 11685 15240 11852
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15528 11852 15853 11880
rect 15528 11840 15534 11852
rect 15841 11849 15853 11852
rect 15887 11849 15899 11883
rect 15841 11843 15899 11849
rect 17865 11883 17923 11889
rect 17865 11849 17877 11883
rect 17911 11880 17923 11883
rect 18414 11880 18420 11892
rect 17911 11852 18420 11880
rect 17911 11849 17923 11852
rect 17865 11843 17923 11849
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 20806 11880 20812 11892
rect 20588 11852 20812 11880
rect 20588 11840 20594 11852
rect 20806 11840 20812 11852
rect 20864 11880 20870 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 20864 11852 21465 11880
rect 20864 11840 20870 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 23106 11880 23112 11892
rect 23067 11852 23112 11880
rect 21453 11843 21511 11849
rect 23106 11840 23112 11852
rect 23164 11840 23170 11892
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11880 23535 11883
rect 23566 11880 23572 11892
rect 23523 11852 23572 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 25041 11883 25099 11889
rect 25041 11849 25053 11883
rect 25087 11880 25099 11883
rect 25866 11880 25872 11892
rect 25087 11852 25872 11880
rect 25087 11849 25099 11852
rect 25041 11843 25099 11849
rect 25866 11840 25872 11852
rect 25924 11840 25930 11892
rect 27154 11840 27160 11892
rect 27212 11880 27218 11892
rect 28077 11883 28135 11889
rect 28077 11880 28089 11883
rect 27212 11852 28089 11880
rect 27212 11840 27218 11852
rect 28077 11849 28089 11852
rect 28123 11849 28135 11883
rect 28077 11843 28135 11849
rect 16298 11812 16304 11824
rect 16259 11784 16304 11812
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 18233 11815 18291 11821
rect 18233 11812 18245 11815
rect 18012 11784 18245 11812
rect 18012 11772 18018 11784
rect 18233 11781 18245 11784
rect 18279 11812 18291 11815
rect 18785 11815 18843 11821
rect 18785 11812 18797 11815
rect 18279 11784 18797 11812
rect 18279 11781 18291 11784
rect 18233 11775 18291 11781
rect 18785 11781 18797 11784
rect 18831 11812 18843 11815
rect 20898 11812 20904 11824
rect 18831 11784 19012 11812
rect 20859 11784 20904 11812
rect 18831 11781 18843 11784
rect 18785 11775 18843 11781
rect 15470 11744 15476 11756
rect 15383 11716 15476 11744
rect 15470 11704 15476 11716
rect 15528 11744 15534 11756
rect 16574 11744 16580 11756
rect 15528 11716 16580 11744
rect 15528 11704 15534 11716
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17494 11744 17500 11756
rect 17083 11716 17500 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 18984 11753 19012 11784
rect 20898 11772 20904 11784
rect 20956 11772 20962 11824
rect 21174 11812 21180 11824
rect 21135 11784 21180 11812
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 21818 11704 21824 11756
rect 21876 11744 21882 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21876 11716 22017 11744
rect 21876 11704 21882 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 23124 11744 23152 11840
rect 24302 11772 24308 11824
rect 24360 11812 24366 11824
rect 24360 11784 24532 11812
rect 24360 11772 24366 11784
rect 24504 11753 24532 11784
rect 25498 11772 25504 11824
rect 25556 11812 25562 11824
rect 25961 11815 26019 11821
rect 25961 11812 25973 11815
rect 25556 11784 25973 11812
rect 25556 11772 25562 11784
rect 25961 11781 25973 11784
rect 26007 11781 26019 11815
rect 25961 11775 26019 11781
rect 24397 11747 24455 11753
rect 24397 11744 24409 11747
rect 23124 11716 24409 11744
rect 22005 11707 22063 11713
rect 24397 11713 24409 11716
rect 24443 11713 24455 11747
rect 24397 11707 24455 11713
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 25682 11704 25688 11756
rect 25740 11744 25746 11756
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25740 11716 26157 11744
rect 25740 11704 25746 11716
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 8921 11679 8979 11685
rect 8921 11676 8933 11679
rect 8812 11648 8933 11676
rect 8812 11636 8818 11648
rect 8921 11645 8933 11648
rect 8967 11645 8979 11679
rect 8921 11639 8979 11645
rect 15197 11679 15255 11685
rect 15197 11645 15209 11679
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 15896 11648 16865 11676
rect 15896 11636 15902 11648
rect 16853 11645 16865 11648
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 20772 11648 21925 11676
rect 20772 11636 20778 11648
rect 21913 11645 21925 11648
rect 21959 11676 21971 11679
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 21959 11648 22477 11676
rect 21959 11645 21971 11648
rect 21913 11639 21971 11645
rect 22465 11645 22477 11648
rect 22511 11645 22523 11679
rect 22465 11639 22523 11645
rect 24118 11636 24124 11688
rect 24176 11676 24182 11688
rect 26418 11685 26424 11688
rect 24305 11679 24363 11685
rect 24305 11676 24317 11679
rect 24176 11648 24317 11676
rect 24176 11636 24182 11648
rect 24305 11645 24317 11648
rect 24351 11645 24363 11679
rect 26412 11676 26424 11685
rect 26379 11648 26424 11676
rect 24305 11639 24363 11645
rect 26412 11639 26424 11648
rect 26418 11636 26424 11639
rect 26476 11636 26482 11688
rect 4332 11611 4390 11617
rect 4332 11577 4344 11611
rect 4378 11608 4390 11611
rect 4706 11608 4712 11620
rect 4378 11580 4712 11608
rect 4378 11577 4390 11580
rect 4332 11571 4390 11577
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 5810 11568 5816 11620
rect 5868 11608 5874 11620
rect 7561 11611 7619 11617
rect 5868 11580 6500 11608
rect 5868 11568 5874 11580
rect 6472 11552 6500 11580
rect 7561 11577 7573 11611
rect 7607 11608 7619 11611
rect 8386 11608 8392 11620
rect 7607 11580 8392 11608
rect 7607 11577 7619 11580
rect 7561 11571 7619 11577
rect 8386 11568 8392 11580
rect 8444 11608 8450 11620
rect 9030 11608 9036 11620
rect 8444 11580 9036 11608
rect 8444 11568 8450 11580
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 14369 11611 14427 11617
rect 14369 11577 14381 11611
rect 14415 11608 14427 11611
rect 14415 11580 15332 11608
rect 14415 11577 14427 11580
rect 14369 11571 14427 11577
rect 15304 11552 15332 11580
rect 16482 11568 16488 11620
rect 16540 11608 16546 11620
rect 16761 11611 16819 11617
rect 16761 11608 16773 11611
rect 16540 11580 16773 11608
rect 16540 11568 16546 11580
rect 16761 11577 16773 11580
rect 16807 11608 16819 11611
rect 18138 11608 18144 11620
rect 16807 11580 18144 11608
rect 16807 11577 16819 11580
rect 16761 11571 16819 11577
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 19150 11568 19156 11620
rect 19208 11617 19214 11620
rect 19208 11611 19272 11617
rect 19208 11577 19226 11611
rect 19260 11577 19272 11611
rect 19208 11571 19272 11577
rect 19208 11568 19214 11571
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 21821 11611 21879 11617
rect 21821 11608 21833 11611
rect 20864 11580 21833 11608
rect 20864 11568 20870 11580
rect 21821 11577 21833 11580
rect 21867 11608 21879 11611
rect 22094 11608 22100 11620
rect 21867 11580 22100 11608
rect 21867 11577 21879 11580
rect 21821 11571 21879 11577
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 24578 11608 24584 11620
rect 22664 11580 24584 11608
rect 4522 11540 4528 11552
rect 3344 11512 4528 11540
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5684 11512 6009 11540
rect 5684 11500 5690 11512
rect 5997 11509 6009 11512
rect 6043 11509 6055 11543
rect 6454 11540 6460 11552
rect 6415 11512 6460 11540
rect 5997 11503 6055 11509
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 7098 11540 7104 11552
rect 7059 11512 7104 11540
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 7466 11540 7472 11552
rect 7427 11512 7472 11540
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 8478 11540 8484 11552
rect 8439 11512 8484 11540
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 14826 11540 14832 11552
rect 14787 11512 14832 11540
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 15286 11540 15292 11552
rect 15247 11512 15292 11540
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 16393 11543 16451 11549
rect 16393 11509 16405 11543
rect 16439 11540 16451 11543
rect 16574 11540 16580 11552
rect 16439 11512 16580 11540
rect 16439 11509 16451 11512
rect 16393 11503 16451 11509
rect 16574 11500 16580 11512
rect 16632 11500 16638 11552
rect 17494 11540 17500 11552
rect 17455 11512 17500 11540
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 20162 11500 20168 11552
rect 20220 11540 20226 11552
rect 20349 11543 20407 11549
rect 20349 11540 20361 11543
rect 20220 11512 20361 11540
rect 20220 11500 20226 11512
rect 20349 11509 20361 11512
rect 20395 11540 20407 11543
rect 21177 11543 21235 11549
rect 21177 11540 21189 11543
rect 20395 11512 21189 11540
rect 20395 11509 20407 11512
rect 20349 11503 20407 11509
rect 21177 11509 21189 11512
rect 21223 11540 21235 11543
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 21223 11512 21281 11540
rect 21223 11509 21235 11512
rect 21177 11503 21235 11509
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21269 11503 21327 11509
rect 21634 11500 21640 11552
rect 21692 11540 21698 11552
rect 22664 11540 22692 11580
rect 24578 11568 24584 11580
rect 24636 11608 24642 11620
rect 25593 11611 25651 11617
rect 25593 11608 25605 11611
rect 24636 11580 25605 11608
rect 24636 11568 24642 11580
rect 25593 11577 25605 11580
rect 25639 11608 25651 11611
rect 26878 11608 26884 11620
rect 25639 11580 26884 11608
rect 25639 11577 25651 11580
rect 25593 11571 25651 11577
rect 26878 11568 26884 11580
rect 26936 11568 26942 11620
rect 21692 11512 22692 11540
rect 21692 11500 21698 11512
rect 22738 11500 22744 11552
rect 22796 11540 22802 11552
rect 23937 11543 23995 11549
rect 23937 11540 23949 11543
rect 22796 11512 23949 11540
rect 22796 11500 22802 11512
rect 23937 11509 23949 11512
rect 23983 11509 23995 11543
rect 23937 11503 23995 11509
rect 26970 11500 26976 11552
rect 27028 11540 27034 11552
rect 27525 11543 27583 11549
rect 27525 11540 27537 11543
rect 27028 11512 27537 11540
rect 27028 11500 27034 11512
rect 27525 11509 27537 11512
rect 27571 11509 27583 11543
rect 27525 11503 27583 11509
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 3697 11339 3755 11345
rect 3697 11336 3709 11339
rect 2372 11308 3709 11336
rect 2372 11296 2378 11308
rect 3697 11305 3709 11308
rect 3743 11305 3755 11339
rect 3697 11299 3755 11305
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 4120 11308 4261 11336
rect 4120 11296 4126 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5592 11308 5825 11336
rect 5592 11296 5598 11308
rect 5813 11305 5825 11308
rect 5859 11336 5871 11339
rect 6270 11336 6276 11348
rect 5859 11308 6276 11336
rect 5859 11305 5871 11308
rect 5813 11299 5871 11305
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6914 11336 6920 11348
rect 6875 11308 6920 11336
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 7524 11308 9321 11336
rect 7524 11296 7530 11308
rect 9309 11305 9321 11308
rect 9355 11305 9367 11339
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 9309 11299 9367 11305
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 10502 11336 10508 11348
rect 10463 11308 10508 11336
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10928 11308 10977 11336
rect 10928 11296 10934 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 11422 11336 11428 11348
rect 11383 11308 11428 11336
rect 10965 11299 11023 11305
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 15470 11336 15476 11348
rect 14967 11308 15476 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 16025 11339 16083 11345
rect 16025 11336 16037 11339
rect 15896 11308 16037 11336
rect 15896 11296 15902 11308
rect 16025 11305 16037 11308
rect 16071 11305 16083 11339
rect 16025 11299 16083 11305
rect 16390 11296 16396 11348
rect 16448 11336 16454 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 16448 11308 16497 11336
rect 16448 11296 16454 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17037 11339 17095 11345
rect 17037 11336 17049 11339
rect 17000 11308 17049 11336
rect 17000 11296 17006 11308
rect 17037 11305 17049 11308
rect 17083 11305 17095 11339
rect 17037 11299 17095 11305
rect 17589 11339 17647 11345
rect 17589 11305 17601 11339
rect 17635 11336 17647 11339
rect 17862 11336 17868 11348
rect 17635 11308 17868 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 1118 11228 1124 11280
rect 1176 11268 1182 11280
rect 2685 11271 2743 11277
rect 2685 11268 2697 11271
rect 1176 11240 2697 11268
rect 1176 11228 1182 11240
rect 2332 11212 2360 11240
rect 2685 11237 2697 11240
rect 2731 11237 2743 11271
rect 3418 11268 3424 11280
rect 3379 11240 3424 11268
rect 2685 11231 2743 11237
rect 3418 11228 3424 11240
rect 3476 11268 3482 11280
rect 3602 11268 3608 11280
rect 3476 11240 3608 11268
rect 3476 11228 3482 11240
rect 3602 11228 3608 11240
rect 3660 11268 3666 11280
rect 4617 11271 4675 11277
rect 4617 11268 4629 11271
rect 3660 11240 4629 11268
rect 3660 11228 3666 11240
rect 4617 11237 4629 11240
rect 4663 11268 4675 11271
rect 4798 11268 4804 11280
rect 4663 11240 4804 11268
rect 4663 11237 4675 11240
rect 4617 11231 4675 11237
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 7282 11277 7288 11280
rect 7276 11268 7288 11277
rect 7243 11240 7288 11268
rect 7276 11231 7288 11240
rect 7282 11228 7288 11231
rect 7340 11228 7346 11280
rect 11330 11268 11336 11280
rect 11243 11240 11336 11268
rect 11330 11228 11336 11240
rect 11388 11268 11394 11280
rect 12434 11268 12440 11280
rect 11388 11240 12440 11268
rect 11388 11228 11394 11240
rect 12434 11228 12440 11240
rect 12492 11228 12498 11280
rect 17052 11268 17080 11299
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 19242 11336 19248 11348
rect 19203 11308 19248 11336
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19610 11336 19616 11348
rect 19392 11308 19616 11336
rect 19392 11296 19398 11308
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 21358 11336 21364 11348
rect 21319 11308 21364 11336
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22738 11336 22744 11348
rect 22152 11308 22197 11336
rect 22699 11308 22744 11336
rect 22152 11296 22158 11308
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 23658 11336 23664 11348
rect 23619 11308 23664 11336
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24305 11339 24363 11345
rect 24305 11305 24317 11339
rect 24351 11336 24363 11339
rect 24394 11336 24400 11348
rect 24351 11308 24400 11336
rect 24351 11305 24363 11308
rect 24305 11299 24363 11305
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25317 11339 25375 11345
rect 25317 11305 25329 11339
rect 25363 11336 25375 11339
rect 25590 11336 25596 11348
rect 25363 11308 25596 11336
rect 25363 11305 25375 11308
rect 25317 11299 25375 11305
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 25682 11296 25688 11348
rect 25740 11336 25746 11348
rect 26145 11339 26203 11345
rect 26145 11336 26157 11339
rect 25740 11308 26157 11336
rect 25740 11296 25746 11308
rect 26145 11305 26157 11308
rect 26191 11305 26203 11339
rect 26145 11299 26203 11305
rect 26510 11296 26516 11348
rect 26568 11336 26574 11348
rect 26973 11339 27031 11345
rect 26973 11336 26985 11339
rect 26568 11308 26985 11336
rect 26568 11296 26574 11308
rect 26973 11305 26985 11308
rect 27019 11336 27031 11339
rect 27614 11336 27620 11348
rect 27019 11308 27620 11336
rect 27019 11305 27031 11308
rect 26973 11299 27031 11305
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 18969 11271 19027 11277
rect 18969 11268 18981 11271
rect 17052 11240 18981 11268
rect 18969 11237 18981 11240
rect 19015 11268 19027 11271
rect 19150 11268 19156 11280
rect 19015 11240 19156 11268
rect 19015 11237 19027 11240
rect 18969 11231 19027 11237
rect 19150 11228 19156 11240
rect 19208 11228 19214 11280
rect 19426 11228 19432 11280
rect 19484 11268 19490 11280
rect 19705 11271 19763 11277
rect 19705 11268 19717 11271
rect 19484 11240 19717 11268
rect 19484 11228 19490 11240
rect 19705 11237 19717 11240
rect 19751 11237 19763 11271
rect 19705 11231 19763 11237
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 24213 11271 24271 11277
rect 24213 11268 24225 11271
rect 23532 11240 24225 11268
rect 23532 11228 23538 11240
rect 24213 11237 24225 11240
rect 24259 11268 24271 11271
rect 25409 11271 25467 11277
rect 25409 11268 25421 11271
rect 24259 11240 25421 11268
rect 24259 11237 24271 11240
rect 24213 11231 24271 11237
rect 25409 11237 25421 11240
rect 25455 11237 25467 11271
rect 26878 11268 26884 11280
rect 26839 11240 26884 11268
rect 25409 11231 25467 11237
rect 26878 11228 26884 11240
rect 26936 11228 26942 11280
rect 2314 11160 2320 11212
rect 2372 11160 2378 11212
rect 2590 11200 2596 11212
rect 2551 11172 2596 11200
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3936 11172 4077 11200
rect 3936 11160 3942 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 5810 11200 5816 11212
rect 5767 11172 5816 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 8478 11200 8484 11212
rect 7024 11172 8484 11200
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1811 11104 2145 11132
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 2133 11101 2145 11104
rect 2179 11132 2191 11135
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 2179 11104 2881 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2869 11101 2881 11104
rect 2915 11132 2927 11135
rect 2958 11132 2964 11144
rect 2915 11104 2964 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5828 11104 5917 11132
rect 2222 11064 2228 11076
rect 2135 11036 2228 11064
rect 2222 11024 2228 11036
rect 2280 11064 2286 11076
rect 4985 11067 5043 11073
rect 4985 11064 4997 11067
rect 2280 11036 4997 11064
rect 2280 11024 2286 11036
rect 4985 11033 4997 11036
rect 5031 11033 5043 11067
rect 5350 11064 5356 11076
rect 5311 11036 5356 11064
rect 4985 11027 5043 11033
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5828 10996 5856 11104
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 7024 11141 7052 11172
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 15838 11160 15844 11212
rect 15896 11200 15902 11212
rect 16393 11203 16451 11209
rect 16393 11200 16405 11203
rect 15896 11172 16405 11200
rect 15896 11160 15902 11172
rect 16393 11169 16405 11172
rect 16439 11200 16451 11203
rect 17402 11200 17408 11212
rect 16439 11172 17408 11200
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 21174 11200 21180 11212
rect 21087 11172 21180 11200
rect 21174 11160 21180 11172
rect 21232 11200 21238 11212
rect 21542 11200 21548 11212
rect 21232 11172 21548 11200
rect 21232 11160 21238 11172
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 22649 11203 22707 11209
rect 22649 11169 22661 11203
rect 22695 11200 22707 11203
rect 23293 11203 23351 11209
rect 23293 11200 23305 11203
rect 22695 11172 23305 11200
rect 22695 11169 22707 11172
rect 22649 11163 22707 11169
rect 23293 11169 23305 11172
rect 23339 11200 23351 11203
rect 23339 11172 23888 11200
rect 23339 11169 23351 11172
rect 23293 11163 23351 11169
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6328 11104 7021 11132
rect 6328 11092 6334 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 7009 11095 7067 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11296 11104 11621 11132
rect 11296 11092 11302 11104
rect 11609 11101 11621 11104
rect 11655 11132 11667 11135
rect 12710 11132 12716 11144
rect 11655 11104 12716 11132
rect 11655 11101 11667 11104
rect 11609 11095 11667 11101
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 16666 11132 16672 11144
rect 16579 11104 16672 11132
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 18414 11132 18420 11144
rect 18279 11104 18420 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11132 19947 11135
rect 20162 11132 20168 11144
rect 19935 11104 20168 11132
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 20162 11092 20168 11104
rect 20220 11092 20226 11144
rect 22922 11132 22928 11144
rect 22883 11104 22928 11132
rect 22922 11092 22928 11104
rect 22980 11092 22986 11144
rect 6457 11067 6515 11073
rect 6457 11033 6469 11067
rect 6503 11064 6515 11067
rect 6638 11064 6644 11076
rect 6503 11036 6644 11064
rect 6503 11033 6515 11036
rect 6457 11027 6515 11033
rect 6638 11024 6644 11036
rect 6696 11064 6702 11076
rect 8389 11067 8447 11073
rect 6696 11036 6868 11064
rect 6696 11024 6702 11036
rect 5132 10968 5856 10996
rect 6840 10996 6868 11036
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 8754 11064 8760 11076
rect 8435 11036 8760 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 7190 10996 7196 11008
rect 6840 10968 7196 10996
rect 5132 10956 5138 10968
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 8846 10956 8852 11008
rect 8904 10996 8910 11008
rect 8941 10999 8999 11005
rect 8941 10996 8953 10999
rect 8904 10968 8953 10996
rect 8904 10956 8910 10968
rect 8941 10965 8953 10968
rect 8987 10965 8999 10999
rect 16684 10996 16712 11092
rect 22281 11067 22339 11073
rect 22281 11033 22293 11067
rect 22327 11064 22339 11067
rect 23290 11064 23296 11076
rect 22327 11036 23296 11064
rect 22327 11033 22339 11036
rect 22281 11027 22339 11033
rect 23290 11024 23296 11036
rect 23348 11024 23354 11076
rect 23860 11073 23888 11172
rect 24302 11092 24308 11144
rect 24360 11132 24366 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 24360 11104 24409 11132
rect 24360 11092 24366 11104
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 26970 11092 26976 11144
rect 27028 11132 27034 11144
rect 27065 11135 27123 11141
rect 27065 11132 27077 11135
rect 27028 11104 27077 11132
rect 27028 11092 27034 11104
rect 27065 11101 27077 11104
rect 27111 11101 27123 11135
rect 27065 11095 27123 11101
rect 23845 11067 23903 11073
rect 23845 11033 23857 11067
rect 23891 11033 23903 11067
rect 23845 11027 23903 11033
rect 26326 11024 26332 11076
rect 26384 11064 26390 11076
rect 26513 11067 26571 11073
rect 26513 11064 26525 11067
rect 26384 11036 26525 11064
rect 26384 11024 26390 11036
rect 26513 11033 26525 11036
rect 26559 11033 26571 11067
rect 26513 11027 26571 11033
rect 16850 10996 16856 11008
rect 16684 10968 16856 10996
rect 8941 10959 8999 10965
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 21818 10996 21824 11008
rect 21779 10968 21824 10996
rect 21818 10956 21824 10968
rect 21876 10956 21882 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 2866 10792 2872 10804
rect 2372 10764 2872 10792
rect 2372 10752 2378 10764
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 3602 10792 3608 10804
rect 3344 10764 3608 10792
rect 2222 10656 2228 10668
rect 2183 10628 2228 10656
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2774 10656 2780 10668
rect 2372 10628 2780 10656
rect 2372 10616 2378 10628
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3344 10665 3372 10764
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4706 10792 4712 10804
rect 4667 10764 4712 10792
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 7466 10792 7472 10804
rect 7147 10764 7472 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8662 10792 8668 10804
rect 8623 10764 8668 10792
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 11238 10792 11244 10804
rect 11199 10764 11244 10792
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11480 10764 11529 10792
rect 11480 10752 11486 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 15838 10792 15844 10804
rect 12308 10764 15844 10792
rect 12308 10752 12314 10764
rect 15838 10752 15844 10764
rect 15896 10792 15902 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15896 10764 16037 10792
rect 15896 10752 15902 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 16390 10792 16396 10804
rect 16351 10764 16396 10792
rect 16025 10755 16083 10761
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 16632 10764 17233 10792
rect 16632 10752 16638 10764
rect 17221 10761 17233 10764
rect 17267 10792 17279 10795
rect 17862 10792 17868 10804
rect 17267 10764 17868 10792
rect 17267 10761 17279 10764
rect 17221 10755 17279 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18104 10764 18245 10792
rect 18104 10752 18110 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 19061 10795 19119 10801
rect 19061 10761 19073 10795
rect 19107 10792 19119 10795
rect 19242 10792 19248 10804
rect 19107 10764 19248 10792
rect 19107 10761 19119 10764
rect 19061 10755 19119 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 20622 10792 20628 10804
rect 19567 10764 20628 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 21266 10792 21272 10804
rect 21227 10764 21272 10792
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 23109 10795 23167 10801
rect 23109 10761 23121 10795
rect 23155 10792 23167 10795
rect 23382 10792 23388 10804
rect 23155 10764 23388 10792
rect 23155 10761 23167 10764
rect 23109 10755 23167 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 24394 10792 24400 10804
rect 23523 10764 24400 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 26878 10752 26884 10804
rect 26936 10792 26942 10804
rect 27157 10795 27215 10801
rect 27157 10792 27169 10795
rect 26936 10764 27169 10792
rect 26936 10752 26942 10764
rect 27157 10761 27169 10764
rect 27203 10761 27215 10795
rect 27157 10755 27215 10761
rect 27614 10752 27620 10804
rect 27672 10792 27678 10804
rect 27893 10795 27951 10801
rect 27893 10792 27905 10795
rect 27672 10764 27905 10792
rect 27672 10752 27678 10764
rect 27893 10761 27905 10764
rect 27939 10761 27951 10795
rect 27893 10755 27951 10761
rect 17681 10727 17739 10733
rect 17681 10693 17693 10727
rect 17727 10724 17739 10727
rect 18414 10724 18420 10736
rect 17727 10696 18420 10724
rect 17727 10693 17739 10696
rect 17681 10687 17739 10693
rect 18414 10684 18420 10696
rect 18472 10684 18478 10736
rect 21174 10724 21180 10736
rect 21135 10696 21180 10724
rect 21174 10684 21180 10696
rect 21232 10684 21238 10736
rect 24854 10684 24860 10736
rect 24912 10724 24918 10736
rect 26145 10727 26203 10733
rect 26145 10724 26157 10727
rect 24912 10696 26157 10724
rect 24912 10684 24918 10696
rect 26145 10693 26157 10696
rect 26191 10693 26203 10727
rect 26145 10687 26203 10693
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 3200 10628 3341 10656
rect 3200 10616 3206 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7650 10656 7656 10668
rect 7340 10628 7656 10656
rect 7340 10616 7346 10628
rect 7650 10616 7656 10628
rect 7708 10656 7714 10668
rect 8113 10659 8171 10665
rect 8113 10656 8125 10659
rect 7708 10628 8125 10656
rect 7708 10616 7714 10628
rect 8113 10625 8125 10628
rect 8159 10656 8171 10659
rect 8846 10656 8852 10668
rect 8159 10628 8852 10656
rect 8159 10625 8171 10628
rect 8113 10619 8171 10625
rect 8846 10616 8852 10628
rect 8904 10656 8910 10668
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 8904 10628 9229 10656
rect 8904 10616 8910 10628
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10656 18751 10659
rect 20162 10656 20168 10668
rect 18739 10628 20168 10656
rect 18739 10625 18751 10628
rect 18693 10619 18751 10625
rect 20162 10616 20168 10628
rect 20220 10656 20226 10668
rect 20220 10628 20668 10656
rect 20220 10616 20226 10628
rect 6273 10591 6331 10597
rect 6273 10557 6285 10591
rect 6319 10588 6331 10591
rect 7466 10588 7472 10600
rect 6319 10560 7472 10588
rect 6319 10557 6331 10560
rect 6273 10551 6331 10557
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10588 8631 10591
rect 8938 10588 8944 10600
rect 8619 10560 8944 10588
rect 8619 10557 8631 10560
rect 8573 10551 8631 10557
rect 8938 10548 8944 10560
rect 8996 10588 9002 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8996 10560 9045 10588
rect 8996 10548 9002 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9033 10551 9091 10557
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 10778 10588 10784 10600
rect 10275 10560 10784 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 19978 10588 19984 10600
rect 19939 10560 19984 10588
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10520 1731 10523
rect 2130 10520 2136 10532
rect 1719 10492 2136 10520
rect 1719 10489 1731 10492
rect 1673 10483 1731 10489
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 3574 10523 3632 10529
rect 3574 10520 3586 10523
rect 3476 10492 3586 10520
rect 3476 10480 3482 10492
rect 3574 10489 3586 10492
rect 3620 10489 3632 10523
rect 5810 10520 5816 10532
rect 5723 10492 5816 10520
rect 3574 10483 3632 10489
rect 5810 10480 5816 10492
rect 5868 10520 5874 10532
rect 6914 10520 6920 10532
rect 5868 10492 6920 10520
rect 5868 10480 5874 10492
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 19429 10523 19487 10529
rect 19429 10489 19441 10523
rect 19475 10520 19487 10523
rect 19886 10520 19892 10532
rect 19475 10492 19892 10520
rect 19475 10489 19487 10492
rect 19429 10483 19487 10489
rect 19886 10480 19892 10492
rect 19944 10480 19950 10532
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 3237 10455 3295 10461
rect 3237 10452 3249 10455
rect 2924 10424 3249 10452
rect 2924 10412 2930 10424
rect 3237 10421 3249 10424
rect 3283 10452 3295 10455
rect 3878 10452 3884 10464
rect 3283 10424 3884 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 4948 10424 6653 10452
rect 4948 10412 4954 10424
rect 6641 10421 6653 10424
rect 6687 10452 6699 10455
rect 7558 10452 7564 10464
rect 6687 10424 7564 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9677 10455 9735 10461
rect 9677 10452 9689 10455
rect 9180 10424 9689 10452
rect 9180 10412 9186 10424
rect 9677 10421 9689 10424
rect 9723 10421 9735 10455
rect 10410 10452 10416 10464
rect 10371 10424 10416 10452
rect 9677 10415 9735 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 20640 10461 20668 10628
rect 21358 10616 21364 10668
rect 21416 10656 21422 10668
rect 21818 10656 21824 10668
rect 21416 10628 21824 10656
rect 21416 10616 21422 10628
rect 21818 10616 21824 10628
rect 21876 10616 21882 10668
rect 23658 10656 23664 10668
rect 23619 10628 23664 10656
rect 23658 10616 23664 10628
rect 23716 10616 23722 10668
rect 26697 10659 26755 10665
rect 26697 10656 26709 10659
rect 25608 10628 26709 10656
rect 21634 10520 21640 10532
rect 21595 10492 21640 10520
rect 21634 10480 21640 10492
rect 21692 10480 21698 10532
rect 22649 10523 22707 10529
rect 22649 10520 22661 10523
rect 21744 10492 22661 10520
rect 20625 10455 20683 10461
rect 20625 10421 20637 10455
rect 20671 10452 20683 10455
rect 20806 10452 20812 10464
rect 20671 10424 20812 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 21744 10461 21772 10492
rect 22649 10489 22661 10492
rect 22695 10489 22707 10523
rect 22649 10483 22707 10489
rect 23382 10480 23388 10532
rect 23440 10520 23446 10532
rect 23906 10523 23964 10529
rect 23906 10520 23918 10523
rect 23440 10492 23918 10520
rect 23440 10480 23446 10492
rect 23906 10489 23918 10492
rect 23952 10520 23964 10523
rect 24302 10520 24308 10532
rect 23952 10492 24308 10520
rect 23952 10489 23964 10492
rect 23906 10483 23964 10489
rect 24302 10480 24308 10492
rect 24360 10520 24366 10532
rect 25608 10529 25636 10628
rect 26697 10625 26709 10628
rect 26743 10656 26755 10659
rect 26970 10656 26976 10668
rect 26743 10628 26976 10656
rect 26743 10625 26755 10628
rect 26697 10619 26755 10625
rect 26970 10616 26976 10628
rect 27028 10656 27034 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27028 10628 27537 10656
rect 27028 10616 27034 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 25958 10588 25964 10600
rect 25919 10560 25964 10588
rect 25958 10548 25964 10560
rect 26016 10588 26022 10600
rect 26513 10591 26571 10597
rect 26513 10588 26525 10591
rect 26016 10560 26525 10588
rect 26016 10548 26022 10560
rect 26513 10557 26525 10560
rect 26559 10588 26571 10591
rect 27154 10588 27160 10600
rect 26559 10560 27160 10588
rect 26559 10557 26571 10560
rect 26513 10551 26571 10557
rect 27154 10548 27160 10560
rect 27212 10548 27218 10600
rect 25593 10523 25651 10529
rect 25593 10520 25605 10523
rect 24360 10492 25605 10520
rect 24360 10480 24366 10492
rect 25593 10489 25605 10492
rect 25639 10489 25651 10523
rect 25593 10483 25651 10489
rect 26605 10523 26663 10529
rect 26605 10489 26617 10523
rect 26651 10520 26663 10523
rect 26694 10520 26700 10532
rect 26651 10492 26700 10520
rect 26651 10489 26663 10492
rect 26605 10483 26663 10489
rect 26694 10480 26700 10492
rect 26752 10480 26758 10532
rect 21729 10455 21787 10461
rect 21729 10452 21741 10455
rect 21600 10424 21741 10452
rect 21600 10412 21606 10424
rect 21729 10421 21741 10424
rect 21775 10421 21787 10455
rect 21729 10415 21787 10421
rect 22373 10455 22431 10461
rect 22373 10421 22385 10455
rect 22419 10452 22431 10455
rect 22922 10452 22928 10464
rect 22419 10424 22928 10452
rect 22419 10421 22431 10424
rect 22373 10415 22431 10421
rect 22922 10412 22928 10424
rect 22980 10452 22986 10464
rect 23750 10452 23756 10464
rect 22980 10424 23756 10452
rect 22980 10412 22986 10424
rect 23750 10412 23756 10424
rect 23808 10452 23814 10464
rect 25041 10455 25099 10461
rect 25041 10452 25053 10455
rect 23808 10424 25053 10452
rect 23808 10412 23814 10424
rect 25041 10421 25053 10424
rect 25087 10421 25099 10455
rect 25041 10415 25099 10421
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 1670 10248 1676 10260
rect 1627 10220 1676 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 5868 10220 6745 10248
rect 5868 10208 5874 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 7650 10248 7656 10260
rect 7611 10220 7656 10248
rect 6733 10211 6791 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 9122 10248 9128 10260
rect 7883 10220 9128 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 11057 10251 11115 10257
rect 11057 10217 11069 10251
rect 11103 10248 11115 10251
rect 11330 10248 11336 10260
rect 11103 10220 11336 10248
rect 11103 10217 11115 10220
rect 11057 10211 11115 10217
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 17957 10251 18015 10257
rect 17957 10217 17969 10251
rect 18003 10248 18015 10251
rect 18046 10248 18052 10260
rect 18003 10220 18052 10248
rect 18003 10217 18015 10220
rect 17957 10211 18015 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18322 10208 18328 10260
rect 18380 10248 18386 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 18380 10220 18429 10248
rect 18380 10208 18386 10220
rect 18417 10217 18429 10220
rect 18463 10248 18475 10251
rect 19150 10248 19156 10260
rect 18463 10220 19156 10248
rect 18463 10217 18475 10220
rect 18417 10211 18475 10217
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 19337 10251 19395 10257
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 19426 10248 19432 10260
rect 19383 10220 19432 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 19794 10248 19800 10260
rect 19755 10220 19800 10248
rect 19794 10208 19800 10220
rect 19852 10208 19858 10260
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 20036 10220 20085 10248
rect 20036 10208 20042 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 21358 10248 21364 10260
rect 21319 10220 21364 10248
rect 20073 10211 20131 10217
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 22002 10248 22008 10260
rect 21963 10220 22008 10248
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22738 10248 22744 10260
rect 22699 10220 22744 10248
rect 22738 10208 22744 10220
rect 22796 10208 22802 10260
rect 23382 10248 23388 10260
rect 23343 10220 23388 10248
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 26237 10251 26295 10257
rect 26237 10217 26249 10251
rect 26283 10248 26295 10251
rect 26694 10248 26700 10260
rect 26283 10220 26700 10248
rect 26283 10217 26295 10220
rect 26237 10211 26295 10217
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 26970 10208 26976 10260
rect 27028 10248 27034 10260
rect 27065 10251 27123 10257
rect 27065 10248 27077 10251
rect 27028 10220 27077 10248
rect 27028 10208 27034 10220
rect 27065 10217 27077 10220
rect 27111 10217 27123 10251
rect 27065 10211 27123 10217
rect 2777 10183 2835 10189
rect 2777 10149 2789 10183
rect 2823 10180 2835 10183
rect 4614 10180 4620 10192
rect 2823 10152 4620 10180
rect 2823 10149 2835 10152
rect 2777 10143 2835 10149
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 7668 10180 7696 10208
rect 8849 10183 8907 10189
rect 8849 10180 8861 10183
rect 7668 10152 8861 10180
rect 8849 10149 8861 10152
rect 8895 10149 8907 10183
rect 8849 10143 8907 10149
rect 21450 10140 21456 10192
rect 21508 10180 21514 10192
rect 21726 10180 21732 10192
rect 21508 10152 21732 10180
rect 21508 10140 21514 10152
rect 21726 10140 21732 10152
rect 21784 10180 21790 10192
rect 22097 10183 22155 10189
rect 22097 10180 22109 10183
rect 21784 10152 22109 10180
rect 21784 10140 21790 10152
rect 22097 10149 22109 10152
rect 22143 10149 22155 10183
rect 23658 10180 23664 10192
rect 22097 10143 22155 10149
rect 23492 10152 23664 10180
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 2590 10112 2596 10124
rect 2363 10084 2596 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 3786 10112 3792 10124
rect 2915 10084 3792 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3786 10072 3792 10084
rect 3844 10072 3850 10124
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5609 10115 5667 10121
rect 5609 10112 5621 10115
rect 5132 10084 5621 10112
rect 5132 10072 5138 10084
rect 5609 10081 5621 10084
rect 5655 10081 5667 10115
rect 5609 10075 5667 10081
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 8205 10115 8263 10121
rect 8205 10112 8217 10115
rect 7892 10084 8217 10112
rect 7892 10072 7898 10084
rect 8205 10081 8217 10084
rect 8251 10081 8263 10115
rect 18322 10112 18328 10124
rect 18283 10084 18328 10112
rect 8205 10075 8263 10081
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 23492 10121 23520 10152
rect 23658 10140 23664 10152
rect 23716 10140 23722 10192
rect 23750 10121 23756 10124
rect 23477 10115 23535 10121
rect 23477 10112 23489 10115
rect 23440 10084 23489 10112
rect 23440 10072 23446 10084
rect 23477 10081 23489 10084
rect 23523 10081 23535 10115
rect 23744 10112 23756 10121
rect 23711 10084 23756 10112
rect 23477 10075 23535 10081
rect 23744 10075 23756 10084
rect 23750 10072 23756 10075
rect 23808 10072 23814 10124
rect 26513 10115 26571 10121
rect 26513 10081 26525 10115
rect 26559 10112 26571 10115
rect 26602 10112 26608 10124
rect 26559 10084 26608 10112
rect 26559 10081 26571 10084
rect 26513 10075 26571 10081
rect 26602 10072 26608 10084
rect 26660 10072 26666 10124
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 2976 9976 3004 10007
rect 4798 10004 4804 10056
rect 4856 10044 4862 10056
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 4856 10016 5365 10044
rect 4856 10004 4862 10016
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 3418 9976 3424 9988
rect 2832 9948 3424 9976
rect 2832 9936 2838 9948
rect 3418 9936 3424 9948
rect 3476 9936 3482 9988
rect 1949 9911 2007 9917
rect 1949 9877 1961 9911
rect 1995 9908 2007 9911
rect 2038 9908 2044 9920
rect 1995 9880 2044 9908
rect 1995 9877 2007 9880
rect 1949 9871 2007 9877
rect 2038 9868 2044 9880
rect 2096 9908 2102 9920
rect 2314 9908 2320 9920
rect 2096 9880 2320 9908
rect 2096 9868 2102 9880
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4249 9911 4307 9917
rect 4249 9908 4261 9911
rect 4120 9880 4261 9908
rect 4120 9868 4126 9880
rect 4249 9877 4261 9880
rect 4295 9877 4307 9911
rect 4249 9871 4307 9877
rect 5074 9868 5080 9920
rect 5132 9908 5138 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 5132 9880 5181 9908
rect 5132 9868 5138 9880
rect 5169 9877 5181 9880
rect 5215 9877 5227 9911
rect 5368 9908 5396 10007
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8168 10016 8309 10044
rect 8168 10004 8174 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8478 10044 8484 10056
rect 8439 10016 8484 10044
rect 8297 10007 8355 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 18506 10004 18512 10056
rect 18564 10044 18570 10056
rect 22278 10044 22284 10056
rect 18564 10016 18609 10044
rect 22239 10016 22284 10044
rect 18564 10004 18570 10016
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 8496 9976 8524 10004
rect 7248 9948 8524 9976
rect 20717 9979 20775 9985
rect 7248 9936 7254 9948
rect 20717 9945 20729 9979
rect 20763 9976 20775 9979
rect 21634 9976 21640 9988
rect 20763 9948 21640 9976
rect 20763 9945 20775 9948
rect 20717 9939 20775 9945
rect 21634 9936 21640 9948
rect 21692 9936 21698 9988
rect 6270 9908 6276 9920
rect 5368 9880 6276 9908
rect 5169 9871 5227 9877
rect 6270 9868 6276 9880
rect 6328 9908 6334 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 6328 9880 7297 9908
rect 6328 9868 6334 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 24857 9911 24915 9917
rect 24857 9877 24869 9911
rect 24903 9908 24915 9911
rect 24946 9908 24952 9920
rect 24903 9880 24952 9908
rect 24903 9877 24915 9880
rect 24857 9871 24915 9877
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 26697 9911 26755 9917
rect 26697 9877 26709 9911
rect 26743 9908 26755 9911
rect 26970 9908 26976 9920
rect 26743 9880 26976 9908
rect 26743 9877 26755 9880
rect 26697 9871 26755 9877
rect 26970 9868 26976 9880
rect 27028 9868 27034 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 3142 9704 3148 9716
rect 2792 9676 3148 9704
rect 2685 9639 2743 9645
rect 2685 9605 2697 9639
rect 2731 9636 2743 9639
rect 2792 9636 2820 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 3476 9676 4200 9704
rect 3476 9664 3482 9676
rect 4172 9645 4200 9676
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 9214 9704 9220 9716
rect 8812 9676 9220 9704
rect 8812 9664 8818 9676
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 18506 9704 18512 9716
rect 17880 9676 18512 9704
rect 2731 9608 2820 9636
rect 4157 9639 4215 9645
rect 2731 9605 2743 9608
rect 2685 9599 2743 9605
rect 4157 9605 4169 9639
rect 4203 9605 4215 9639
rect 4157 9599 4215 9605
rect 2700 9568 2728 9599
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 4801 9639 4859 9645
rect 4801 9636 4813 9639
rect 4304 9608 4813 9636
rect 4304 9596 4310 9608
rect 4801 9605 4813 9608
rect 4847 9636 4859 9639
rect 4982 9636 4988 9648
rect 4847 9608 4988 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 5442 9636 5448 9648
rect 5403 9608 5448 9636
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5592 9608 5825 9636
rect 5592 9596 5598 9608
rect 5813 9605 5825 9608
rect 5859 9605 5871 9639
rect 6822 9636 6828 9648
rect 6783 9608 6828 9636
rect 5813 9599 5871 9605
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 8386 9636 8392 9648
rect 6932 9608 7512 9636
rect 8347 9608 8392 9636
rect 2608 9540 2728 9568
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1443 9472 1961 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1949 9469 1961 9472
rect 1995 9500 2007 9503
rect 2130 9500 2136 9512
rect 1995 9472 2136 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2608 9432 2636 9540
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5552 9500 5580 9596
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6932 9568 6960 9608
rect 6687 9540 6960 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7484 9577 7512 9608
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 9401 9639 9459 9645
rect 9401 9636 9413 9639
rect 8536 9608 9413 9636
rect 8536 9596 8542 9608
rect 9401 9605 9413 9608
rect 9447 9605 9459 9639
rect 9401 9599 9459 9605
rect 17129 9639 17187 9645
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 17494 9636 17500 9648
rect 17175 9608 17500 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 17494 9596 17500 9608
rect 17552 9636 17558 9648
rect 17880 9636 17908 9676
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 19150 9704 19156 9716
rect 19111 9676 19156 9704
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 21542 9664 21548 9716
rect 21600 9704 21606 9716
rect 21637 9707 21695 9713
rect 21637 9704 21649 9707
rect 21600 9676 21649 9704
rect 21600 9664 21606 9676
rect 21637 9673 21649 9676
rect 21683 9673 21695 9707
rect 21637 9667 21695 9673
rect 26602 9664 26608 9716
rect 26660 9704 26666 9716
rect 26973 9707 27031 9713
rect 26973 9704 26985 9707
rect 26660 9676 26985 9704
rect 26660 9664 26666 9676
rect 26973 9673 26985 9676
rect 27019 9673 27031 9707
rect 26973 9667 27031 9673
rect 18138 9636 18144 9648
rect 17552 9608 17908 9636
rect 18099 9608 18144 9636
rect 17552 9596 17558 9608
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 19702 9636 19708 9648
rect 19663 9608 19708 9636
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 20346 9596 20352 9648
rect 20404 9596 20410 9648
rect 23109 9639 23167 9645
rect 23109 9605 23121 9639
rect 23155 9636 23167 9639
rect 23382 9636 23388 9648
rect 23155 9608 23388 9636
rect 23155 9605 23167 9608
rect 23109 9599 23167 9605
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 23842 9636 23848 9648
rect 23803 9608 23848 9636
rect 23842 9596 23848 9608
rect 23900 9596 23906 9648
rect 26329 9639 26387 9645
rect 26329 9605 26341 9639
rect 26375 9636 26387 9639
rect 26878 9636 26884 9648
rect 26375 9608 26884 9636
rect 26375 9605 26387 9608
rect 26329 9599 26387 9605
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 7064 9540 7297 9568
rect 7064 9528 7070 9540
rect 7285 9537 7297 9540
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7650 9568 7656 9580
rect 7515 9540 7656 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7650 9528 7656 9540
rect 7708 9568 7714 9580
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 7708 9540 8953 9568
rect 7708 9528 7714 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 17773 9571 17831 9577
rect 17773 9568 17785 9571
rect 17092 9540 17785 9568
rect 17092 9528 17098 9540
rect 17773 9537 17785 9540
rect 17819 9568 17831 9571
rect 18414 9568 18420 9580
rect 17819 9540 18420 9568
rect 17819 9537 17831 9540
rect 17773 9531 17831 9537
rect 18414 9528 18420 9540
rect 18472 9568 18478 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 18472 9540 18613 9568
rect 18472 9528 18478 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 19242 9568 19248 9580
rect 18831 9540 19248 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 5307 9472 5580 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 2792 9432 2820 9463
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6788 9472 7205 9500
rect 6788 9460 6794 9472
rect 7193 9469 7205 9472
rect 7239 9500 7251 9503
rect 8846 9500 8852 9512
rect 7239 9472 8852 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 17497 9503 17555 9509
rect 17497 9500 17509 9503
rect 16908 9472 17509 9500
rect 16908 9460 16914 9472
rect 17497 9469 17509 9472
rect 17543 9500 17555 9503
rect 18800 9500 18828 9531
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19852 9540 20269 9568
rect 19852 9528 19858 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 20070 9500 20076 9512
rect 17543 9472 18828 9500
rect 19983 9472 20076 9500
rect 17543 9469 17555 9472
rect 17497 9463 17555 9469
rect 20070 9460 20076 9472
rect 20128 9500 20134 9512
rect 20364 9500 20392 9596
rect 20806 9568 20812 9580
rect 20719 9540 20812 9568
rect 20806 9528 20812 9540
rect 20864 9568 20870 9580
rect 22278 9568 22284 9580
rect 20864 9540 22284 9568
rect 20864 9528 20870 9540
rect 22278 9528 22284 9540
rect 22336 9568 22342 9580
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 22336 9540 22661 9568
rect 22336 9528 22342 9540
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9568 23535 9571
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 23523 9540 24501 9568
rect 23523 9537 23535 9540
rect 23477 9531 23535 9537
rect 24489 9537 24501 9540
rect 24535 9568 24547 9571
rect 24946 9568 24952 9580
rect 24535 9540 24952 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 20128 9472 20392 9500
rect 21177 9503 21235 9509
rect 20128 9460 20134 9472
rect 21177 9469 21189 9503
rect 21223 9500 21235 9503
rect 21818 9500 21824 9512
rect 21223 9472 21824 9500
rect 21223 9469 21235 9472
rect 21177 9463 21235 9469
rect 21818 9460 21824 9472
rect 21876 9500 21882 9512
rect 26436 9509 26464 9608
rect 26878 9596 26884 9608
rect 26936 9596 26942 9648
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21876 9472 22109 9500
rect 21876 9460 21882 9472
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 26421 9503 26479 9509
rect 26421 9469 26433 9503
rect 26467 9469 26479 9503
rect 26421 9463 26479 9469
rect 27430 9460 27436 9512
rect 27488 9500 27494 9512
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27488 9472 27537 9500
rect 27488 9460 27494 9472
rect 27525 9469 27537 9472
rect 27571 9500 27583 9503
rect 28077 9503 28135 9509
rect 28077 9500 28089 9503
rect 27571 9472 28089 9500
rect 27571 9469 27583 9472
rect 27525 9463 27583 9469
rect 28077 9469 28089 9472
rect 28123 9469 28135 9503
rect 28077 9463 28135 9469
rect 2608 9404 2820 9432
rect 3044 9435 3102 9441
rect 3044 9401 3056 9435
rect 3090 9432 3102 9435
rect 3418 9432 3424 9444
rect 3090 9404 3424 9432
rect 3090 9401 3102 9404
rect 3044 9395 3102 9401
rect 3418 9392 3424 9404
rect 3476 9392 3482 9444
rect 8297 9435 8355 9441
rect 8297 9401 8309 9435
rect 8343 9432 8355 9435
rect 8754 9432 8760 9444
rect 8343 9404 8760 9432
rect 8343 9401 8355 9404
rect 8297 9395 8355 9401
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 21450 9432 21456 9444
rect 21411 9404 21456 9432
rect 21450 9392 21456 9404
rect 21508 9432 21514 9444
rect 22005 9435 22063 9441
rect 22005 9432 22017 9435
rect 21508 9404 22017 9432
rect 21508 9392 21514 9404
rect 22005 9401 22017 9404
rect 22051 9401 22063 9435
rect 22005 9395 22063 9401
rect 23474 9392 23480 9444
rect 23532 9432 23538 9444
rect 24210 9432 24216 9444
rect 23532 9404 24216 9432
rect 23532 9392 23538 9404
rect 24210 9392 24216 9404
rect 24268 9392 24274 9444
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 1670 9364 1676 9376
rect 1627 9336 1676 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 4982 9324 4988 9376
rect 5040 9364 5046 9376
rect 5077 9367 5135 9373
rect 5077 9364 5089 9367
rect 5040 9336 5089 9364
rect 5040 9324 5046 9336
rect 5077 9333 5089 9336
rect 5123 9333 5135 9367
rect 5077 9327 5135 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5592 9336 6193 9364
rect 5592 9324 5598 9336
rect 6181 9333 6193 9336
rect 6227 9364 6239 9367
rect 6270 9364 6276 9376
rect 6227 9336 6276 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7340 9336 7849 9364
rect 7340 9324 7346 9336
rect 7837 9333 7849 9336
rect 7883 9364 7895 9367
rect 8110 9364 8116 9376
rect 7883 9336 8116 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8628 9336 8861 9364
rect 8628 9324 8634 9336
rect 8849 9333 8861 9336
rect 8895 9333 8907 9367
rect 8849 9327 8907 9333
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18012 9336 18521 9364
rect 18012 9324 18018 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 19613 9367 19671 9373
rect 19613 9333 19625 9367
rect 19659 9364 19671 9367
rect 20162 9364 20168 9376
rect 19659 9336 20168 9364
rect 19659 9333 19671 9336
rect 19613 9327 19671 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 24305 9367 24363 9373
rect 24305 9333 24317 9367
rect 24351 9364 24363 9367
rect 24486 9364 24492 9376
rect 24351 9336 24492 9364
rect 24351 9333 24363 9336
rect 24305 9327 24363 9333
rect 24486 9324 24492 9336
rect 24544 9324 24550 9376
rect 26605 9367 26663 9373
rect 26605 9333 26617 9367
rect 26651 9364 26663 9367
rect 26786 9364 26792 9376
rect 26651 9336 26792 9364
rect 26651 9333 26663 9336
rect 26605 9327 26663 9333
rect 26786 9324 26792 9336
rect 26844 9324 26850 9376
rect 27709 9367 27767 9373
rect 27709 9333 27721 9367
rect 27755 9364 27767 9367
rect 27798 9364 27804 9376
rect 27755 9336 27804 9364
rect 27755 9333 27767 9336
rect 27709 9327 27767 9333
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2038 9160 2044 9172
rect 1995 9132 2044 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2774 9160 2780 9172
rect 2363 9132 2780 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2774 9120 2780 9132
rect 2832 9120 2838 9172
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 2924 9132 2969 9160
rect 2924 9120 2930 9132
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3844 9132 4077 9160
rect 3844 9120 3850 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 5408 9132 5457 9160
rect 5408 9120 5414 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 6972 9132 8125 9160
rect 6972 9120 6978 9132
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 8113 9123 8171 9129
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8904 9132 8953 9160
rect 8904 9120 8910 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 17865 9163 17923 9169
rect 17865 9129 17877 9163
rect 17911 9160 17923 9163
rect 18322 9160 18328 9172
rect 17911 9132 18328 9160
rect 17911 9129 17923 9132
rect 17865 9123 17923 9129
rect 18322 9120 18328 9132
rect 18380 9160 18386 9172
rect 18509 9163 18567 9169
rect 18509 9160 18521 9163
rect 18380 9132 18521 9160
rect 18380 9120 18386 9132
rect 18509 9129 18521 9132
rect 18555 9129 18567 9163
rect 18509 9123 18567 9129
rect 18874 9120 18880 9172
rect 18932 9160 18938 9172
rect 18969 9163 19027 9169
rect 18969 9160 18981 9163
rect 18932 9132 18981 9160
rect 18932 9120 18938 9132
rect 18969 9129 18981 9132
rect 19015 9129 19027 9163
rect 18969 9123 19027 9129
rect 19797 9163 19855 9169
rect 19797 9129 19809 9163
rect 19843 9160 19855 9163
rect 20070 9160 20076 9172
rect 19843 9132 20076 9160
rect 19843 9129 19855 9132
rect 19797 9123 19855 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 21726 9160 21732 9172
rect 21687 9132 21732 9160
rect 21726 9120 21732 9132
rect 21784 9120 21790 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 23937 9163 23995 9169
rect 22152 9132 22197 9160
rect 22152 9120 22158 9132
rect 23937 9129 23949 9163
rect 23983 9160 23995 9163
rect 24486 9160 24492 9172
rect 23983 9132 24492 9160
rect 23983 9129 23995 9132
rect 23937 9123 23995 9129
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 24854 9160 24860 9172
rect 24815 9132 24860 9160
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 24949 9163 25007 9169
rect 24949 9129 24961 9163
rect 24995 9160 25007 9163
rect 25038 9160 25044 9172
rect 24995 9132 25044 9160
rect 24995 9129 25007 9132
rect 24949 9123 25007 9129
rect 25038 9120 25044 9132
rect 25096 9160 25102 9172
rect 26142 9160 26148 9172
rect 25096 9132 26148 9160
rect 25096 9120 25102 9132
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 2590 9052 2596 9104
rect 2648 9092 2654 9104
rect 2884 9092 2912 9120
rect 2648 9064 2912 9092
rect 2648 9052 2654 9064
rect 17954 9052 17960 9104
rect 18012 9092 18018 9104
rect 18141 9095 18199 9101
rect 18141 9092 18153 9095
rect 18012 9064 18153 9092
rect 18012 9052 18018 9064
rect 18141 9061 18153 9064
rect 18187 9061 18199 9095
rect 24210 9092 24216 9104
rect 24171 9064 24216 9092
rect 18141 9055 18199 9061
rect 24210 9052 24216 9064
rect 24268 9052 24274 9104
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3881 9027 3939 9033
rect 2832 8996 2877 9024
rect 2832 8984 2838 8996
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 4430 9024 4436 9036
rect 3927 8996 4436 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 5896 9027 5954 9033
rect 5896 8993 5908 9027
rect 5942 9024 5954 9027
rect 6270 9024 6276 9036
rect 5942 8996 6276 9024
rect 5942 8993 5954 8996
rect 5896 8987 5954 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 18598 8984 18604 9036
rect 18656 9024 18662 9036
rect 18877 9027 18935 9033
rect 18877 9024 18889 9027
rect 18656 8996 18889 9024
rect 18656 8984 18662 8996
rect 18877 8993 18889 8996
rect 18923 8993 18935 9027
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 18877 8987 18935 8993
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2096 8928 3065 8956
rect 2096 8916 2102 8928
rect 3053 8925 3065 8928
rect 3099 8956 3111 8959
rect 3510 8956 3516 8968
rect 3099 8928 3516 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 4522 8956 4528 8968
rect 4483 8928 4528 8956
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 5592 8928 5641 8956
rect 5592 8916 5598 8928
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 19153 8959 19211 8965
rect 19153 8925 19165 8959
rect 19199 8956 19211 8959
rect 19242 8956 19248 8968
rect 19199 8928 19248 8956
rect 19199 8925 19211 8928
rect 19153 8919 19211 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 23569 8959 23627 8965
rect 23569 8925 23581 8959
rect 23615 8956 23627 8959
rect 23750 8956 23756 8968
rect 23615 8928 23756 8956
rect 23615 8925 23627 8928
rect 23569 8919 23627 8925
rect 23750 8916 23756 8928
rect 23808 8956 23814 8968
rect 25133 8959 25191 8965
rect 25133 8956 25145 8959
rect 23808 8928 25145 8956
rect 23808 8916 23814 8928
rect 25133 8925 25145 8928
rect 25179 8956 25191 8959
rect 25222 8956 25228 8968
rect 25179 8928 25228 8956
rect 25179 8925 25191 8928
rect 25133 8919 25191 8925
rect 25222 8916 25228 8928
rect 25280 8916 25286 8968
rect 3418 8888 3424 8900
rect 3331 8860 3424 8888
rect 3418 8848 3424 8860
rect 3476 8888 3482 8900
rect 4724 8888 4752 8916
rect 3476 8860 4752 8888
rect 3476 8848 3482 8860
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8820 2467 8823
rect 2866 8820 2872 8832
rect 2455 8792 2872 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 5074 8820 5080 8832
rect 5035 8792 5080 8820
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 6730 8780 6736 8832
rect 6788 8820 6794 8832
rect 7009 8823 7067 8829
rect 7009 8820 7021 8823
rect 6788 8792 7021 8820
rect 6788 8780 6794 8792
rect 7009 8789 7021 8792
rect 7055 8789 7067 8823
rect 7834 8820 7840 8832
rect 7795 8792 7840 8820
rect 7009 8783 7067 8789
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 26694 8820 26700 8832
rect 26655 8792 26700 8820
rect 26694 8780 26700 8792
rect 26752 8780 26758 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4522 8616 4528 8628
rect 4120 8588 4528 8616
rect 4120 8576 4126 8588
rect 4522 8576 4528 8588
rect 4580 8616 4586 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 4580 8588 6837 8616
rect 4580 8576 4586 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 18598 8616 18604 8628
rect 18559 8588 18604 8616
rect 6825 8579 6883 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 18874 8616 18880 8628
rect 18835 8588 18880 8616
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 19242 8616 19248 8628
rect 19203 8588 19248 8616
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 24121 8619 24179 8625
rect 24121 8585 24133 8619
rect 24167 8616 24179 8619
rect 25038 8616 25044 8628
rect 24167 8588 25044 8616
rect 24167 8585 24179 8588
rect 24121 8579 24179 8585
rect 25038 8576 25044 8588
rect 25096 8576 25102 8628
rect 25222 8616 25228 8628
rect 25183 8588 25228 8616
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 25498 8616 25504 8628
rect 25459 8588 25504 8616
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26568 8588 27353 8616
rect 26568 8576 26574 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27706 8616 27712 8628
rect 27667 8588 27712 8616
rect 27341 8579 27399 8585
rect 27706 8576 27712 8588
rect 27764 8576 27770 8628
rect 1854 8508 1860 8560
rect 1912 8548 1918 8560
rect 4614 8548 4620 8560
rect 1912 8520 2084 8548
rect 4575 8520 4620 8548
rect 1912 8508 1918 8520
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2056 8489 2084 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 24397 8551 24455 8557
rect 4816 8520 5304 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 3568 8452 3617 8480
rect 3568 8440 3574 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 4203 8452 4537 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4525 8449 4537 8452
rect 4571 8480 4583 8483
rect 4706 8480 4712 8492
rect 4571 8452 4712 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4706 8440 4712 8452
rect 4764 8480 4770 8492
rect 4816 8480 4844 8520
rect 5074 8480 5080 8492
rect 4764 8452 4844 8480
rect 5035 8452 5080 8480
rect 4764 8440 4770 8452
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5276 8489 5304 8520
rect 24397 8517 24409 8551
rect 24443 8548 24455 8551
rect 25130 8548 25136 8560
rect 24443 8520 25136 8548
rect 24443 8517 24455 8520
rect 24397 8511 24455 8517
rect 25130 8508 25136 8520
rect 25188 8508 25194 8560
rect 26602 8548 26608 8560
rect 26563 8520 26608 8548
rect 26602 8508 26608 8520
rect 26660 8508 26666 8560
rect 27065 8551 27123 8557
rect 27065 8517 27077 8551
rect 27111 8548 27123 8551
rect 27246 8548 27252 8560
rect 27111 8520 27252 8548
rect 27111 8517 27123 8520
rect 27065 8511 27123 8517
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5810 8480 5816 8492
rect 5307 8452 5816 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6788 8452 7389 8480
rect 6788 8440 6794 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 7377 8443 7435 8449
rect 24228 8452 24869 8480
rect 1762 8372 1768 8424
rect 1820 8412 1826 8424
rect 1857 8415 1915 8421
rect 1857 8412 1869 8415
rect 1820 8384 1869 8412
rect 1820 8372 1826 8384
rect 1857 8381 1869 8384
rect 1903 8381 1915 8415
rect 1964 8412 1992 8440
rect 2590 8412 2596 8424
rect 1964 8384 2596 8412
rect 1857 8375 1915 8381
rect 1872 8344 1900 8375
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 2774 8412 2780 8424
rect 2700 8384 2780 8412
rect 2700 8344 2728 8384
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 3234 8412 3240 8424
rect 3007 8384 3240 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3234 8372 3240 8384
rect 3292 8412 3298 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3292 8384 3433 8412
rect 3292 8372 3298 8384
rect 3421 8381 3433 8384
rect 3467 8412 3479 8415
rect 3786 8412 3792 8424
rect 3467 8384 3792 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 5350 8412 5356 8424
rect 5031 8384 5356 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 7190 8412 7196 8424
rect 7151 8384 7196 8412
rect 7190 8372 7196 8384
rect 7248 8412 7254 8424
rect 24228 8421 24256 8452
rect 24857 8449 24869 8452
rect 24903 8480 24915 8483
rect 25682 8480 25688 8492
rect 24903 8452 25688 8480
rect 24903 8449 24915 8452
rect 24857 8443 24915 8449
rect 25682 8440 25688 8452
rect 25740 8440 25746 8492
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 7248 8384 8217 8412
rect 7248 8372 7254 8384
rect 8205 8381 8217 8384
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 24213 8415 24271 8421
rect 24213 8381 24225 8415
rect 24259 8381 24271 8415
rect 25314 8412 25320 8424
rect 25275 8384 25320 8412
rect 24213 8375 24271 8381
rect 25314 8372 25320 8384
rect 25372 8412 25378 8424
rect 25869 8415 25927 8421
rect 25869 8412 25881 8415
rect 25372 8384 25881 8412
rect 25372 8372 25378 8384
rect 25869 8381 25881 8384
rect 25915 8381 25927 8415
rect 25869 8375 25927 8381
rect 26421 8415 26479 8421
rect 26421 8381 26433 8415
rect 26467 8412 26479 8415
rect 27080 8412 27108 8511
rect 27246 8508 27252 8520
rect 27304 8508 27310 8560
rect 27522 8412 27528 8424
rect 26467 8384 27108 8412
rect 27483 8384 27528 8412
rect 26467 8381 26479 8384
rect 26421 8375 26479 8381
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27580 8384 28089 8412
rect 27580 8372 27586 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 1872 8316 2728 8344
rect 3513 8347 3571 8353
rect 3513 8313 3525 8347
rect 3559 8344 3571 8347
rect 3694 8344 3700 8356
rect 3559 8316 3700 8344
rect 3559 8313 3571 8316
rect 3513 8307 3571 8313
rect 3694 8304 3700 8316
rect 3752 8304 3758 8356
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 5592 8316 5733 8344
rect 5592 8304 5598 8316
rect 5721 8313 5733 8316
rect 5767 8344 5779 8347
rect 5902 8344 5908 8356
rect 5767 8316 5908 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 6270 8344 6276 8356
rect 6135 8316 6276 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 6270 8304 6276 8316
rect 6328 8304 6334 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 6972 8316 7297 8344
rect 6972 8304 6978 8316
rect 7285 8313 7297 8316
rect 7331 8344 7343 8347
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 7331 8316 7849 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 7837 8313 7849 8316
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 1489 8279 1547 8285
rect 1489 8245 1501 8279
rect 1535 8276 1547 8279
rect 1762 8276 1768 8288
rect 1535 8248 1768 8276
rect 1535 8245 1547 8248
rect 1489 8239 1547 8245
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 3050 8276 3056 8288
rect 3011 8248 3056 8276
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 5868 8248 6561 8276
rect 5868 8236 5874 8248
rect 6549 8245 6561 8248
rect 6595 8276 6607 8279
rect 6730 8276 6736 8288
rect 6595 8248 6736 8276
rect 6595 8245 6607 8248
rect 6549 8239 6607 8245
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1673 8075 1731 8081
rect 1673 8072 1685 8075
rect 1452 8044 1685 8072
rect 1452 8032 1458 8044
rect 1673 8041 1685 8044
rect 1719 8041 1731 8075
rect 1673 8035 1731 8041
rect 1688 8004 1716 8035
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 2130 8072 2136 8084
rect 1820 8044 2136 8072
rect 1820 8032 1826 8044
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2958 8072 2964 8084
rect 2823 8044 2964 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3510 8072 3516 8084
rect 3471 8044 3516 8072
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4062 8072 4068 8084
rect 3927 8044 4068 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4246 8072 4252 8084
rect 4207 8044 4252 8072
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5261 8075 5319 8081
rect 5261 8072 5273 8075
rect 5132 8044 5273 8072
rect 5132 8032 5138 8044
rect 5261 8041 5273 8044
rect 5307 8041 5319 8075
rect 5261 8035 5319 8041
rect 5629 8075 5687 8081
rect 5629 8041 5641 8075
rect 5675 8072 5687 8075
rect 5718 8072 5724 8084
rect 5675 8044 5724 8072
rect 5675 8041 5687 8044
rect 5629 8035 5687 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 24762 8072 24768 8084
rect 24627 8044 24768 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 25501 8075 25559 8081
rect 25501 8041 25513 8075
rect 25547 8072 25559 8075
rect 25590 8072 25596 8084
rect 25547 8044 25596 8072
rect 25547 8041 25559 8044
rect 25501 8035 25559 8041
rect 25590 8032 25596 8044
rect 25648 8032 25654 8084
rect 26326 8032 26332 8084
rect 26384 8072 26390 8084
rect 26510 8072 26516 8084
rect 26384 8044 26516 8072
rect 26384 8032 26390 8044
rect 26510 8032 26516 8044
rect 26568 8032 26574 8084
rect 2314 8004 2320 8016
rect 1688 7976 2320 8004
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 3145 8007 3203 8013
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 3694 8004 3700 8016
rect 3191 7976 3700 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 2038 7936 2044 7948
rect 1999 7908 2044 7936
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7868 2286 7880
rect 2682 7868 2688 7880
rect 2280 7840 2688 7868
rect 2280 7828 2286 7840
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 1394 7692 1400 7744
rect 1452 7732 1458 7744
rect 1578 7732 1584 7744
rect 1452 7704 1584 7732
rect 1452 7692 1458 7704
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 3160 7732 3188 7967
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4154 7936 4160 7948
rect 4111 7908 4160 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4154 7896 4160 7908
rect 4212 7936 4218 7948
rect 4890 7936 4896 7948
rect 4212 7908 4896 7936
rect 4212 7896 4218 7908
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 5592 7908 5733 7936
rect 5592 7896 5598 7908
rect 5721 7905 5733 7908
rect 5767 7936 5779 7939
rect 6362 7936 6368 7948
rect 5767 7908 6368 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7936 7251 7939
rect 7834 7936 7840 7948
rect 7239 7908 7840 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 25314 7936 25320 7948
rect 25275 7908 25320 7936
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 26513 7939 26571 7945
rect 26513 7905 26525 7939
rect 26559 7936 26571 7939
rect 27062 7936 27068 7948
rect 26559 7908 27068 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 27062 7896 27068 7908
rect 27120 7896 27126 7948
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5810 7868 5816 7880
rect 5040 7840 5816 7868
rect 5040 7828 5046 7840
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7282 7868 7288 7880
rect 6972 7840 7288 7868
rect 6972 7828 6978 7840
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7466 7868 7472 7880
rect 7427 7840 7472 7868
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 4801 7803 4859 7809
rect 4801 7769 4813 7803
rect 4847 7800 4859 7803
rect 4847 7772 5396 7800
rect 4847 7769 4859 7772
rect 4801 7763 4859 7769
rect 5368 7744 5396 7772
rect 2740 7704 3188 7732
rect 2740 7692 2746 7704
rect 4982 7692 4988 7744
rect 5040 7732 5046 7744
rect 5077 7735 5135 7741
rect 5077 7732 5089 7735
rect 5040 7704 5089 7732
rect 5040 7692 5046 7704
rect 5077 7701 5089 7704
rect 5123 7701 5135 7735
rect 5077 7695 5135 7701
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 6825 7735 6883 7741
rect 6825 7732 6837 7735
rect 5408 7704 6837 7732
rect 5408 7692 5414 7704
rect 6825 7701 6837 7704
rect 6871 7701 6883 7735
rect 6825 7695 6883 7701
rect 26326 7692 26332 7744
rect 26384 7732 26390 7744
rect 26697 7735 26755 7741
rect 26697 7732 26709 7735
rect 26384 7704 26709 7732
rect 26384 7692 26390 7704
rect 26697 7701 26709 7704
rect 26743 7701 26755 7735
rect 26697 7695 26755 7701
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2406 7528 2412 7540
rect 2096 7500 2412 7528
rect 2096 7488 2102 7500
rect 2406 7488 2412 7500
rect 2464 7528 2470 7540
rect 3053 7531 3111 7537
rect 3053 7528 3065 7531
rect 2464 7500 3065 7528
rect 2464 7488 2470 7500
rect 3053 7497 3065 7500
rect 3099 7497 3111 7531
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 3053 7491 3111 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4488 7500 4905 7528
rect 4488 7488 4494 7500
rect 4893 7497 4905 7500
rect 4939 7497 4951 7531
rect 4893 7491 4951 7497
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 5905 7531 5963 7537
rect 5905 7528 5917 7531
rect 5776 7500 5917 7528
rect 5776 7488 5782 7500
rect 5905 7497 5917 7500
rect 5951 7497 5963 7531
rect 6546 7528 6552 7540
rect 6507 7500 6552 7528
rect 5905 7491 5963 7497
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 25314 7528 25320 7540
rect 25275 7500 25320 7528
rect 25314 7488 25320 7500
rect 25372 7488 25378 7540
rect 27062 7488 27068 7540
rect 27120 7528 27126 7540
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 27120 7500 27353 7528
rect 27120 7488 27126 7500
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 1578 7460 1584 7472
rect 1539 7432 1584 7460
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 2222 7420 2228 7472
rect 2280 7460 2286 7472
rect 2317 7463 2375 7469
rect 2317 7460 2329 7463
rect 2280 7432 2329 7460
rect 2280 7420 2286 7432
rect 2317 7429 2329 7432
rect 2363 7429 2375 7463
rect 2317 7423 2375 7429
rect 4982 7420 4988 7472
rect 5040 7460 5046 7472
rect 5040 7432 5488 7460
rect 5040 7420 5046 7432
rect 2958 7392 2964 7404
rect 2871 7364 2964 7392
rect 2958 7352 2964 7364
rect 3016 7392 3022 7404
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 3016 7364 3617 7392
rect 3016 7352 3022 7364
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 5350 7392 5356 7404
rect 5311 7364 5356 7392
rect 3605 7355 3663 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5460 7401 5488 7432
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 6564 7392 6592 7488
rect 27706 7460 27712 7472
rect 27667 7432 27712 7460
rect 27706 7420 27712 7432
rect 27764 7420 27770 7472
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 6564 7364 7297 7392
rect 5445 7355 5503 7361
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7466 7392 7472 7404
rect 7427 7364 7472 7392
rect 7285 7355 7343 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7324 1458 7336
rect 1949 7327 2007 7333
rect 1949 7324 1961 7327
rect 1452 7296 1961 7324
rect 1452 7284 1458 7296
rect 1949 7293 1961 7296
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3418 7324 3424 7336
rect 3108 7296 3424 7324
rect 3108 7284 3114 7296
rect 3418 7284 3424 7296
rect 3476 7324 3482 7336
rect 3513 7327 3571 7333
rect 3513 7324 3525 7327
rect 3476 7296 3525 7324
rect 3476 7284 3482 7296
rect 3513 7293 3525 7296
rect 3559 7293 3571 7327
rect 3513 7287 3571 7293
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 5258 7324 5264 7336
rect 4847 7296 5264 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 26418 7324 26424 7336
rect 26379 7296 26424 7324
rect 26418 7284 26424 7296
rect 26476 7324 26482 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26476 7296 26985 7324
rect 26476 7284 26482 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 27522 7324 27528 7336
rect 27483 7296 27528 7324
rect 26973 7287 27031 7293
rect 27522 7284 27528 7296
rect 27580 7324 27586 7336
rect 28077 7327 28135 7333
rect 28077 7324 28089 7327
rect 27580 7296 28089 7324
rect 27580 7284 27586 7296
rect 28077 7293 28089 7296
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 2866 7148 2872 7200
rect 2924 7188 2930 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 2924 7160 3433 7188
rect 2924 7148 2930 7160
rect 3421 7157 3433 7160
rect 3467 7188 3479 7191
rect 3786 7188 3792 7200
rect 3467 7160 3792 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 3786 7148 3792 7160
rect 3844 7148 3850 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7834 7188 7840 7200
rect 7795 7160 7840 7188
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 26605 7191 26663 7197
rect 26605 7157 26617 7191
rect 26651 7188 26663 7191
rect 26878 7188 26884 7200
rect 26651 7160 26884 7188
rect 26651 7157 26663 7160
rect 26605 7151 26663 7157
rect 26878 7148 26884 7160
rect 26936 7148 26942 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 3418 6984 3424 6996
rect 3379 6956 3424 6984
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 3786 6984 3792 6996
rect 3747 6956 3792 6984
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4982 6984 4988 6996
rect 4943 6956 4988 6984
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5442 6984 5448 6996
rect 5403 6956 5448 6984
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7190 6984 7196 6996
rect 7151 6956 7196 6984
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 2958 6916 2964 6928
rect 2424 6888 2964 6916
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 1949 6851 2007 6857
rect 1949 6848 1961 6851
rect 1912 6820 1961 6848
rect 1912 6808 1918 6820
rect 1949 6817 1961 6820
rect 1995 6848 2007 6851
rect 2424 6848 2452 6888
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 5534 6916 5540 6928
rect 5460 6888 5540 6916
rect 1995 6820 2452 6848
rect 2501 6851 2559 6857
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 2501 6817 2513 6851
rect 2547 6848 2559 6851
rect 3510 6848 3516 6860
rect 2547 6820 3516 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4338 6848 4344 6860
rect 4111 6820 4344 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 5350 6848 5356 6860
rect 5263 6820 5356 6848
rect 5350 6808 5356 6820
rect 5408 6848 5414 6860
rect 5460 6848 5488 6888
rect 5534 6876 5540 6888
rect 5592 6876 5598 6928
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 7524 6888 7665 6916
rect 7524 6876 7530 6888
rect 7653 6885 7665 6888
rect 7699 6916 7711 6919
rect 8294 6916 8300 6928
rect 7699 6888 8300 6916
rect 7699 6885 7711 6888
rect 7653 6879 7711 6885
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 5810 6848 5816 6860
rect 5408 6820 5488 6848
rect 5771 6820 5816 6848
rect 5408 6808 5414 6820
rect 5810 6808 5816 6820
rect 5868 6848 5874 6860
rect 6454 6848 6460 6860
rect 5868 6820 6460 6848
rect 5868 6808 5874 6820
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 26510 6848 26516 6860
rect 26471 6820 26516 6848
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2590 6780 2596 6792
rect 2455 6752 2596 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2832 6752 3065 6780
rect 2832 6740 2838 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5592 6752 5917 6780
rect 5592 6740 5598 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6270 6780 6276 6792
rect 6135 6752 6276 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 2498 6672 2504 6724
rect 2556 6712 2562 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2556 6684 2697 6712
rect 2556 6672 2562 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 4212 6616 4261 6644
rect 4212 6604 4218 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 4249 6607 4307 6613
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 26694 6644 26700 6656
rect 26655 6616 26700 6644
rect 26694 6604 26700 6616
rect 26752 6604 26758 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 2409 6443 2467 6449
rect 2409 6440 2421 6443
rect 1452 6412 2421 6440
rect 1452 6400 1458 6412
rect 2409 6409 2421 6412
rect 2455 6440 2467 6443
rect 2682 6440 2688 6452
rect 2455 6412 2688 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 3142 6440 3148 6452
rect 3103 6412 3148 6440
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 4249 6443 4307 6449
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 4338 6440 4344 6452
rect 4295 6412 4344 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 6270 6440 6276 6452
rect 6183 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6440 6334 6452
rect 7466 6440 7472 6452
rect 6328 6412 7472 6440
rect 6328 6400 6334 6412
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 26602 6440 26608 6452
rect 26563 6412 26608 6440
rect 26602 6400 26608 6412
rect 26660 6400 26666 6452
rect 1578 6372 1584 6384
rect 1539 6344 1584 6372
rect 1578 6332 1584 6344
rect 1636 6332 1642 6384
rect 2038 6372 2044 6384
rect 1999 6344 2044 6372
rect 2038 6332 2044 6344
rect 2096 6332 2102 6384
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2056 6236 2084 6332
rect 3160 6304 3188 6400
rect 26510 6332 26516 6384
rect 26568 6372 26574 6384
rect 26973 6375 27031 6381
rect 26973 6372 26985 6375
rect 26568 6344 26985 6372
rect 26568 6332 26574 6344
rect 26973 6341 26985 6344
rect 27019 6341 27031 6375
rect 26973 6335 27031 6341
rect 2516 6276 3188 6304
rect 26329 6307 26387 6313
rect 2516 6245 2544 6276
rect 26329 6273 26341 6307
rect 26375 6304 26387 6307
rect 27154 6304 27160 6316
rect 26375 6276 27160 6304
rect 26375 6273 26387 6276
rect 26329 6267 26387 6273
rect 1443 6208 2084 6236
rect 2501 6239 2559 6245
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 3510 6236 3516 6248
rect 3471 6208 3516 6236
rect 2501 6199 2559 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 26436 6245 26464 6276
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 26421 6239 26479 6245
rect 3660 6208 3705 6236
rect 3660 6196 3666 6208
rect 26421 6205 26433 6239
rect 26467 6236 26479 6239
rect 26467 6208 26501 6236
rect 26467 6205 26479 6208
rect 26421 6199 26479 6205
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2685 6103 2743 6109
rect 2685 6100 2697 6103
rect 2280 6072 2697 6100
rect 2280 6060 2286 6072
rect 2685 6069 2697 6072
rect 2731 6069 2743 6103
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 2685 6063 2743 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 5810 6100 5816 6112
rect 5771 6072 5816 6100
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2041 5899 2099 5905
rect 2041 5865 2053 5899
rect 2087 5896 2099 5899
rect 2130 5896 2136 5908
rect 2087 5868 2136 5896
rect 2087 5865 2099 5868
rect 2041 5859 2099 5865
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 3602 5896 3608 5908
rect 3563 5868 3608 5896
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 2314 5788 2320 5840
rect 2372 5828 2378 5840
rect 3053 5831 3111 5837
rect 3053 5828 3065 5831
rect 2372 5800 3065 5828
rect 2372 5788 2378 5800
rect 3053 5797 3065 5800
rect 3099 5797 3111 5831
rect 3053 5791 3111 5797
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 1762 5760 1768 5772
rect 1443 5732 1768 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2498 5760 2504 5772
rect 2459 5732 2504 5760
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 26510 5760 26516 5772
rect 26471 5732 26516 5760
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 26694 5624 26700 5636
rect 26655 5596 26700 5624
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 2498 5352 2504 5364
rect 2459 5324 2504 5352
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26568 5324 27353 5352
rect 26568 5312 26574 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 27341 5315 27399 5321
rect 2038 5216 2044 5228
rect 1412 5188 2044 5216
rect 1412 5157 1440 5188
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 26418 5148 26424 5160
rect 26379 5120 26424 5148
rect 1397 5111 1455 5117
rect 26418 5108 26424 5120
rect 26476 5148 26482 5160
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26476 5120 26985 5148
rect 26476 5108 26482 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1762 4808 1768 4820
rect 1719 4780 1768 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 7190 2505 7196 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7184 2496 7196 2505
rect 6779 2468 7196 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7184 2459 7196 2468
rect 7190 2456 7196 2459
rect 7248 2456 7254 2508
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6288 2400 6929 2428
rect 4982 2252 4988 2304
rect 5040 2292 5046 2304
rect 5718 2292 5724 2304
rect 5040 2264 5724 2292
rect 5040 2252 5046 2264
rect 5718 2252 5724 2264
rect 5776 2292 5782 2304
rect 6288 2301 6316 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 6273 2295 6331 2301
rect 6273 2292 6285 2295
rect 5776 2264 6285 2292
rect 5776 2252 5782 2264
rect 6273 2261 6285 2264
rect 6319 2261 6331 2295
rect 6273 2255 6331 2261
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3332 22516 3384 22568
rect 7932 22516 7984 22568
rect 2964 22108 3016 22160
rect 13636 22108 13688 22160
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 27160 21088 27212 21140
rect 29000 21020 29052 21072
rect 23848 20952 23900 21004
rect 4068 20748 4120 20800
rect 5724 20748 5776 20800
rect 15568 20791 15620 20800
rect 15568 20757 15577 20791
rect 15577 20757 15611 20791
rect 15611 20757 15620 20791
rect 15568 20748 15620 20757
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 21272 20748 21324 20800
rect 25504 20748 25556 20800
rect 25780 20748 25832 20800
rect 26608 20748 26660 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 940 20544 992 20596
rect 8208 20544 8260 20596
rect 10232 20544 10284 20596
rect 14004 20544 14056 20596
rect 15844 20544 15896 20596
rect 17776 20544 17828 20596
rect 19616 20544 19668 20596
rect 21548 20544 21600 20596
rect 25228 20544 25280 20596
rect 4988 20519 5040 20528
rect 4988 20485 4997 20519
rect 4997 20485 5031 20519
rect 5031 20485 5040 20519
rect 4988 20476 5040 20485
rect 15568 20408 15620 20460
rect 19248 20408 19300 20460
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 4160 20340 4212 20392
rect 2412 20204 2464 20256
rect 7840 20204 7892 20256
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 14924 20340 14976 20392
rect 18052 20383 18104 20392
rect 14556 20315 14608 20324
rect 14556 20281 14565 20315
rect 14565 20281 14599 20315
rect 14599 20281 14608 20315
rect 14556 20272 14608 20281
rect 16396 20272 16448 20324
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 20720 20383 20772 20392
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 25780 20272 25832 20324
rect 9956 20204 10008 20256
rect 14004 20247 14056 20256
rect 14004 20213 14013 20247
rect 14013 20213 14047 20247
rect 14047 20213 14056 20247
rect 14004 20204 14056 20213
rect 14924 20247 14976 20256
rect 14924 20213 14933 20247
rect 14933 20213 14967 20247
rect 14967 20213 14976 20247
rect 14924 20204 14976 20213
rect 15108 20247 15160 20256
rect 15108 20213 15117 20247
rect 15117 20213 15151 20247
rect 15151 20213 15160 20247
rect 15108 20204 15160 20213
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 19156 20247 19208 20256
rect 19156 20213 19165 20247
rect 19165 20213 19199 20247
rect 19199 20213 19208 20247
rect 19156 20204 19208 20213
rect 19524 20247 19576 20256
rect 19524 20213 19533 20247
rect 19533 20213 19567 20247
rect 19567 20213 19576 20247
rect 19524 20204 19576 20213
rect 19616 20247 19668 20256
rect 19616 20213 19625 20247
rect 19625 20213 19659 20247
rect 19659 20213 19668 20247
rect 19616 20204 19668 20213
rect 23848 20204 23900 20256
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 25228 20204 25280 20256
rect 25504 20247 25556 20256
rect 25504 20213 25513 20247
rect 25513 20213 25547 20247
rect 25547 20213 25556 20247
rect 25504 20204 25556 20213
rect 25872 20247 25924 20256
rect 25872 20213 25881 20247
rect 25881 20213 25915 20247
rect 25915 20213 25924 20247
rect 25872 20204 25924 20213
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 15108 20000 15160 20052
rect 15476 20000 15528 20052
rect 17500 20000 17552 20052
rect 25504 19932 25556 19984
rect 11612 19864 11664 19916
rect 15200 19864 15252 19916
rect 16488 19864 16540 19916
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 24400 19864 24452 19916
rect 25044 19864 25096 19916
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 9036 19660 9088 19712
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11428 19660 11480 19712
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 15844 19839 15896 19848
rect 12532 19796 12584 19805
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 18604 19796 18656 19848
rect 25044 19728 25096 19780
rect 11980 19703 12032 19712
rect 11980 19669 11989 19703
rect 11989 19669 12023 19703
rect 12023 19669 12032 19703
rect 11980 19660 12032 19669
rect 12808 19660 12860 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 18328 19660 18380 19712
rect 19616 19660 19668 19712
rect 24768 19703 24820 19712
rect 24768 19669 24777 19703
rect 24777 19669 24811 19703
rect 24811 19669 24820 19703
rect 25412 19796 25464 19848
rect 26148 19796 26200 19848
rect 26516 19839 26568 19848
rect 26516 19805 26525 19839
rect 26525 19805 26559 19839
rect 26559 19805 26568 19839
rect 26516 19796 26568 19805
rect 25872 19703 25924 19712
rect 24768 19660 24820 19669
rect 25872 19669 25881 19703
rect 25881 19669 25915 19703
rect 25915 19669 25924 19703
rect 25872 19660 25924 19669
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 14004 19456 14056 19508
rect 24124 19456 24176 19508
rect 8760 19388 8812 19440
rect 9588 19388 9640 19440
rect 9496 19320 9548 19372
rect 10876 19320 10928 19372
rect 11336 19363 11388 19372
rect 3056 19252 3108 19304
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 12532 19320 12584 19372
rect 12348 19252 12400 19304
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 16488 19320 16540 19372
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 18236 19320 18288 19372
rect 18972 19252 19024 19304
rect 21824 19295 21876 19304
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 24216 19252 24268 19304
rect 25412 19456 25464 19508
rect 25872 19456 25924 19508
rect 25504 19388 25556 19440
rect 25044 19363 25096 19372
rect 25044 19329 25053 19363
rect 25053 19329 25087 19363
rect 25087 19329 25096 19363
rect 25044 19320 25096 19329
rect 2136 19184 2188 19236
rect 9588 19184 9640 19236
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 1952 19116 2004 19168
rect 2964 19159 3016 19168
rect 2964 19125 2973 19159
rect 2973 19125 3007 19159
rect 3007 19125 3016 19159
rect 2964 19116 3016 19125
rect 3240 19159 3292 19168
rect 3240 19125 3249 19159
rect 3249 19125 3283 19159
rect 3283 19125 3292 19159
rect 3240 19116 3292 19125
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 10692 19116 10744 19168
rect 11612 19116 11664 19168
rect 15108 19184 15160 19236
rect 18144 19184 18196 19236
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 13544 19159 13596 19168
rect 12900 19116 12952 19125
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 15200 19116 15252 19168
rect 15844 19116 15896 19168
rect 18604 19184 18656 19236
rect 19708 19184 19760 19236
rect 20260 19184 20312 19236
rect 18972 19159 19024 19168
rect 18972 19125 18981 19159
rect 18981 19125 19015 19159
rect 19015 19125 19024 19159
rect 18972 19116 19024 19125
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 22008 19159 22060 19168
rect 22008 19125 22017 19159
rect 22017 19125 22051 19159
rect 22051 19125 22060 19159
rect 22008 19116 22060 19125
rect 23756 19116 23808 19168
rect 27344 19320 27396 19372
rect 26516 19252 26568 19304
rect 25320 19116 25372 19168
rect 25688 19116 25740 19168
rect 27344 19159 27396 19168
rect 27344 19125 27353 19159
rect 27353 19125 27387 19159
rect 27387 19125 27396 19159
rect 27344 19116 27396 19125
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 3240 18912 3292 18964
rect 8760 18955 8812 18964
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 10324 18955 10376 18964
rect 10324 18921 10333 18955
rect 10333 18921 10367 18955
rect 10367 18921 10376 18955
rect 10324 18912 10376 18921
rect 11336 18955 11388 18964
rect 11336 18921 11345 18955
rect 11345 18921 11379 18955
rect 11379 18921 11388 18955
rect 11336 18912 11388 18921
rect 12532 18912 12584 18964
rect 15476 18955 15528 18964
rect 15476 18921 15485 18955
rect 15485 18921 15519 18955
rect 15519 18921 15528 18955
rect 15476 18912 15528 18921
rect 19156 18912 19208 18964
rect 21456 18912 21508 18964
rect 22468 18955 22520 18964
rect 22468 18921 22477 18955
rect 22477 18921 22511 18955
rect 22511 18921 22520 18955
rect 22468 18912 22520 18921
rect 25320 18955 25372 18964
rect 25320 18921 25329 18955
rect 25329 18921 25363 18955
rect 25363 18921 25372 18955
rect 25320 18912 25372 18921
rect 25780 18912 25832 18964
rect 26976 18955 27028 18964
rect 26976 18921 26985 18955
rect 26985 18921 27019 18955
rect 27019 18921 27028 18955
rect 26976 18912 27028 18921
rect 16856 18844 16908 18896
rect 24216 18887 24268 18896
rect 24216 18853 24250 18887
rect 24250 18853 24268 18887
rect 24216 18844 24268 18853
rect 1676 18776 1728 18828
rect 2688 18776 2740 18828
rect 2780 18776 2832 18828
rect 3424 18776 3476 18828
rect 5264 18819 5316 18828
rect 5264 18785 5273 18819
rect 5273 18785 5307 18819
rect 5307 18785 5316 18819
rect 5264 18776 5316 18785
rect 6460 18776 6512 18828
rect 8576 18819 8628 18828
rect 8576 18785 8585 18819
rect 8585 18785 8619 18819
rect 8619 18785 8628 18819
rect 8576 18776 8628 18785
rect 9036 18776 9088 18828
rect 9680 18776 9732 18828
rect 10692 18819 10744 18828
rect 10692 18785 10701 18819
rect 10701 18785 10735 18819
rect 10735 18785 10744 18819
rect 10692 18776 10744 18785
rect 17132 18776 17184 18828
rect 19432 18776 19484 18828
rect 22008 18776 22060 18828
rect 24676 18776 24728 18828
rect 26700 18776 26752 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 5172 18708 5224 18760
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 10784 18708 10836 18717
rect 11888 18751 11940 18760
rect 10600 18640 10652 18692
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 16948 18751 17000 18760
rect 16948 18717 16957 18751
rect 16957 18717 16991 18751
rect 16991 18717 17000 18751
rect 16948 18708 17000 18717
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 3332 18615 3384 18624
rect 3332 18581 3341 18615
rect 3341 18581 3375 18615
rect 3375 18581 3384 18615
rect 3332 18572 3384 18581
rect 3516 18572 3568 18624
rect 4160 18572 4212 18624
rect 22468 18640 22520 18692
rect 12992 18572 13044 18624
rect 15200 18572 15252 18624
rect 16304 18615 16356 18624
rect 16304 18581 16313 18615
rect 16313 18581 16347 18615
rect 16347 18581 16356 18615
rect 16304 18572 16356 18581
rect 18604 18572 18656 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 21548 18572 21600 18624
rect 27344 18708 27396 18760
rect 28172 18708 28224 18760
rect 23480 18615 23532 18624
rect 23480 18581 23489 18615
rect 23489 18581 23523 18615
rect 23523 18581 23532 18615
rect 23480 18572 23532 18581
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 9496 18368 9548 18420
rect 10324 18368 10376 18420
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12348 18368 12400 18420
rect 12716 18368 12768 18420
rect 16488 18411 16540 18420
rect 16488 18377 16497 18411
rect 16497 18377 16531 18411
rect 16531 18377 16540 18411
rect 16488 18368 16540 18377
rect 16948 18368 17000 18420
rect 17776 18411 17828 18420
rect 17776 18377 17785 18411
rect 17785 18377 17819 18411
rect 17819 18377 17828 18411
rect 17776 18368 17828 18377
rect 18144 18368 18196 18420
rect 3516 18300 3568 18352
rect 4896 18300 4948 18352
rect 5356 18300 5408 18352
rect 1584 18232 1636 18284
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 1676 18164 1728 18216
rect 2964 18164 3016 18216
rect 3240 18164 3292 18216
rect 5080 18232 5132 18284
rect 19156 18275 19208 18284
rect 19156 18241 19165 18275
rect 19165 18241 19199 18275
rect 19199 18241 19208 18275
rect 19156 18232 19208 18241
rect 19432 18232 19484 18284
rect 20444 18368 20496 18420
rect 21456 18411 21508 18420
rect 21456 18377 21465 18411
rect 21465 18377 21499 18411
rect 21499 18377 21508 18411
rect 21456 18368 21508 18377
rect 23112 18411 23164 18420
rect 23112 18377 23121 18411
rect 23121 18377 23155 18411
rect 23155 18377 23164 18411
rect 23112 18368 23164 18377
rect 26424 18368 26476 18420
rect 26976 18368 27028 18420
rect 24952 18300 25004 18352
rect 25412 18300 25464 18352
rect 20260 18232 20312 18284
rect 21548 18232 21600 18284
rect 23480 18232 23532 18284
rect 24768 18232 24820 18284
rect 4896 18164 4948 18216
rect 5172 18164 5224 18216
rect 8484 18164 8536 18216
rect 12348 18164 12400 18216
rect 12532 18164 12584 18216
rect 15016 18207 15068 18216
rect 15016 18173 15025 18207
rect 15025 18173 15059 18207
rect 15059 18173 15068 18207
rect 15016 18164 15068 18173
rect 5356 18139 5408 18148
rect 1860 18028 1912 18080
rect 2872 18071 2924 18080
rect 2872 18037 2881 18071
rect 2881 18037 2915 18071
rect 2915 18037 2924 18071
rect 2872 18028 2924 18037
rect 3516 18071 3568 18080
rect 3516 18037 3525 18071
rect 3525 18037 3559 18071
rect 3559 18037 3568 18071
rect 3516 18028 3568 18037
rect 4252 18028 4304 18080
rect 4988 18071 5040 18080
rect 4988 18037 4997 18071
rect 4997 18037 5031 18071
rect 5031 18037 5040 18071
rect 4988 18028 5040 18037
rect 5356 18105 5365 18139
rect 5365 18105 5399 18139
rect 5399 18105 5408 18139
rect 5356 18096 5408 18105
rect 13912 18096 13964 18148
rect 14280 18096 14332 18148
rect 15844 18096 15896 18148
rect 20352 18164 20404 18216
rect 20904 18164 20956 18216
rect 22008 18164 22060 18216
rect 23112 18164 23164 18216
rect 20536 18096 20588 18148
rect 20812 18096 20864 18148
rect 22652 18096 22704 18148
rect 22744 18096 22796 18148
rect 6460 18071 6512 18080
rect 6460 18037 6469 18071
rect 6469 18037 6503 18071
rect 6503 18037 6512 18071
rect 6460 18028 6512 18037
rect 7656 18071 7708 18080
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 8116 18071 8168 18080
rect 8116 18037 8125 18071
rect 8125 18037 8159 18071
rect 8159 18037 8168 18071
rect 8116 18028 8168 18037
rect 8484 18071 8536 18080
rect 8484 18037 8493 18071
rect 8493 18037 8527 18071
rect 8527 18037 8536 18071
rect 8484 18028 8536 18037
rect 12808 18028 12860 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 16948 18028 17000 18080
rect 17132 18028 17184 18080
rect 17868 18028 17920 18080
rect 18972 18028 19024 18080
rect 20168 18028 20220 18080
rect 21916 18028 21968 18080
rect 22100 18028 22152 18080
rect 23940 18071 23992 18080
rect 23940 18037 23949 18071
rect 23949 18037 23983 18071
rect 23983 18037 23992 18071
rect 23940 18028 23992 18037
rect 24032 18028 24084 18080
rect 24676 18028 24728 18080
rect 25412 18096 25464 18148
rect 26700 18096 26752 18148
rect 28172 18071 28224 18080
rect 28172 18037 28181 18071
rect 28181 18037 28215 18071
rect 28215 18037 28224 18071
rect 28172 18028 28224 18037
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 4344 17824 4396 17876
rect 5264 17824 5316 17876
rect 9036 17867 9088 17876
rect 9036 17833 9045 17867
rect 9045 17833 9079 17867
rect 9079 17833 9088 17867
rect 9036 17824 9088 17833
rect 9680 17824 9732 17876
rect 10784 17824 10836 17876
rect 11980 17824 12032 17876
rect 12440 17824 12492 17876
rect 13636 17867 13688 17876
rect 13636 17833 13645 17867
rect 13645 17833 13679 17867
rect 13679 17833 13688 17867
rect 13636 17824 13688 17833
rect 15108 17824 15160 17876
rect 15568 17824 15620 17876
rect 17776 17867 17828 17876
rect 17776 17833 17785 17867
rect 17785 17833 17819 17867
rect 17819 17833 17828 17867
rect 17776 17824 17828 17833
rect 17960 17824 18012 17876
rect 18144 17824 18196 17876
rect 18236 17824 18288 17876
rect 20168 17824 20220 17876
rect 20352 17867 20404 17876
rect 20352 17833 20361 17867
rect 20361 17833 20395 17867
rect 20395 17833 20404 17867
rect 20352 17824 20404 17833
rect 22008 17867 22060 17876
rect 22008 17833 22017 17867
rect 22017 17833 22051 17867
rect 22051 17833 22060 17867
rect 22008 17824 22060 17833
rect 2044 17756 2096 17808
rect 2964 17756 3016 17808
rect 9404 17756 9456 17808
rect 10692 17799 10744 17808
rect 10692 17765 10701 17799
rect 10701 17765 10735 17799
rect 10735 17765 10744 17799
rect 10692 17756 10744 17765
rect 11336 17756 11388 17808
rect 5080 17688 5132 17740
rect 8392 17731 8444 17740
rect 8392 17697 8401 17731
rect 8401 17697 8435 17731
rect 8435 17697 8444 17731
rect 8392 17688 8444 17697
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 1492 17663 1544 17672
rect 1492 17629 1501 17663
rect 1501 17629 1535 17663
rect 1535 17629 1544 17663
rect 1492 17620 1544 17629
rect 3884 17620 3936 17672
rect 7748 17620 7800 17672
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 9864 17620 9916 17672
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 12164 17663 12216 17672
rect 10232 17620 10284 17629
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 13820 17756 13872 17808
rect 16580 17756 16632 17808
rect 18788 17756 18840 17808
rect 25688 17756 25740 17808
rect 14372 17688 14424 17740
rect 15016 17688 15068 17740
rect 18512 17688 18564 17740
rect 21364 17688 21416 17740
rect 22376 17731 22428 17740
rect 22376 17697 22410 17731
rect 22410 17697 22428 17731
rect 22376 17688 22428 17697
rect 25780 17688 25832 17740
rect 26424 17688 26476 17740
rect 27804 17688 27856 17740
rect 14280 17620 14332 17672
rect 16304 17620 16356 17672
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 18420 17620 18472 17672
rect 2688 17552 2740 17604
rect 10968 17552 11020 17604
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 25504 17663 25556 17672
rect 20444 17552 20496 17604
rect 6368 17527 6420 17536
rect 6368 17493 6377 17527
rect 6377 17493 6411 17527
rect 6411 17493 6420 17527
rect 6368 17484 6420 17493
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 8116 17484 8168 17536
rect 8576 17484 8628 17536
rect 10416 17484 10468 17536
rect 12808 17527 12860 17536
rect 12808 17493 12817 17527
rect 12817 17493 12851 17527
rect 12851 17493 12860 17527
rect 12808 17484 12860 17493
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 21548 17527 21600 17536
rect 21548 17493 21557 17527
rect 21557 17493 21591 17527
rect 21591 17493 21600 17527
rect 21548 17484 21600 17493
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 27436 17620 27488 17672
rect 24124 17552 24176 17604
rect 25596 17552 25648 17604
rect 22284 17484 22336 17536
rect 24032 17527 24084 17536
rect 24032 17493 24041 17527
rect 24041 17493 24075 17527
rect 24075 17493 24084 17527
rect 24032 17484 24084 17493
rect 25228 17484 25280 17536
rect 25412 17484 25464 17536
rect 26332 17527 26384 17536
rect 26332 17493 26341 17527
rect 26341 17493 26375 17527
rect 26375 17493 26384 17527
rect 26332 17484 26384 17493
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 2964 17323 3016 17332
rect 2964 17289 2973 17323
rect 2973 17289 3007 17323
rect 3007 17289 3016 17323
rect 2964 17280 3016 17289
rect 5080 17280 5132 17332
rect 5540 17280 5592 17332
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 8392 17280 8444 17332
rect 9772 17280 9824 17332
rect 13544 17280 13596 17332
rect 14372 17280 14424 17332
rect 10692 17212 10744 17264
rect 1492 17144 1544 17196
rect 10968 17187 11020 17196
rect 1860 17119 1912 17128
rect 1860 17085 1894 17119
rect 1894 17085 1912 17119
rect 1860 17076 1912 17085
rect 2320 17076 2372 17128
rect 3884 17076 3936 17128
rect 4344 17119 4396 17128
rect 4344 17085 4378 17119
rect 4378 17085 4396 17119
rect 4344 17076 4396 17085
rect 7932 17076 7984 17128
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 12808 17212 12860 17264
rect 15016 17280 15068 17332
rect 16580 17280 16632 17332
rect 20444 17323 20496 17332
rect 20444 17289 20453 17323
rect 20453 17289 20487 17323
rect 20487 17289 20496 17323
rect 20444 17280 20496 17289
rect 21364 17323 21416 17332
rect 21364 17289 21373 17323
rect 21373 17289 21407 17323
rect 21407 17289 21416 17323
rect 21364 17280 21416 17289
rect 21824 17323 21876 17332
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 13636 17144 13688 17196
rect 18512 17212 18564 17264
rect 22284 17212 22336 17264
rect 24676 17280 24728 17332
rect 25320 17280 25372 17332
rect 26516 17323 26568 17332
rect 26516 17289 26525 17323
rect 26525 17289 26559 17323
rect 26559 17289 26568 17323
rect 26516 17280 26568 17289
rect 10048 17076 10100 17128
rect 12072 17076 12124 17128
rect 15108 17119 15160 17128
rect 3516 16983 3568 16992
rect 3516 16949 3525 16983
rect 3525 16949 3559 16983
rect 3559 16949 3568 16983
rect 6644 17008 6696 17060
rect 7748 17008 7800 17060
rect 8576 17008 8628 17060
rect 10416 17008 10468 17060
rect 3516 16940 3568 16949
rect 6828 16940 6880 16992
rect 7656 16940 7708 16992
rect 9404 16983 9456 16992
rect 9404 16949 9413 16983
rect 9413 16949 9447 16983
rect 9447 16949 9456 16983
rect 9404 16940 9456 16949
rect 9864 16940 9916 16992
rect 11336 16940 11388 16992
rect 15108 17085 15142 17119
rect 15142 17085 15160 17119
rect 15108 17076 15160 17085
rect 15384 17076 15436 17128
rect 18788 17119 18840 17128
rect 18788 17085 18822 17119
rect 18822 17085 18840 17119
rect 12072 16940 12124 16992
rect 12532 16940 12584 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 14280 16983 14332 16992
rect 14280 16949 14289 16983
rect 14289 16949 14323 16983
rect 14323 16949 14332 16983
rect 14280 16940 14332 16949
rect 15844 16940 15896 16992
rect 16396 16940 16448 16992
rect 18788 17076 18840 17085
rect 21640 17008 21692 17060
rect 25412 17144 25464 17196
rect 27528 17144 27580 17196
rect 28172 17144 28224 17196
rect 26332 17076 26384 17128
rect 24124 17008 24176 17060
rect 27252 17008 27304 17060
rect 27436 17008 27488 17060
rect 18972 16940 19024 16992
rect 19064 16940 19116 16992
rect 20260 16940 20312 16992
rect 22192 16983 22244 16992
rect 22192 16949 22201 16983
rect 22201 16949 22235 16983
rect 22235 16949 22244 16983
rect 22192 16940 22244 16949
rect 25504 16940 25556 16992
rect 26424 16983 26476 16992
rect 26424 16949 26433 16983
rect 26433 16949 26467 16983
rect 26467 16949 26476 16983
rect 26424 16940 26476 16949
rect 27804 16940 27856 16992
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 2780 16736 2832 16788
rect 4436 16779 4488 16788
rect 4436 16745 4445 16779
rect 4445 16745 4479 16779
rect 4479 16745 4488 16779
rect 4436 16736 4488 16745
rect 5540 16779 5592 16788
rect 5540 16745 5549 16779
rect 5549 16745 5583 16779
rect 5583 16745 5592 16779
rect 5540 16736 5592 16745
rect 6736 16736 6788 16788
rect 6920 16736 6972 16788
rect 8300 16736 8352 16788
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 13820 16736 13872 16788
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 16304 16736 16356 16788
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 17316 16779 17368 16788
rect 17316 16745 17325 16779
rect 17325 16745 17359 16779
rect 17359 16745 17368 16779
rect 17960 16779 18012 16788
rect 17316 16736 17368 16745
rect 17960 16745 17969 16779
rect 17969 16745 18003 16779
rect 18003 16745 18012 16779
rect 17960 16736 18012 16745
rect 18512 16779 18564 16788
rect 18512 16745 18521 16779
rect 18521 16745 18555 16779
rect 18555 16745 18564 16779
rect 18512 16736 18564 16745
rect 19432 16736 19484 16788
rect 21824 16736 21876 16788
rect 22192 16736 22244 16788
rect 24124 16779 24176 16788
rect 24124 16745 24133 16779
rect 24133 16745 24167 16779
rect 24167 16745 24176 16779
rect 24124 16736 24176 16745
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25504 16736 25556 16788
rect 26240 16736 26292 16788
rect 26332 16736 26384 16788
rect 2596 16668 2648 16720
rect 7472 16711 7524 16720
rect 7472 16677 7481 16711
rect 7481 16677 7515 16711
rect 7515 16677 7524 16711
rect 7472 16668 7524 16677
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 2780 16600 2832 16609
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 3700 16532 3752 16584
rect 4528 16575 4580 16584
rect 1492 16464 1544 16516
rect 2780 16464 2832 16516
rect 3516 16464 3568 16516
rect 4528 16541 4537 16575
rect 4537 16541 4571 16575
rect 4571 16541 4580 16575
rect 4528 16532 4580 16541
rect 5540 16600 5592 16652
rect 10324 16668 10376 16720
rect 10968 16668 11020 16720
rect 12440 16668 12492 16720
rect 13452 16643 13504 16652
rect 5632 16532 5684 16584
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 7656 16532 7708 16584
rect 7748 16532 7800 16584
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 22008 16668 22060 16720
rect 22100 16668 22152 16720
rect 25228 16711 25280 16720
rect 25228 16677 25237 16711
rect 25237 16677 25271 16711
rect 25271 16677 25280 16711
rect 25228 16668 25280 16677
rect 15660 16643 15712 16652
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 9864 16575 9916 16584
rect 8576 16532 8628 16541
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 10232 16532 10284 16584
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 13636 16532 13688 16584
rect 13820 16532 13872 16584
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16672 16600 16724 16652
rect 15752 16532 15804 16584
rect 11704 16464 11756 16516
rect 14280 16464 14332 16516
rect 18144 16600 18196 16652
rect 25780 16600 25832 16652
rect 26884 16643 26936 16652
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 19064 16575 19116 16584
rect 19064 16541 19073 16575
rect 19073 16541 19107 16575
rect 19107 16541 19116 16575
rect 19064 16532 19116 16541
rect 21548 16532 21600 16584
rect 25320 16575 25372 16584
rect 7932 16439 7984 16448
rect 7932 16405 7941 16439
rect 7941 16405 7975 16439
rect 7975 16405 7984 16439
rect 7932 16396 7984 16405
rect 8484 16396 8536 16448
rect 8668 16396 8720 16448
rect 15568 16396 15620 16448
rect 18512 16396 18564 16448
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 25320 16532 25372 16541
rect 25412 16575 25464 16584
rect 25412 16541 25421 16575
rect 25421 16541 25455 16575
rect 25455 16541 25464 16575
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 25412 16532 25464 16541
rect 25504 16464 25556 16516
rect 25872 16464 25924 16516
rect 21916 16396 21968 16448
rect 22284 16396 22336 16448
rect 22376 16396 22428 16448
rect 23756 16439 23808 16448
rect 23756 16405 23765 16439
rect 23765 16405 23799 16439
rect 23799 16405 23808 16439
rect 23756 16396 23808 16405
rect 26332 16396 26384 16448
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 3332 16192 3384 16244
rect 4436 16192 4488 16244
rect 5264 16192 5316 16244
rect 6460 16192 6512 16244
rect 8300 16192 8352 16244
rect 9864 16235 9916 16244
rect 9864 16201 9873 16235
rect 9873 16201 9907 16235
rect 9907 16201 9916 16235
rect 9864 16192 9916 16201
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 12164 16192 12216 16244
rect 16396 16192 16448 16244
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 18144 16192 18196 16244
rect 21180 16192 21232 16244
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 24860 16192 24912 16244
rect 27528 16235 27580 16244
rect 27528 16201 27537 16235
rect 27537 16201 27571 16235
rect 27571 16201 27580 16235
rect 27528 16192 27580 16201
rect 14648 16167 14700 16176
rect 2320 16056 2372 16108
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 3700 16099 3752 16108
rect 3700 16065 3709 16099
rect 3709 16065 3743 16099
rect 3743 16065 3752 16099
rect 3700 16056 3752 16065
rect 1768 15988 1820 16040
rect 2688 15988 2740 16040
rect 4712 15988 4764 16040
rect 10600 16056 10652 16108
rect 11980 16056 12032 16108
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 14648 16133 14657 16167
rect 14657 16133 14691 16167
rect 14691 16133 14700 16167
rect 14648 16124 14700 16133
rect 17316 16124 17368 16176
rect 21364 16124 21416 16176
rect 25504 16124 25556 16176
rect 15568 16056 15620 16108
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 6368 15988 6420 16040
rect 6828 15988 6880 16040
rect 7472 15988 7524 16040
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 12992 16031 13044 16040
rect 2872 15920 2924 15972
rect 5080 15963 5132 15972
rect 5080 15929 5089 15963
rect 5089 15929 5123 15963
rect 5123 15929 5132 15963
rect 5080 15920 5132 15929
rect 5816 15920 5868 15972
rect 8668 15920 8720 15972
rect 12992 15997 13026 16031
rect 13026 15997 13044 16031
rect 12992 15988 13044 15997
rect 14648 15988 14700 16040
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 15476 15920 15528 15972
rect 16396 15920 16448 15972
rect 17132 15920 17184 15972
rect 18512 15988 18564 16040
rect 22468 15988 22520 16040
rect 18972 15920 19024 15972
rect 23756 15988 23808 16040
rect 26148 16031 26200 16040
rect 26148 15997 26157 16031
rect 26157 15997 26191 16031
rect 26191 15997 26200 16031
rect 26148 15988 26200 15997
rect 24952 15920 25004 15972
rect 25872 15920 25924 15972
rect 26332 15920 26384 15972
rect 1584 15852 1636 15904
rect 3516 15895 3568 15904
rect 3516 15861 3525 15895
rect 3525 15861 3559 15895
rect 3559 15861 3568 15895
rect 3516 15852 3568 15861
rect 3792 15852 3844 15904
rect 4528 15852 4580 15904
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 7196 15895 7248 15904
rect 6552 15852 6604 15861
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 11520 15852 11572 15904
rect 12440 15852 12492 15904
rect 15016 15895 15068 15904
rect 15016 15861 15025 15895
rect 15025 15861 15059 15895
rect 15059 15861 15068 15895
rect 15016 15852 15068 15861
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 19340 15852 19392 15904
rect 21548 15852 21600 15904
rect 21732 15895 21784 15904
rect 21732 15861 21741 15895
rect 21741 15861 21775 15895
rect 21775 15861 21784 15895
rect 21732 15852 21784 15861
rect 21916 15852 21968 15904
rect 22100 15852 22152 15904
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 3700 15648 3752 15700
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 6920 15648 6972 15700
rect 5172 15580 5224 15632
rect 13820 15648 13872 15700
rect 15752 15648 15804 15700
rect 18420 15691 18472 15700
rect 18420 15657 18429 15691
rect 18429 15657 18463 15691
rect 18463 15657 18472 15691
rect 18420 15648 18472 15657
rect 21364 15648 21416 15700
rect 21548 15580 21600 15632
rect 22836 15580 22888 15632
rect 25320 15648 25372 15700
rect 24216 15580 24268 15632
rect 25412 15580 25464 15632
rect 26424 15580 26476 15632
rect 26976 15623 27028 15632
rect 26976 15589 26985 15623
rect 26985 15589 27019 15623
rect 27019 15589 27028 15623
rect 26976 15580 27028 15589
rect 2136 15555 2188 15564
rect 2136 15521 2145 15555
rect 2145 15521 2179 15555
rect 2179 15521 2188 15555
rect 2136 15512 2188 15521
rect 8392 15555 8444 15564
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 2504 15444 2556 15496
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2872 15308 2924 15360
rect 4712 15351 4764 15360
rect 4712 15317 4721 15351
rect 4721 15317 4755 15351
rect 4755 15317 4764 15351
rect 4712 15308 4764 15317
rect 8208 15444 8260 15496
rect 10324 15512 10376 15564
rect 11612 15512 11664 15564
rect 11704 15512 11756 15564
rect 13636 15512 13688 15564
rect 15568 15555 15620 15564
rect 15568 15521 15602 15555
rect 15602 15521 15620 15555
rect 15568 15512 15620 15521
rect 18788 15555 18840 15564
rect 18788 15521 18797 15555
rect 18797 15521 18831 15555
rect 18831 15521 18840 15555
rect 18788 15512 18840 15521
rect 22008 15512 22060 15564
rect 22560 15512 22612 15564
rect 24584 15512 24636 15564
rect 26240 15512 26292 15564
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 10876 15487 10928 15496
rect 8576 15444 8628 15453
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 4988 15308 5040 15360
rect 5724 15308 5776 15360
rect 6920 15308 6972 15360
rect 9588 15376 9640 15428
rect 7748 15308 7800 15360
rect 8116 15308 8168 15360
rect 8484 15308 8536 15360
rect 9680 15308 9732 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 11980 15308 12032 15360
rect 13452 15308 13504 15360
rect 13636 15308 13688 15360
rect 17960 15444 18012 15496
rect 19064 15444 19116 15496
rect 21732 15444 21784 15496
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 26332 15444 26384 15496
rect 27528 15444 27580 15496
rect 25412 15376 25464 15428
rect 16304 15308 16356 15360
rect 16580 15308 16632 15360
rect 17408 15308 17460 15360
rect 18420 15308 18472 15360
rect 21456 15308 21508 15360
rect 24124 15308 24176 15360
rect 26332 15308 26384 15360
rect 26976 15308 27028 15360
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 3700 15104 3752 15156
rect 3792 15104 3844 15156
rect 2780 15036 2832 15088
rect 3056 15036 3108 15088
rect 6828 15104 6880 15156
rect 8208 15104 8260 15156
rect 11612 15147 11664 15156
rect 11612 15113 11621 15147
rect 11621 15113 11655 15147
rect 11655 15113 11664 15147
rect 11612 15104 11664 15113
rect 11888 15104 11940 15156
rect 13176 15147 13228 15156
rect 13176 15113 13185 15147
rect 13185 15113 13219 15147
rect 13219 15113 13228 15147
rect 13176 15104 13228 15113
rect 18420 15147 18472 15156
rect 18420 15113 18429 15147
rect 18429 15113 18463 15147
rect 18463 15113 18472 15147
rect 18420 15104 18472 15113
rect 21640 15104 21692 15156
rect 25320 15104 25372 15156
rect 1492 14900 1544 14952
rect 9128 15036 9180 15088
rect 11980 15079 12032 15088
rect 11980 15045 11989 15079
rect 11989 15045 12023 15079
rect 12023 15045 12032 15079
rect 11980 15036 12032 15045
rect 7564 15011 7616 15020
rect 3792 14900 3844 14952
rect 4068 14900 4120 14952
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 8208 14968 8260 15020
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 21456 15036 21508 15088
rect 25044 15036 25096 15088
rect 26424 15104 26476 15156
rect 13912 14968 13964 15020
rect 14832 14968 14884 15020
rect 15384 14968 15436 15020
rect 15752 14968 15804 15020
rect 16488 14968 16540 15020
rect 19064 15011 19116 15020
rect 19064 14977 19073 15011
rect 19073 14977 19107 15011
rect 19107 14977 19116 15011
rect 19064 14968 19116 14977
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 23480 14968 23532 15020
rect 24124 15011 24176 15020
rect 4988 14900 5040 14952
rect 5632 14900 5684 14952
rect 5816 14900 5868 14952
rect 9680 14900 9732 14952
rect 2504 14832 2556 14884
rect 4712 14832 4764 14884
rect 5080 14832 5132 14884
rect 6552 14832 6604 14884
rect 9312 14832 9364 14884
rect 9864 14875 9916 14884
rect 9864 14841 9898 14875
rect 9898 14841 9916 14875
rect 9864 14832 9916 14841
rect 21732 14900 21784 14952
rect 1216 14764 1268 14816
rect 2228 14764 2280 14816
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 5172 14764 5224 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7656 14764 7708 14816
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 10324 14764 10376 14816
rect 10600 14764 10652 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 19340 14875 19392 14884
rect 19340 14841 19374 14875
rect 19374 14841 19392 14875
rect 19340 14832 19392 14841
rect 20352 14832 20404 14884
rect 22008 14900 22060 14952
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 14832 14807 14884 14816
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 15108 14764 15160 14816
rect 15384 14807 15436 14816
rect 15384 14773 15393 14807
rect 15393 14773 15427 14807
rect 15427 14773 15436 14807
rect 15384 14764 15436 14773
rect 16212 14764 16264 14816
rect 17868 14807 17920 14816
rect 17868 14773 17877 14807
rect 17877 14773 17911 14807
rect 17911 14773 17920 14807
rect 17868 14764 17920 14773
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 22560 14764 22612 14816
rect 23480 14807 23532 14816
rect 23480 14773 23489 14807
rect 23489 14773 23523 14807
rect 23523 14773 23532 14807
rect 23480 14764 23532 14773
rect 26148 14943 26200 14952
rect 26148 14909 26157 14943
rect 26157 14909 26191 14943
rect 26191 14909 26200 14943
rect 26148 14900 26200 14909
rect 25412 14832 25464 14884
rect 26332 14832 26384 14884
rect 24584 14764 24636 14816
rect 27528 14807 27580 14816
rect 27528 14773 27537 14807
rect 27537 14773 27571 14807
rect 27571 14773 27580 14807
rect 27528 14764 27580 14773
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 2504 14560 2556 14612
rect 3700 14560 3752 14612
rect 4988 14560 5040 14612
rect 6828 14560 6880 14612
rect 7196 14560 7248 14612
rect 10232 14560 10284 14612
rect 11704 14603 11756 14612
rect 11704 14569 11713 14603
rect 11713 14569 11747 14603
rect 11747 14569 11756 14603
rect 11704 14560 11756 14569
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 15384 14560 15436 14612
rect 18788 14560 18840 14612
rect 20352 14603 20404 14612
rect 20352 14569 20361 14603
rect 20361 14569 20395 14603
rect 20395 14569 20404 14603
rect 20352 14560 20404 14569
rect 24124 14560 24176 14612
rect 24860 14560 24912 14612
rect 26332 14560 26384 14612
rect 26608 14560 26660 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2780 14424 2832 14476
rect 4804 14424 4856 14476
rect 5724 14492 5776 14544
rect 9220 14492 9272 14544
rect 9588 14492 9640 14544
rect 9772 14492 9824 14544
rect 10140 14492 10192 14544
rect 16396 14535 16448 14544
rect 16396 14501 16430 14535
rect 16430 14501 16448 14535
rect 16396 14492 16448 14501
rect 19708 14535 19760 14544
rect 19708 14501 19717 14535
rect 19717 14501 19751 14535
rect 19751 14501 19760 14535
rect 19708 14492 19760 14501
rect 20536 14492 20588 14544
rect 23664 14492 23716 14544
rect 25136 14492 25188 14544
rect 25504 14535 25556 14544
rect 25504 14501 25513 14535
rect 25513 14501 25547 14535
rect 25547 14501 25556 14535
rect 25504 14492 25556 14501
rect 6184 14424 6236 14476
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 10692 14424 10744 14476
rect 10876 14424 10928 14476
rect 11244 14424 11296 14476
rect 13084 14424 13136 14476
rect 16212 14424 16264 14476
rect 19616 14467 19668 14476
rect 19616 14433 19625 14467
rect 19625 14433 19659 14467
rect 19659 14433 19668 14467
rect 19616 14424 19668 14433
rect 21088 14424 21140 14476
rect 26884 14467 26936 14476
rect 26884 14433 26893 14467
rect 26893 14433 26927 14467
rect 26927 14433 26936 14467
rect 26884 14424 26936 14433
rect 8852 14356 8904 14408
rect 9864 14356 9916 14408
rect 10600 14399 10652 14408
rect 10600 14365 10609 14399
rect 10609 14365 10643 14399
rect 10643 14365 10652 14399
rect 10600 14356 10652 14365
rect 19892 14399 19944 14408
rect 9036 14331 9088 14340
rect 9036 14297 9045 14331
rect 9045 14297 9079 14331
rect 9079 14297 9088 14331
rect 9036 14288 9088 14297
rect 9956 14288 10008 14340
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 4068 14220 4120 14272
rect 5632 14220 5684 14272
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 7932 14263 7984 14272
rect 7932 14229 7941 14263
rect 7941 14229 7975 14263
rect 7975 14229 7984 14263
rect 7932 14220 7984 14229
rect 9680 14220 9732 14272
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 21456 14356 21508 14408
rect 24032 14356 24084 14408
rect 26148 14399 26200 14408
rect 19340 14288 19392 14340
rect 11980 14220 12032 14272
rect 14832 14220 14884 14272
rect 15568 14220 15620 14272
rect 17500 14263 17552 14272
rect 17500 14229 17509 14263
rect 17509 14229 17543 14263
rect 17543 14229 17552 14263
rect 17500 14220 17552 14229
rect 18696 14263 18748 14272
rect 18696 14229 18705 14263
rect 18705 14229 18739 14263
rect 18739 14229 18748 14263
rect 18696 14220 18748 14229
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 19800 14220 19852 14272
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 22560 14220 22612 14272
rect 24308 14220 24360 14272
rect 26148 14365 26157 14399
rect 26157 14365 26191 14399
rect 26191 14365 26200 14399
rect 26148 14356 26200 14365
rect 26608 14356 26660 14408
rect 27160 14399 27212 14408
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 2136 14016 2188 14068
rect 3056 14059 3108 14068
rect 3056 14025 3065 14059
rect 3065 14025 3099 14059
rect 3099 14025 3108 14059
rect 3056 14016 3108 14025
rect 3976 14016 4028 14068
rect 4804 14016 4856 14068
rect 4988 14016 5040 14068
rect 7288 14016 7340 14068
rect 7932 14016 7984 14068
rect 8668 14016 8720 14068
rect 3240 13948 3292 14000
rect 5540 13948 5592 14000
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 2964 13880 3016 13932
rect 3884 13880 3936 13932
rect 4344 13880 4396 13932
rect 2596 13812 2648 13864
rect 4160 13812 4212 13864
rect 5080 13880 5132 13932
rect 6000 13880 6052 13932
rect 8116 13880 8168 13932
rect 6276 13855 6328 13864
rect 6276 13821 6285 13855
rect 6285 13821 6319 13855
rect 6319 13821 6328 13855
rect 6276 13812 6328 13821
rect 7196 13855 7248 13864
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 8484 13812 8536 13864
rect 10600 14016 10652 14068
rect 11244 14059 11296 14068
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 11980 14016 12032 14068
rect 14740 14016 14792 14068
rect 12440 13991 12492 14000
rect 12440 13957 12449 13991
rect 12449 13957 12483 13991
rect 12483 13957 12492 13991
rect 12440 13948 12492 13957
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 13268 13880 13320 13932
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 12716 13812 12768 13864
rect 15384 14016 15436 14068
rect 16396 14016 16448 14068
rect 16672 14016 16724 14068
rect 17684 14016 17736 14068
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 18236 14016 18288 14068
rect 18788 14016 18840 14068
rect 19616 14059 19668 14068
rect 19616 14025 19625 14059
rect 19625 14025 19659 14059
rect 19659 14025 19668 14059
rect 19616 14016 19668 14025
rect 21364 14016 21416 14068
rect 21456 14016 21508 14068
rect 21732 14059 21784 14068
rect 21732 14025 21741 14059
rect 21741 14025 21775 14059
rect 21775 14025 21784 14059
rect 21732 14016 21784 14025
rect 22836 14059 22888 14068
rect 22836 14025 22845 14059
rect 22845 14025 22879 14059
rect 22879 14025 22888 14059
rect 22836 14016 22888 14025
rect 23664 14016 23716 14068
rect 24032 14059 24084 14068
rect 24032 14025 24041 14059
rect 24041 14025 24075 14059
rect 24075 14025 24084 14059
rect 24032 14016 24084 14025
rect 25872 14016 25924 14068
rect 27160 14016 27212 14068
rect 18880 13948 18932 14000
rect 20812 13948 20864 14000
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 20352 13880 20404 13932
rect 26608 13948 26660 14000
rect 26792 13923 26844 13932
rect 26792 13889 26801 13923
rect 26801 13889 26835 13923
rect 26835 13889 26844 13923
rect 26792 13880 26844 13889
rect 27528 13923 27580 13932
rect 27528 13889 27537 13923
rect 27537 13889 27571 13923
rect 27571 13889 27580 13923
rect 27528 13880 27580 13889
rect 27712 13880 27764 13932
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 16304 13812 16356 13864
rect 11336 13787 11388 13796
rect 11336 13753 11345 13787
rect 11345 13753 11379 13787
rect 11379 13753 11388 13787
rect 11336 13744 11388 13753
rect 18788 13812 18840 13864
rect 19616 13812 19668 13864
rect 20260 13812 20312 13864
rect 22744 13812 22796 13864
rect 24308 13812 24360 13864
rect 17040 13744 17092 13796
rect 20444 13744 20496 13796
rect 21088 13744 21140 13796
rect 23940 13744 23992 13796
rect 27620 13744 27672 13796
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 2780 13676 2832 13728
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 5264 13676 5316 13728
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 12256 13719 12308 13728
rect 5632 13676 5684 13685
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 12992 13676 13044 13728
rect 14924 13676 14976 13728
rect 17684 13676 17736 13728
rect 18696 13676 18748 13728
rect 19248 13676 19300 13728
rect 20536 13719 20588 13728
rect 20536 13685 20545 13719
rect 20545 13685 20579 13719
rect 20579 13685 20588 13719
rect 20536 13676 20588 13685
rect 22100 13719 22152 13728
rect 22100 13685 22109 13719
rect 22109 13685 22143 13719
rect 22143 13685 22152 13719
rect 22100 13676 22152 13685
rect 25964 13676 26016 13728
rect 26792 13676 26844 13728
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 3976 13472 4028 13524
rect 1860 13404 1912 13456
rect 3700 13447 3752 13456
rect 3700 13413 3709 13447
rect 3709 13413 3743 13447
rect 3743 13413 3752 13447
rect 3700 13404 3752 13413
rect 5448 13472 5500 13524
rect 5724 13472 5776 13524
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 8852 13515 8904 13524
rect 8852 13481 8861 13515
rect 8861 13481 8895 13515
rect 8895 13481 8904 13515
rect 8852 13472 8904 13481
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 10232 13515 10284 13524
rect 10232 13481 10241 13515
rect 10241 13481 10275 13515
rect 10275 13481 10284 13515
rect 10232 13472 10284 13481
rect 12716 13515 12768 13524
rect 12716 13481 12725 13515
rect 12725 13481 12759 13515
rect 12759 13481 12768 13515
rect 12716 13472 12768 13481
rect 13084 13515 13136 13524
rect 13084 13481 13093 13515
rect 13093 13481 13127 13515
rect 13127 13481 13136 13515
rect 13084 13472 13136 13481
rect 13728 13472 13780 13524
rect 14924 13472 14976 13524
rect 15108 13472 15160 13524
rect 19892 13472 19944 13524
rect 20352 13515 20404 13524
rect 20352 13481 20361 13515
rect 20361 13481 20395 13515
rect 20395 13481 20404 13515
rect 20352 13472 20404 13481
rect 20536 13472 20588 13524
rect 21732 13472 21784 13524
rect 22100 13472 22152 13524
rect 23940 13472 23992 13524
rect 25412 13472 25464 13524
rect 25872 13472 25924 13524
rect 26884 13472 26936 13524
rect 26976 13515 27028 13524
rect 26976 13481 26985 13515
rect 26985 13481 27019 13515
rect 27019 13481 27028 13515
rect 26976 13472 27028 13481
rect 27712 13472 27764 13524
rect 5356 13404 5408 13456
rect 6460 13404 6512 13456
rect 6736 13404 6788 13456
rect 11704 13404 11756 13456
rect 13636 13404 13688 13456
rect 15476 13404 15528 13456
rect 17500 13404 17552 13456
rect 19708 13447 19760 13456
rect 19708 13413 19717 13447
rect 19717 13413 19751 13447
rect 19751 13413 19760 13447
rect 19708 13404 19760 13413
rect 1492 13336 1544 13388
rect 2504 13336 2556 13388
rect 15016 13336 15068 13388
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 4528 13268 4580 13320
rect 4896 13268 4948 13320
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 5724 13268 5776 13320
rect 5908 13268 5960 13320
rect 6276 13268 6328 13320
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 13176 13311 13228 13320
rect 6000 13200 6052 13252
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 20352 13268 20404 13320
rect 21456 13404 21508 13456
rect 23020 13404 23072 13456
rect 21916 13336 21968 13388
rect 24308 13404 24360 13456
rect 23756 13268 23808 13320
rect 26884 13379 26936 13388
rect 26884 13345 26893 13379
rect 26893 13345 26927 13379
rect 26927 13345 26936 13379
rect 26884 13336 26936 13345
rect 25964 13268 26016 13320
rect 27068 13311 27120 13320
rect 27068 13277 27077 13311
rect 27077 13277 27111 13311
rect 27111 13277 27120 13311
rect 27068 13268 27120 13277
rect 15292 13243 15344 13252
rect 15292 13209 15301 13243
rect 15301 13209 15335 13243
rect 15335 13209 15344 13243
rect 15292 13200 15344 13209
rect 2780 13175 2832 13184
rect 2780 13141 2789 13175
rect 2789 13141 2823 13175
rect 2823 13141 2832 13175
rect 2780 13132 2832 13141
rect 2964 13132 3016 13184
rect 4620 13132 4672 13184
rect 5264 13132 5316 13184
rect 7288 13132 7340 13184
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 11428 13132 11480 13184
rect 12808 13132 12860 13184
rect 12992 13132 13044 13184
rect 16948 13132 17000 13184
rect 17316 13132 17368 13184
rect 18420 13175 18472 13184
rect 18420 13141 18429 13175
rect 18429 13141 18463 13175
rect 18463 13141 18472 13175
rect 18420 13132 18472 13141
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 20996 13132 21048 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 2872 12928 2924 12980
rect 3700 12928 3752 12980
rect 5172 12928 5224 12980
rect 5448 12928 5500 12980
rect 6276 12928 6328 12980
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 11060 12928 11112 12980
rect 11520 12928 11572 12980
rect 13176 12928 13228 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 14556 12928 14608 12980
rect 15016 12971 15068 12980
rect 2504 12903 2556 12912
rect 2504 12869 2513 12903
rect 2513 12869 2547 12903
rect 2547 12869 2556 12903
rect 2504 12860 2556 12869
rect 8484 12860 8536 12912
rect 6460 12792 6512 12844
rect 7380 12792 7432 12844
rect 2964 12767 3016 12776
rect 2964 12733 2998 12767
rect 2998 12733 3016 12767
rect 2964 12724 3016 12733
rect 1216 12656 1268 12708
rect 1492 12588 1544 12640
rect 6552 12656 6604 12708
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 5448 12588 5500 12640
rect 7656 12724 7708 12776
rect 6828 12656 6880 12708
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 8668 12656 8720 12708
rect 11520 12792 11572 12844
rect 13360 12792 13412 12844
rect 9956 12724 10008 12776
rect 12624 12724 12676 12776
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 10876 12656 10928 12708
rect 15016 12937 15025 12971
rect 15025 12937 15059 12971
rect 15059 12937 15068 12971
rect 15016 12928 15068 12937
rect 15844 12928 15896 12980
rect 17132 12971 17184 12980
rect 17132 12937 17141 12971
rect 17141 12937 17175 12971
rect 17175 12937 17184 12971
rect 17132 12928 17184 12937
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 17960 12928 18012 12980
rect 20628 12928 20680 12980
rect 20812 12928 20864 12980
rect 22100 12928 22152 12980
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 23756 12860 23808 12912
rect 15200 12792 15252 12844
rect 15016 12724 15068 12776
rect 15752 12792 15804 12844
rect 17040 12792 17092 12844
rect 19156 12835 19208 12844
rect 16488 12724 16540 12776
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 20444 12792 20496 12844
rect 20996 12835 21048 12844
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 17776 12656 17828 12708
rect 19064 12699 19116 12708
rect 19064 12665 19073 12699
rect 19073 12665 19107 12699
rect 19107 12665 19116 12699
rect 19064 12656 19116 12665
rect 20812 12724 20864 12776
rect 22192 12724 22244 12776
rect 21640 12656 21692 12708
rect 23664 12656 23716 12708
rect 25320 12928 25372 12980
rect 26884 12928 26936 12980
rect 24032 12860 24084 12912
rect 26976 12860 27028 12912
rect 27068 12835 27120 12844
rect 27068 12801 27077 12835
rect 27077 12801 27111 12835
rect 27111 12801 27120 12835
rect 27068 12792 27120 12801
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 25412 12767 25464 12776
rect 25412 12733 25446 12767
rect 25446 12733 25464 12767
rect 25412 12724 25464 12733
rect 25688 12656 25740 12708
rect 8300 12588 8352 12640
rect 10784 12588 10836 12640
rect 11612 12588 11664 12640
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12440 12588 12492 12597
rect 16488 12631 16540 12640
rect 16488 12597 16497 12631
rect 16497 12597 16531 12631
rect 16531 12597 16540 12631
rect 16488 12588 16540 12597
rect 20720 12588 20772 12640
rect 21272 12588 21324 12640
rect 22192 12588 22244 12640
rect 22468 12631 22520 12640
rect 22468 12597 22477 12631
rect 22477 12597 22511 12631
rect 22511 12597 22520 12631
rect 22468 12588 22520 12597
rect 26424 12588 26476 12640
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 2504 12384 2556 12436
rect 2964 12384 3016 12436
rect 4804 12384 4856 12436
rect 2228 12316 2280 12368
rect 3240 12316 3292 12368
rect 5080 12316 5132 12368
rect 5448 12316 5500 12368
rect 6368 12384 6420 12436
rect 7840 12384 7892 12436
rect 10692 12384 10744 12436
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 13268 12384 13320 12436
rect 15016 12427 15068 12436
rect 15016 12393 15025 12427
rect 15025 12393 15059 12427
rect 15059 12393 15068 12427
rect 15016 12384 15068 12393
rect 15200 12384 15252 12436
rect 15568 12384 15620 12436
rect 16304 12384 16356 12436
rect 17776 12384 17828 12436
rect 21916 12384 21968 12436
rect 22560 12384 22612 12436
rect 24676 12427 24728 12436
rect 24676 12393 24685 12427
rect 24685 12393 24719 12427
rect 24719 12393 24728 12427
rect 24676 12384 24728 12393
rect 25412 12384 25464 12436
rect 7012 12316 7064 12368
rect 11520 12316 11572 12368
rect 15108 12316 15160 12368
rect 18420 12316 18472 12368
rect 21456 12316 21508 12368
rect 25596 12316 25648 12368
rect 26700 12316 26752 12368
rect 27436 12316 27488 12368
rect 2872 12248 2924 12300
rect 3608 12248 3660 12300
rect 5908 12291 5960 12300
rect 5908 12257 5917 12291
rect 5917 12257 5951 12291
rect 5951 12257 5960 12291
rect 5908 12248 5960 12257
rect 6368 12248 6420 12300
rect 6644 12248 6696 12300
rect 7104 12248 7156 12300
rect 10140 12291 10192 12300
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 5632 12180 5684 12232
rect 5816 12180 5868 12232
rect 6460 12180 6512 12232
rect 6920 12180 6972 12232
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 10508 12248 10560 12300
rect 10876 12248 10928 12300
rect 11336 12291 11388 12300
rect 11336 12257 11345 12291
rect 11345 12257 11379 12291
rect 11379 12257 11388 12291
rect 11336 12248 11388 12257
rect 15476 12248 15528 12300
rect 17040 12248 17092 12300
rect 17132 12248 17184 12300
rect 17960 12248 18012 12300
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 21180 12291 21232 12300
rect 21180 12257 21214 12291
rect 21214 12257 21232 12291
rect 21180 12248 21232 12257
rect 23572 12291 23624 12300
rect 23572 12257 23581 12291
rect 23581 12257 23615 12291
rect 23615 12257 23624 12291
rect 23572 12248 23624 12257
rect 24124 12291 24176 12300
rect 24124 12257 24133 12291
rect 24133 12257 24167 12291
rect 24167 12257 24176 12291
rect 24124 12248 24176 12257
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 16948 12223 17000 12232
rect 6736 12112 6788 12164
rect 9864 12112 9916 12164
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 24952 12180 25004 12232
rect 25136 12223 25188 12232
rect 25136 12189 25145 12223
rect 25145 12189 25179 12223
rect 25179 12189 25188 12223
rect 25136 12180 25188 12189
rect 25872 12248 25924 12300
rect 26884 12291 26936 12300
rect 26884 12257 26893 12291
rect 26893 12257 26927 12291
rect 26927 12257 26936 12291
rect 26884 12248 26936 12257
rect 25504 12180 25556 12232
rect 26608 12180 26660 12232
rect 27160 12223 27212 12232
rect 27160 12189 27169 12223
rect 27169 12189 27203 12223
rect 27203 12189 27212 12223
rect 27160 12180 27212 12189
rect 10600 12112 10652 12164
rect 15752 12112 15804 12164
rect 26424 12112 26476 12164
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 4712 12044 4764 12053
rect 6460 12044 6512 12096
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 7380 12044 7432 12096
rect 7656 12044 7708 12096
rect 8760 12044 8812 12096
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 10324 12044 10376 12096
rect 10692 12044 10744 12096
rect 10784 12044 10836 12096
rect 11704 12044 11756 12096
rect 13084 12044 13136 12096
rect 15844 12044 15896 12096
rect 19156 12044 19208 12096
rect 20536 12087 20588 12096
rect 20536 12053 20545 12087
rect 20545 12053 20579 12087
rect 20579 12053 20588 12087
rect 20536 12044 20588 12053
rect 23756 12087 23808 12096
rect 23756 12053 23765 12087
rect 23765 12053 23799 12087
rect 23799 12053 23808 12087
rect 23756 12044 23808 12053
rect 24308 12044 24360 12096
rect 26516 12087 26568 12096
rect 26516 12053 26525 12087
rect 26525 12053 26559 12087
rect 26559 12053 26568 12087
rect 26516 12044 26568 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2228 11840 2280 11892
rect 2596 11840 2648 11892
rect 3608 11840 3660 11892
rect 4804 11840 4856 11892
rect 7748 11840 7800 11892
rect 9956 11840 10008 11892
rect 10232 11840 10284 11892
rect 10876 11840 10928 11892
rect 11336 11883 11388 11892
rect 11336 11849 11345 11883
rect 11345 11849 11379 11883
rect 11379 11849 11388 11883
rect 11336 11840 11388 11849
rect 11520 11840 11572 11892
rect 13912 11840 13964 11892
rect 2504 11772 2556 11824
rect 3424 11772 3476 11824
rect 10600 11815 10652 11824
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 10600 11781 10609 11815
rect 10609 11781 10643 11815
rect 10643 11781 10652 11815
rect 10600 11772 10652 11781
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 8484 11636 8536 11688
rect 8760 11636 8812 11688
rect 15476 11840 15528 11892
rect 18420 11840 18472 11892
rect 20536 11840 20588 11892
rect 20812 11840 20864 11892
rect 23112 11883 23164 11892
rect 23112 11849 23121 11883
rect 23121 11849 23155 11883
rect 23155 11849 23164 11883
rect 23112 11840 23164 11849
rect 23572 11840 23624 11892
rect 25872 11840 25924 11892
rect 27160 11840 27212 11892
rect 16304 11815 16356 11824
rect 16304 11781 16313 11815
rect 16313 11781 16347 11815
rect 16347 11781 16356 11815
rect 16304 11772 16356 11781
rect 17960 11772 18012 11824
rect 20904 11815 20956 11824
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 16580 11704 16632 11756
rect 17500 11704 17552 11756
rect 20904 11781 20913 11815
rect 20913 11781 20947 11815
rect 20947 11781 20956 11815
rect 20904 11772 20956 11781
rect 21180 11815 21232 11824
rect 21180 11781 21189 11815
rect 21189 11781 21223 11815
rect 21223 11781 21232 11815
rect 21180 11772 21232 11781
rect 21824 11704 21876 11756
rect 24308 11772 24360 11824
rect 25504 11772 25556 11824
rect 25688 11704 25740 11756
rect 15844 11636 15896 11688
rect 20720 11636 20772 11688
rect 24124 11636 24176 11688
rect 26424 11679 26476 11688
rect 26424 11645 26458 11679
rect 26458 11645 26476 11679
rect 26424 11636 26476 11645
rect 4712 11568 4764 11620
rect 5816 11568 5868 11620
rect 8392 11568 8444 11620
rect 9036 11568 9088 11620
rect 16488 11568 16540 11620
rect 18144 11568 18196 11620
rect 19156 11568 19208 11620
rect 20812 11568 20864 11620
rect 22100 11568 22152 11620
rect 4528 11500 4580 11552
rect 5632 11500 5684 11552
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 7104 11543 7156 11552
rect 7104 11509 7113 11543
rect 7113 11509 7147 11543
rect 7147 11509 7156 11543
rect 7104 11500 7156 11509
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 7472 11500 7524 11509
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 8484 11500 8536 11509
rect 14832 11543 14884 11552
rect 14832 11509 14841 11543
rect 14841 11509 14875 11543
rect 14875 11509 14884 11543
rect 14832 11500 14884 11509
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 16580 11500 16632 11552
rect 17500 11543 17552 11552
rect 17500 11509 17509 11543
rect 17509 11509 17543 11543
rect 17543 11509 17552 11543
rect 17500 11500 17552 11509
rect 20168 11500 20220 11552
rect 21640 11500 21692 11552
rect 24584 11568 24636 11620
rect 26884 11568 26936 11620
rect 22744 11500 22796 11552
rect 26976 11500 27028 11552
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2320 11296 2372 11348
rect 4068 11296 4120 11348
rect 5540 11296 5592 11348
rect 6276 11296 6328 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 7472 11296 7524 11348
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 10508 11339 10560 11348
rect 10508 11305 10517 11339
rect 10517 11305 10551 11339
rect 10551 11305 10560 11339
rect 10508 11296 10560 11305
rect 10876 11296 10928 11348
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 15476 11296 15528 11348
rect 15844 11296 15896 11348
rect 16396 11296 16448 11348
rect 16948 11296 17000 11348
rect 1124 11228 1176 11280
rect 3424 11271 3476 11280
rect 3424 11237 3433 11271
rect 3433 11237 3467 11271
rect 3467 11237 3476 11271
rect 3424 11228 3476 11237
rect 3608 11228 3660 11280
rect 4804 11228 4856 11280
rect 7288 11271 7340 11280
rect 7288 11237 7322 11271
rect 7322 11237 7340 11271
rect 7288 11228 7340 11237
rect 11336 11271 11388 11280
rect 11336 11237 11345 11271
rect 11345 11237 11379 11271
rect 11379 11237 11388 11271
rect 11336 11228 11388 11237
rect 12440 11228 12492 11280
rect 17868 11296 17920 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19340 11296 19392 11348
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 22100 11339 22152 11348
rect 22100 11305 22109 11339
rect 22109 11305 22143 11339
rect 22143 11305 22152 11339
rect 22744 11339 22796 11348
rect 22100 11296 22152 11305
rect 22744 11305 22753 11339
rect 22753 11305 22787 11339
rect 22787 11305 22796 11339
rect 22744 11296 22796 11305
rect 23664 11339 23716 11348
rect 23664 11305 23673 11339
rect 23673 11305 23707 11339
rect 23707 11305 23716 11339
rect 23664 11296 23716 11305
rect 24400 11296 24452 11348
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 25596 11296 25648 11348
rect 25688 11296 25740 11348
rect 26516 11296 26568 11348
rect 27620 11296 27672 11348
rect 19156 11228 19208 11280
rect 19432 11228 19484 11280
rect 23480 11228 23532 11280
rect 26884 11271 26936 11280
rect 26884 11237 26893 11271
rect 26893 11237 26927 11271
rect 26927 11237 26936 11271
rect 26884 11228 26936 11237
rect 2320 11160 2372 11212
rect 2596 11203 2648 11212
rect 2596 11169 2605 11203
rect 2605 11169 2639 11203
rect 2639 11169 2648 11203
rect 2596 11160 2648 11169
rect 3884 11160 3936 11212
rect 5816 11160 5868 11212
rect 2964 11092 3016 11144
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 5356 11067 5408 11076
rect 5356 11033 5365 11067
rect 5365 11033 5399 11067
rect 5399 11033 5408 11067
rect 5356 11024 5408 11033
rect 5080 10956 5132 11008
rect 6276 11092 6328 11144
rect 8484 11160 8536 11212
rect 15844 11160 15896 11212
rect 17408 11160 17460 11212
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 21180 11203 21232 11212
rect 21180 11169 21189 11203
rect 21189 11169 21223 11203
rect 21223 11169 21232 11203
rect 21180 11160 21232 11169
rect 21548 11160 21600 11212
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11244 11092 11296 11144
rect 12716 11092 12768 11144
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18420 11092 18472 11144
rect 20168 11092 20220 11144
rect 22928 11135 22980 11144
rect 22928 11101 22937 11135
rect 22937 11101 22971 11135
rect 22971 11101 22980 11135
rect 22928 11092 22980 11101
rect 6644 11024 6696 11076
rect 8760 11024 8812 11076
rect 7196 10956 7248 11008
rect 8852 10956 8904 11008
rect 23296 11024 23348 11076
rect 24308 11092 24360 11144
rect 26976 11092 27028 11144
rect 26332 11024 26384 11076
rect 16856 10956 16908 11008
rect 21824 10999 21876 11008
rect 21824 10965 21833 10999
rect 21833 10965 21867 10999
rect 21867 10965 21876 10999
rect 21824 10956 21876 10965
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 2320 10752 2372 10804
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 2780 10616 2832 10668
rect 3148 10616 3200 10668
rect 3608 10752 3660 10804
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 7472 10752 7524 10804
rect 8668 10795 8720 10804
rect 8668 10761 8677 10795
rect 8677 10761 8711 10795
rect 8711 10761 8720 10795
rect 8668 10752 8720 10761
rect 11244 10795 11296 10804
rect 11244 10761 11253 10795
rect 11253 10761 11287 10795
rect 11287 10761 11296 10795
rect 11244 10752 11296 10761
rect 11428 10752 11480 10804
rect 12256 10752 12308 10804
rect 15844 10752 15896 10804
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 16580 10752 16632 10804
rect 17868 10752 17920 10804
rect 18052 10752 18104 10804
rect 19248 10752 19300 10804
rect 20628 10752 20680 10804
rect 21272 10795 21324 10804
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 23388 10752 23440 10804
rect 24400 10752 24452 10804
rect 26884 10752 26936 10804
rect 27620 10752 27672 10804
rect 18420 10684 18472 10736
rect 21180 10727 21232 10736
rect 21180 10693 21189 10727
rect 21189 10693 21223 10727
rect 21223 10693 21232 10727
rect 21180 10684 21232 10693
rect 24860 10684 24912 10736
rect 7288 10616 7340 10668
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 8852 10616 8904 10668
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 8944 10548 8996 10600
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 2136 10523 2188 10532
rect 2136 10489 2145 10523
rect 2145 10489 2179 10523
rect 2179 10489 2188 10523
rect 2136 10480 2188 10489
rect 3424 10480 3476 10532
rect 5816 10523 5868 10532
rect 5816 10489 5825 10523
rect 5825 10489 5859 10523
rect 5859 10489 5868 10523
rect 5816 10480 5868 10489
rect 6920 10480 6972 10532
rect 19892 10523 19944 10532
rect 19892 10489 19901 10523
rect 19901 10489 19935 10523
rect 19935 10489 19944 10523
rect 19892 10480 19944 10489
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 2872 10412 2924 10464
rect 3884 10412 3936 10464
rect 4896 10412 4948 10464
rect 7564 10455 7616 10464
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 21364 10616 21416 10668
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 23664 10659 23716 10668
rect 23664 10625 23673 10659
rect 23673 10625 23707 10659
rect 23707 10625 23716 10659
rect 23664 10616 23716 10625
rect 21640 10523 21692 10532
rect 21640 10489 21649 10523
rect 21649 10489 21683 10523
rect 21683 10489 21692 10523
rect 21640 10480 21692 10489
rect 20812 10412 20864 10464
rect 21548 10412 21600 10464
rect 23388 10480 23440 10532
rect 24308 10480 24360 10532
rect 26976 10616 27028 10668
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 27160 10548 27212 10600
rect 26700 10480 26752 10532
rect 22928 10412 22980 10464
rect 23756 10412 23808 10464
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 1676 10208 1728 10260
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 5816 10208 5868 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 9128 10208 9180 10260
rect 11336 10208 11388 10260
rect 18052 10208 18104 10260
rect 18328 10208 18380 10260
rect 19156 10208 19208 10260
rect 19432 10208 19484 10260
rect 19800 10251 19852 10260
rect 19800 10217 19809 10251
rect 19809 10217 19843 10251
rect 19843 10217 19852 10251
rect 19800 10208 19852 10217
rect 19984 10208 20036 10260
rect 21364 10251 21416 10260
rect 21364 10217 21373 10251
rect 21373 10217 21407 10251
rect 21407 10217 21416 10251
rect 21364 10208 21416 10217
rect 22008 10251 22060 10260
rect 22008 10217 22017 10251
rect 22017 10217 22051 10251
rect 22051 10217 22060 10251
rect 22008 10208 22060 10217
rect 22744 10251 22796 10260
rect 22744 10217 22753 10251
rect 22753 10217 22787 10251
rect 22787 10217 22796 10251
rect 22744 10208 22796 10217
rect 23388 10251 23440 10260
rect 23388 10217 23397 10251
rect 23397 10217 23431 10251
rect 23431 10217 23440 10251
rect 23388 10208 23440 10217
rect 26700 10208 26752 10260
rect 26976 10208 27028 10260
rect 4620 10183 4672 10192
rect 4620 10149 4629 10183
rect 4629 10149 4663 10183
rect 4663 10149 4672 10183
rect 4620 10140 4672 10149
rect 21456 10140 21508 10192
rect 21732 10140 21784 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2596 10072 2648 10124
rect 3792 10115 3844 10124
rect 3792 10081 3801 10115
rect 3801 10081 3835 10115
rect 3835 10081 3844 10115
rect 3792 10072 3844 10081
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 5080 10072 5132 10124
rect 7840 10072 7892 10124
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 23388 10072 23440 10124
rect 23664 10140 23716 10192
rect 23756 10115 23808 10124
rect 23756 10081 23790 10115
rect 23790 10081 23808 10115
rect 23756 10072 23808 10081
rect 26608 10072 26660 10124
rect 2780 9936 2832 9988
rect 4804 10004 4856 10056
rect 3424 9979 3476 9988
rect 3424 9945 3433 9979
rect 3433 9945 3467 9979
rect 3467 9945 3476 9979
rect 3424 9936 3476 9945
rect 2044 9868 2096 9920
rect 2320 9868 2372 9920
rect 4068 9868 4120 9920
rect 5080 9868 5132 9920
rect 8116 10004 8168 10056
rect 8484 10047 8536 10056
rect 8484 10013 8493 10047
rect 8493 10013 8527 10047
rect 8527 10013 8536 10047
rect 8484 10004 8536 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 22284 10047 22336 10056
rect 18512 10004 18564 10013
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 7196 9936 7248 9988
rect 21640 9979 21692 9988
rect 21640 9945 21649 9979
rect 21649 9945 21683 9979
rect 21683 9945 21692 9979
rect 21640 9936 21692 9945
rect 6276 9868 6328 9920
rect 24952 9868 25004 9920
rect 26976 9868 27028 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 3148 9664 3200 9716
rect 3424 9664 3476 9716
rect 8760 9664 8812 9716
rect 9220 9664 9272 9716
rect 4252 9596 4304 9648
rect 4988 9596 5040 9648
rect 5448 9639 5500 9648
rect 5448 9605 5457 9639
rect 5457 9605 5491 9639
rect 5491 9605 5500 9639
rect 5448 9596 5500 9605
rect 5540 9596 5592 9648
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 8392 9639 8444 9648
rect 2136 9460 2188 9512
rect 7012 9528 7064 9580
rect 8392 9605 8401 9639
rect 8401 9605 8435 9639
rect 8435 9605 8444 9639
rect 8392 9596 8444 9605
rect 8484 9596 8536 9648
rect 17500 9596 17552 9648
rect 18512 9664 18564 9716
rect 19156 9707 19208 9716
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 21548 9664 21600 9716
rect 26608 9664 26660 9716
rect 18144 9639 18196 9648
rect 18144 9605 18153 9639
rect 18153 9605 18187 9639
rect 18187 9605 18196 9639
rect 18144 9596 18196 9605
rect 19708 9639 19760 9648
rect 19708 9605 19717 9639
rect 19717 9605 19751 9639
rect 19751 9605 19760 9639
rect 19708 9596 19760 9605
rect 20352 9596 20404 9648
rect 23388 9596 23440 9648
rect 23848 9639 23900 9648
rect 23848 9605 23857 9639
rect 23857 9605 23891 9639
rect 23891 9605 23900 9639
rect 23848 9596 23900 9605
rect 7656 9528 7708 9580
rect 17040 9528 17092 9580
rect 18420 9528 18472 9580
rect 6736 9460 6788 9512
rect 8852 9460 8904 9512
rect 16856 9460 16908 9512
rect 19248 9528 19300 9580
rect 19800 9528 19852 9580
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 22284 9571 22336 9580
rect 20812 9528 20864 9537
rect 22284 9537 22293 9571
rect 22293 9537 22327 9571
rect 22327 9537 22336 9571
rect 22284 9528 22336 9537
rect 24952 9528 25004 9580
rect 20076 9460 20128 9469
rect 21824 9460 21876 9512
rect 26884 9596 26936 9648
rect 27436 9460 27488 9512
rect 3424 9392 3476 9444
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 8760 9392 8812 9401
rect 21456 9435 21508 9444
rect 21456 9401 21465 9435
rect 21465 9401 21499 9435
rect 21499 9401 21508 9435
rect 21456 9392 21508 9401
rect 23480 9392 23532 9444
rect 24216 9435 24268 9444
rect 24216 9401 24225 9435
rect 24225 9401 24259 9435
rect 24259 9401 24268 9435
rect 24216 9392 24268 9401
rect 1676 9324 1728 9376
rect 4988 9324 5040 9376
rect 5540 9324 5592 9376
rect 6276 9324 6328 9376
rect 7288 9324 7340 9376
rect 8116 9324 8168 9376
rect 8576 9324 8628 9376
rect 17960 9324 18012 9376
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 24492 9324 24544 9376
rect 26792 9324 26844 9376
rect 27804 9324 27856 9376
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 2044 9120 2096 9172
rect 2780 9120 2832 9172
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3792 9120 3844 9172
rect 5356 9120 5408 9172
rect 6920 9120 6972 9172
rect 8852 9120 8904 9172
rect 18328 9120 18380 9172
rect 18880 9120 18932 9172
rect 20076 9120 20128 9172
rect 21732 9163 21784 9172
rect 21732 9129 21741 9163
rect 21741 9129 21775 9163
rect 21775 9129 21784 9163
rect 21732 9120 21784 9129
rect 22100 9163 22152 9172
rect 22100 9129 22109 9163
rect 22109 9129 22143 9163
rect 22143 9129 22152 9163
rect 22100 9120 22152 9129
rect 24492 9163 24544 9172
rect 24492 9129 24501 9163
rect 24501 9129 24535 9163
rect 24535 9129 24544 9163
rect 24492 9120 24544 9129
rect 24860 9163 24912 9172
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 25044 9120 25096 9172
rect 26148 9120 26200 9172
rect 2596 9052 2648 9104
rect 17960 9052 18012 9104
rect 24216 9095 24268 9104
rect 24216 9061 24225 9095
rect 24225 9061 24259 9095
rect 24259 9061 24268 9095
rect 24216 9052 24268 9061
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 6276 8984 6328 9036
rect 18604 8984 18656 9036
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 2044 8916 2096 8968
rect 3516 8916 3568 8968
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5540 8916 5592 8968
rect 19248 8916 19300 8968
rect 23756 8916 23808 8968
rect 25228 8916 25280 8968
rect 3424 8891 3476 8900
rect 3424 8857 3433 8891
rect 3433 8857 3467 8891
rect 3467 8857 3476 8891
rect 3424 8848 3476 8857
rect 2872 8780 2924 8832
rect 5080 8823 5132 8832
rect 5080 8789 5089 8823
rect 5089 8789 5123 8823
rect 5123 8789 5132 8823
rect 5080 8780 5132 8789
rect 6736 8780 6788 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 26700 8823 26752 8832
rect 26700 8789 26709 8823
rect 26709 8789 26743 8823
rect 26743 8789 26752 8823
rect 26700 8780 26752 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 4068 8576 4120 8628
rect 4528 8576 4580 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 18880 8619 18932 8628
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 19248 8619 19300 8628
rect 19248 8585 19257 8619
rect 19257 8585 19291 8619
rect 19291 8585 19300 8619
rect 19248 8576 19300 8585
rect 25044 8576 25096 8628
rect 25228 8619 25280 8628
rect 25228 8585 25237 8619
rect 25237 8585 25271 8619
rect 25271 8585 25280 8619
rect 25228 8576 25280 8585
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 26516 8576 26568 8628
rect 27712 8619 27764 8628
rect 27712 8585 27721 8619
rect 27721 8585 27755 8619
rect 27755 8585 27764 8619
rect 27712 8576 27764 8585
rect 1860 8508 1912 8560
rect 4620 8551 4672 8560
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 4620 8517 4629 8551
rect 4629 8517 4663 8551
rect 4663 8517 4672 8551
rect 4620 8508 4672 8517
rect 3516 8440 3568 8492
rect 4712 8440 4764 8492
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 25136 8508 25188 8560
rect 26608 8551 26660 8560
rect 26608 8517 26617 8551
rect 26617 8517 26651 8551
rect 26651 8517 26660 8551
rect 26608 8508 26660 8517
rect 5816 8440 5868 8492
rect 6736 8440 6788 8492
rect 1768 8372 1820 8424
rect 2596 8372 2648 8424
rect 2780 8372 2832 8424
rect 3240 8372 3292 8424
rect 3792 8372 3844 8424
rect 5356 8372 5408 8424
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 25688 8440 25740 8492
rect 7196 8372 7248 8381
rect 25320 8415 25372 8424
rect 25320 8381 25329 8415
rect 25329 8381 25363 8415
rect 25363 8381 25372 8415
rect 25320 8372 25372 8381
rect 27252 8508 27304 8560
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 3700 8304 3752 8356
rect 5540 8304 5592 8356
rect 5908 8304 5960 8356
rect 6276 8304 6328 8356
rect 6920 8304 6972 8356
rect 1768 8236 1820 8288
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 5816 8236 5868 8288
rect 6736 8236 6788 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1400 8032 1452 8084
rect 1768 8032 1820 8084
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 2964 8032 3016 8084
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 4068 8032 4120 8084
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 5080 8032 5132 8084
rect 5724 8032 5776 8084
rect 24768 8032 24820 8084
rect 25596 8032 25648 8084
rect 26332 8032 26384 8084
rect 26516 8032 26568 8084
rect 2320 7964 2372 8016
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2044 7896 2096 7905
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2688 7828 2740 7880
rect 1400 7692 1452 7744
rect 1584 7692 1636 7744
rect 2688 7692 2740 7744
rect 3700 7964 3752 8016
rect 4160 7896 4212 7948
rect 4896 7896 4948 7948
rect 5540 7896 5592 7948
rect 6368 7896 6420 7948
rect 7840 7896 7892 7948
rect 25320 7939 25372 7948
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 27068 7896 27120 7948
rect 4988 7828 5040 7880
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 6920 7828 6972 7880
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 4988 7692 5040 7744
rect 5356 7692 5408 7744
rect 26332 7692 26384 7744
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 2044 7488 2096 7540
rect 2412 7488 2464 7540
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 4436 7488 4488 7540
rect 5724 7488 5776 7540
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 25320 7531 25372 7540
rect 25320 7497 25329 7531
rect 25329 7497 25363 7531
rect 25363 7497 25372 7531
rect 25320 7488 25372 7497
rect 27068 7488 27120 7540
rect 1584 7463 1636 7472
rect 1584 7429 1593 7463
rect 1593 7429 1627 7463
rect 1627 7429 1636 7463
rect 1584 7420 1636 7429
rect 2228 7420 2280 7472
rect 4988 7420 5040 7472
rect 2964 7395 3016 7404
rect 2964 7361 2973 7395
rect 2973 7361 3007 7395
rect 3007 7361 3016 7395
rect 2964 7352 3016 7361
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 27712 7463 27764 7472
rect 27712 7429 27721 7463
rect 27721 7429 27755 7463
rect 27755 7429 27764 7463
rect 27712 7420 27764 7429
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 3056 7284 3108 7336
rect 3424 7284 3476 7336
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 26424 7327 26476 7336
rect 26424 7293 26433 7327
rect 26433 7293 26467 7327
rect 26467 7293 26476 7327
rect 26424 7284 26476 7293
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 2872 7148 2924 7200
rect 3792 7148 3844 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 26884 7148 26936 7200
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 3424 6987 3476 6996
rect 3424 6953 3433 6987
rect 3433 6953 3467 6987
rect 3467 6953 3476 6987
rect 3424 6944 3476 6953
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 4988 6987 5040 6996
rect 4988 6953 4997 6987
rect 4997 6953 5031 6987
rect 5031 6953 5040 6987
rect 4988 6944 5040 6953
rect 5448 6987 5500 6996
rect 5448 6953 5457 6987
rect 5457 6953 5491 6987
rect 5491 6953 5500 6987
rect 5448 6944 5500 6953
rect 7196 6987 7248 6996
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 1860 6808 1912 6860
rect 2964 6876 3016 6928
rect 3516 6808 3568 6860
rect 4344 6808 4396 6860
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5540 6876 5592 6928
rect 7472 6876 7524 6928
rect 8300 6876 8352 6928
rect 5816 6851 5868 6860
rect 5356 6808 5408 6817
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 6460 6808 6512 6860
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 2596 6740 2648 6792
rect 2780 6740 2832 6792
rect 5540 6740 5592 6792
rect 6276 6740 6328 6792
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 2504 6672 2556 6724
rect 4160 6604 4212 6656
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1400 6400 1452 6452
rect 2688 6400 2740 6452
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 4344 6400 4396 6452
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 7472 6400 7524 6452
rect 26608 6443 26660 6452
rect 26608 6409 26617 6443
rect 26617 6409 26651 6443
rect 26651 6409 26660 6443
rect 26608 6400 26660 6409
rect 1584 6375 1636 6384
rect 1584 6341 1593 6375
rect 1593 6341 1627 6375
rect 1627 6341 1636 6375
rect 1584 6332 1636 6341
rect 2044 6375 2096 6384
rect 2044 6341 2053 6375
rect 2053 6341 2087 6375
rect 2087 6341 2096 6375
rect 2044 6332 2096 6341
rect 26516 6332 26568 6384
rect 3516 6239 3568 6248
rect 3516 6205 3525 6239
rect 3525 6205 3559 6239
rect 3559 6205 3568 6239
rect 3516 6196 3568 6205
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 27160 6264 27212 6316
rect 3608 6196 3660 6205
rect 2228 6060 2280 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2136 5856 2188 5908
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 2320 5788 2372 5840
rect 1768 5720 1820 5772
rect 2504 5763 2556 5772
rect 2504 5729 2513 5763
rect 2513 5729 2547 5763
rect 2547 5729 2556 5763
rect 2504 5720 2556 5729
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 26700 5627 26752 5636
rect 26700 5593 26709 5627
rect 26709 5593 26743 5627
rect 26743 5593 26752 5627
rect 26700 5584 26752 5593
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 26516 5312 26568 5364
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 1768 4768 1820 4820
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2044 2932 2096 2984
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 7196 2499 7248 2508
rect 7196 2465 7230 2499
rect 7230 2465 7248 2499
rect 7196 2456 7248 2465
rect 4988 2252 5040 2304
rect 5724 2252 5776 2304
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 938 23520 994 24000
rect 2778 23520 2834 24000
rect 2962 23624 3018 23633
rect 2962 23559 3018 23568
rect 952 20602 980 23520
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1122 15328 1178 15337
rect 1122 15263 1178 15272
rect 1136 11286 1164 15263
rect 1216 14816 1268 14822
rect 1216 14758 1268 14764
rect 1228 12714 1256 14758
rect 1412 12730 1440 20431
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 18834 1716 19654
rect 2136 19236 2188 19242
rect 2136 19178 2188 19184
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1504 17202 1532 17614
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1504 16522 1532 17138
rect 1492 16516 1544 16522
rect 1492 16458 1544 16464
rect 1596 16250 1624 18226
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 16794 1716 18158
rect 1780 16833 1808 19110
rect 1964 18290 1992 19110
rect 2148 18766 2176 19178
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 18290 2176 18702
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2148 18170 2176 18226
rect 2056 18142 2176 18170
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1872 17134 1900 18022
rect 2056 17814 2084 18142
rect 2044 17808 2096 17814
rect 2044 17750 2096 17756
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 1766 16824 1822 16833
rect 1676 16788 1728 16794
rect 1766 16759 1822 16768
rect 1676 16730 1728 16736
rect 2332 16590 2360 17070
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 2332 16114 2360 16526
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1596 15366 1624 15846
rect 1780 15706 1808 15982
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1504 14482 1532 14894
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 13394 1532 14418
rect 1596 13433 1624 15302
rect 2148 14074 2176 15506
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2240 14822 2268 15438
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2226 14104 2282 14113
rect 2136 14068 2188 14074
rect 2226 14039 2282 14048
rect 2136 14010 2188 14016
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1860 13456 1912 13462
rect 1582 13424 1638 13433
rect 1492 13388 1544 13394
rect 1860 13398 1912 13404
rect 1582 13359 1638 13368
rect 1492 13330 1544 13336
rect 1216 12708 1268 12714
rect 1412 12702 1624 12730
rect 1216 12650 1268 12656
rect 1228 12345 1256 12650
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1214 12336 1270 12345
rect 1214 12271 1270 12280
rect 1124 11280 1176 11286
rect 1124 11222 1176 11228
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 8090 1440 10066
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1412 7342 1440 7686
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 6458 1440 6802
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1504 3913 1532 12582
rect 1596 7750 1624 12702
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1674 10296 1730 10305
rect 1674 10231 1676 10240
rect 1728 10231 1730 10240
rect 1676 10202 1728 10208
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1584 7472 1636 7478
rect 1582 7440 1584 7449
rect 1636 7440 1638 7449
rect 1582 7375 1638 7384
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 6730 1624 6831
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1584 6384 1636 6390
rect 1582 6352 1584 6361
rect 1636 6352 1638 6361
rect 1582 6287 1638 6296
rect 1582 5672 1638 5681
rect 1582 5607 1584 5616
rect 1636 5607 1638 5616
rect 1584 5578 1636 5584
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 5030 1624 5063
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1688 4457 1716 9318
rect 1780 8430 1808 10406
rect 1872 8566 1900 13398
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1780 8090 1808 8230
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1766 7304 1822 7313
rect 1766 7239 1822 7248
rect 1780 5778 1808 7239
rect 1872 6866 1900 8502
rect 1964 8498 1992 13670
rect 2042 13560 2098 13569
rect 2042 13495 2098 13504
rect 2056 10418 2084 13495
rect 2134 12608 2190 12617
rect 2134 12543 2190 12552
rect 2148 11762 2176 12543
rect 2240 12374 2268 14039
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 2240 11898 2268 12310
rect 2332 12102 2360 13670
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2332 11354 2360 12038
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2240 10674 2268 11018
rect 2332 10810 2360 11154
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2134 10568 2190 10577
rect 2134 10503 2136 10512
rect 2188 10503 2190 10512
rect 2136 10474 2188 10480
rect 2056 10390 2176 10418
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9178 2084 9862
rect 2148 9518 2176 10390
rect 2332 9926 2360 10610
rect 2424 10266 2452 20198
rect 2792 18834 2820 23520
rect 2976 22166 3004 23559
rect 4618 23520 4674 24000
rect 6550 23520 6606 24000
rect 8390 23520 8446 24000
rect 10230 23520 10286 24000
rect 12162 23520 12218 24000
rect 14002 23520 14058 24000
rect 15934 23520 15990 24000
rect 17774 23520 17830 24000
rect 19614 23520 19670 24000
rect 21546 23520 21602 24000
rect 23386 23520 23442 24000
rect 25042 23624 25098 23633
rect 25042 23559 25098 23568
rect 3330 23080 3386 23089
rect 3330 23015 3386 23024
rect 3344 22574 3372 23015
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3146 22400 3202 22409
rect 3146 22335 3202 22344
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 2962 19544 3018 19553
rect 2962 19479 3018 19488
rect 2976 19174 3004 19479
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2700 18714 2728 18770
rect 2700 18686 2820 18714
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2608 16114 2636 16662
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2608 16017 2636 16050
rect 2700 16046 2728 17546
rect 2792 16794 2820 18686
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2976 18222 3004 18566
rect 3068 18426 3096 19246
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17882 2912 18022
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2964 17808 3016 17814
rect 2964 17750 3016 17756
rect 2976 17338 3004 17750
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2778 16688 2834 16697
rect 2778 16623 2780 16632
rect 2832 16623 2834 16632
rect 2780 16594 2832 16600
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2688 16040 2740 16046
rect 2594 16008 2650 16017
rect 2688 15982 2740 15988
rect 2594 15943 2650 15952
rect 2792 15706 2820 16458
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 14890 2544 15438
rect 2792 15094 2820 15642
rect 2884 15366 2912 15914
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 2516 14618 2544 14826
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2608 13705 2636 13806
rect 2792 13734 2820 14418
rect 2884 13977 2912 15302
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 3068 14074 3096 15030
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2870 13968 2926 13977
rect 2870 13903 2926 13912
rect 2964 13932 3016 13938
rect 2780 13728 2832 13734
rect 2594 13696 2650 13705
rect 2780 13670 2832 13676
rect 2594 13631 2650 13640
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2516 12918 2544 13330
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 2516 12442 2544 12854
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2516 11830 2544 12378
rect 2608 11898 2636 13631
rect 2792 13190 2820 13670
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 12764 2820 13126
rect 2884 12986 2912 13903
rect 2964 13874 3016 13880
rect 2976 13190 3004 13874
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2976 12782 3004 13126
rect 2700 12736 2820 12764
rect 2964 12776 3016 12782
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2594 11248 2650 11257
rect 2594 11183 2596 11192
rect 2648 11183 2650 11192
rect 2596 11154 2648 11160
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2608 10130 2636 11154
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2608 9761 2636 10066
rect 2594 9752 2650 9761
rect 2594 9687 2650 9696
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2056 8974 2084 9114
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2608 8634 2636 9046
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2502 8120 2558 8129
rect 2136 8084 2188 8090
rect 2502 8055 2558 8064
rect 2136 8026 2188 8032
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2056 7546 2084 7890
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 2042 6488 2098 6497
rect 2042 6423 2098 6432
rect 2056 6390 2084 6423
rect 2044 6384 2096 6390
rect 2044 6326 2096 6332
rect 2148 5914 2176 8026
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7478 2268 7822
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1780 4826 1808 5714
rect 2042 5264 2098 5273
rect 2042 5199 2044 5208
rect 2096 5199 2098 5208
rect 2044 5170 2096 5176
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1674 4448 1730 4457
rect 1674 4383 1730 4392
rect 2042 4040 2098 4049
rect 2042 3975 2098 3984
rect 1490 3904 1546 3913
rect 1490 3839 1546 3848
rect 2056 3194 2084 3975
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2689 1624 2790
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 2240 377 2268 6054
rect 2332 5846 2360 7958
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2424 5914 2452 7482
rect 2516 6730 2544 8055
rect 2608 6798 2636 8366
rect 2700 7886 2728 12736
rect 2964 12718 3016 12724
rect 2976 12594 3004 12718
rect 2792 12566 3004 12594
rect 2792 10674 2820 12566
rect 2976 12442 3004 12566
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2870 12336 2926 12345
rect 2870 12271 2872 12280
rect 2924 12271 2926 12280
rect 2872 12242 2924 12248
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11762 3004 12174
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 11150 3004 11698
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 3160 11098 3188 22335
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 4080 20806 4108 21791
rect 4434 21312 4490 21321
rect 4434 21247 4490 21256
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3606 20632 3662 20641
rect 3606 20567 3662 20576
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3252 18970 3280 19110
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3252 18222 3280 18906
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3344 16250 3372 18566
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3330 15872 3386 15881
rect 3330 15807 3386 15816
rect 3344 14113 3372 15807
rect 3330 14104 3386 14113
rect 3330 14039 3386 14048
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 3252 12374 3280 13942
rect 3436 12424 3464 18770
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3528 18358 3556 18566
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3528 18086 3556 18294
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3528 16522 3556 16934
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 3516 15904 3568 15910
rect 3620 15892 3648 20567
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4172 19258 4200 20334
rect 3988 19230 4200 19258
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3896 17134 3924 17614
rect 3884 17128 3936 17134
rect 3790 17096 3846 17105
rect 3884 17070 3936 17076
rect 3790 17031 3846 17040
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3712 16114 3740 16526
rect 3804 16153 3832 17031
rect 3882 16960 3938 16969
rect 3882 16895 3938 16904
rect 3790 16144 3846 16153
rect 3700 16108 3752 16114
rect 3790 16079 3846 16088
rect 3700 16050 3752 16056
rect 3568 15864 3648 15892
rect 3516 15846 3568 15852
rect 3712 15706 3740 16050
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3712 15162 3740 15642
rect 3804 15162 3832 15846
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3896 15042 3924 16895
rect 3620 15014 3924 15042
rect 3514 14512 3570 14521
rect 3514 14447 3570 14456
rect 3344 12396 3464 12424
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3160 11070 3280 11098
rect 2870 10840 2926 10849
rect 2870 10775 2872 10784
rect 2924 10775 2926 10784
rect 2872 10746 2924 10752
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2792 9178 2820 9930
rect 2884 9178 2912 10406
rect 3160 9722 3188 10610
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2778 9072 2834 9081
rect 2778 9007 2780 9016
rect 2832 9007 2834 9016
rect 2780 8978 2832 8984
rect 2792 8922 2820 8978
rect 2792 8894 3004 8922
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2700 6458 2728 7686
rect 2792 6798 2820 8366
rect 2884 7206 2912 8774
rect 2976 8090 3004 8894
rect 3252 8430 3280 11070
rect 3344 10305 3372 12396
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 11286 3464 11766
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3330 10296 3386 10305
rect 3330 10231 3386 10240
rect 3436 9994 3464 10474
rect 3528 10033 3556 14447
rect 3620 12306 3648 15014
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14618 3740 14758
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3804 13682 3832 14894
rect 3884 14272 3936 14278
rect 3882 14240 3884 14249
rect 3936 14240 3938 14249
rect 3882 14175 3938 14184
rect 3896 13938 3924 14175
rect 3988 14074 4016 19230
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4066 18320 4122 18329
rect 4066 18255 4122 18264
rect 4080 14958 4108 18255
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4172 14385 4200 18566
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4158 14376 4214 14385
rect 4158 14311 4214 14320
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3976 13728 4028 13734
rect 3804 13654 3924 13682
rect 3976 13670 4028 13676
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3712 12986 3740 13398
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3620 11898 3648 12242
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3620 10810 3648 11222
rect 3896 11218 3924 13654
rect 3988 13530 4016 13670
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4080 11665 4108 14214
rect 4172 13870 4200 14311
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4264 12617 4292 18022
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4356 17134 4384 17818
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4448 16946 4476 21247
rect 4632 19553 4660 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 4988 20528 5040 20534
rect 4986 20496 4988 20505
rect 5040 20496 5042 20505
rect 4986 20431 5042 20440
rect 4618 19544 4674 19553
rect 4618 19479 4674 19488
rect 4802 19272 4858 19281
rect 4802 19207 4858 19216
rect 4618 17912 4674 17921
rect 4618 17847 4674 17856
rect 4356 16918 4476 16946
rect 4356 14793 4384 16918
rect 4434 16824 4490 16833
rect 4434 16759 4436 16768
rect 4488 16759 4490 16768
rect 4436 16730 4488 16736
rect 4448 16250 4476 16730
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4540 15910 4568 16526
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4434 15600 4490 15609
rect 4434 15535 4490 15544
rect 4342 14784 4398 14793
rect 4342 14719 4398 14728
rect 4356 13938 4384 14719
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4250 12608 4306 12617
rect 4250 12543 4306 12552
rect 4448 12345 4476 15535
rect 4540 13326 4568 15846
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4632 13190 4660 17847
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4724 15366 4752 15982
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4724 14890 4752 15302
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4816 14482 4844 19207
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4908 18222 4936 18294
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4816 14074 4844 14418
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4908 13410 4936 18158
rect 4988 18080 5040 18086
rect 4986 18048 4988 18057
rect 5040 18048 5042 18057
rect 4986 17983 5042 17992
rect 5092 17746 5120 18226
rect 5184 18222 5212 18702
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5092 17338 5120 17682
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5078 16416 5134 16425
rect 5078 16351 5134 16360
rect 5092 15978 5120 16351
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 5184 15638 5212 18158
rect 5276 17882 5304 18770
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5368 18154 5396 18294
rect 5736 18193 5764 20742
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 6564 20505 6592 23520
rect 8404 23474 8432 23520
rect 8312 23446 8432 23474
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 6550 20496 6606 20505
rect 6550 20431 6606 20440
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 6734 19136 6790 19145
rect 6734 19071 6790 19080
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5722 18184 5778 18193
rect 5356 18148 5408 18154
rect 5722 18119 5778 18128
rect 5356 18090 5408 18096
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5276 16250 5304 17818
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5552 16794 5580 17274
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5000 14958 5028 15302
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 5000 14618 5028 14894
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4724 13382 4936 13410
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4724 13002 4752 13382
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4540 12974 4752 13002
rect 4434 12336 4490 12345
rect 4356 12294 4434 12322
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3698 10568 3754 10577
rect 3698 10503 3754 10512
rect 3514 10024 3570 10033
rect 3424 9988 3476 9994
rect 3514 9959 3570 9968
rect 3424 9930 3476 9936
rect 3436 9722 3464 9930
rect 3606 9752 3662 9761
rect 3424 9716 3476 9722
rect 3606 9687 3662 9696
rect 3424 9658 3476 9664
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3436 8906 3464 9386
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3528 8498 3556 8910
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2976 6934 3004 7346
rect 3068 7342 3096 8230
rect 3528 8090 3556 8434
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3436 7002 3464 7278
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 3146 6896 3202 6905
rect 3146 6831 3202 6840
rect 3516 6860 3568 6866
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 3160 6458 3188 6831
rect 3516 6802 3568 6808
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3528 6254 3556 6802
rect 3620 6254 3648 9687
rect 3712 8362 3740 10503
rect 3896 10470 3924 11154
rect 3884 10464 3936 10470
rect 4080 10441 4108 11290
rect 4264 11121 4292 12038
rect 4250 11112 4306 11121
rect 4250 11047 4306 11056
rect 3884 10406 3936 10412
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 4068 10124 4120 10130
rect 4120 10084 4292 10112
rect 4068 10066 4120 10072
rect 3804 9178 3832 10066
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4080 9353 4108 9862
rect 4264 9654 4292 10084
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3790 8936 3846 8945
rect 3790 8871 3846 8880
rect 3804 8430 3832 8871
rect 4250 8664 4306 8673
rect 4068 8628 4120 8634
rect 4250 8599 4306 8608
rect 4068 8570 4120 8576
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3712 8022 3740 8298
rect 4080 8090 4108 8570
rect 4264 8090 4292 8599
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7546 4200 7890
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3804 7002 3832 7142
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 4356 6866 4384 12294
rect 4434 12271 4490 12280
rect 4540 12209 4568 12974
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4526 12200 4582 12209
rect 4526 12135 4582 12144
rect 4540 11558 4568 12135
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11626 4752 12038
rect 4816 11898 4844 12378
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4724 10810 4752 11562
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4448 7546 4476 8978
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8634 4568 8910
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4632 8566 4660 10134
rect 4816 10062 4844 11222
rect 4908 10470 4936 13262
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4724 8498 4752 8910
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4908 7954 4936 10406
rect 5000 9654 5028 14010
rect 5092 13938 5120 14826
rect 5184 14822 5212 15574
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5184 12986 5212 14758
rect 5552 14090 5580 16594
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5644 15910 5672 16526
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5644 15609 5672 15846
rect 5630 15600 5686 15609
rect 5630 15535 5686 15544
rect 5736 15450 5764 18119
rect 6472 18086 6500 18770
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 6380 16046 6408 17478
rect 6472 16250 6500 18022
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5644 15422 5764 15450
rect 5644 14958 5672 15422
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5736 14550 5764 15302
rect 5828 15065 5856 15914
rect 6552 15904 6604 15910
rect 6550 15872 6552 15881
rect 6604 15872 6606 15881
rect 6550 15807 6606 15816
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 5814 15056 5870 15065
rect 5814 14991 5870 15000
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5632 14272 5684 14278
rect 5736 14249 5764 14486
rect 5632 14214 5684 14220
rect 5722 14240 5778 14249
rect 5460 14062 5580 14090
rect 5264 13728 5316 13734
rect 5460 13682 5488 14062
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5264 13670 5316 13676
rect 5276 13326 5304 13670
rect 5368 13654 5488 13682
rect 5368 13462 5396 13654
rect 5448 13524 5500 13530
rect 5552 13512 5580 13942
rect 5644 13734 5672 14214
rect 5722 14175 5778 14184
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 13569 5672 13670
rect 5500 13484 5580 13512
rect 5630 13560 5686 13569
rect 5736 13530 5764 14175
rect 5828 13682 5856 14894
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6184 14476 6236 14482
rect 6236 14436 6316 14464
rect 6184 14418 6236 14424
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5828 13654 5948 13682
rect 5814 13560 5870 13569
rect 5630 13495 5686 13504
rect 5724 13524 5776 13530
rect 5448 13466 5500 13472
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5264 13320 5316 13326
rect 5262 13288 5264 13297
rect 5448 13320 5500 13326
rect 5316 13288 5318 13297
rect 5448 13262 5500 13268
rect 5262 13223 5318 13232
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 5092 11268 5120 12310
rect 5184 11393 5212 12582
rect 5170 11384 5226 11393
rect 5170 11319 5226 11328
rect 5092 11240 5212 11268
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10130 5120 10950
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9926 5120 10066
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5092 9466 5120 9862
rect 5000 9438 5120 9466
rect 5000 9382 5028 9438
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5000 7886 5028 9318
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 8498 5120 8774
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 8090 5120 8434
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5000 7750 5028 7822
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 5000 7478 5028 7686
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 5000 7002 5028 7414
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5184 6905 5212 11240
rect 5276 7342 5304 13126
rect 5460 12986 5488 13262
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5644 12753 5672 13495
rect 5814 13495 5870 13504
rect 5724 13466 5776 13472
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5630 12744 5686 12753
rect 5630 12679 5686 12688
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5460 12374 5488 12582
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5644 11558 5672 12174
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5368 9178 5396 11018
rect 5552 10826 5580 11290
rect 5460 10810 5580 10826
rect 5448 10804 5580 10810
rect 5500 10798 5580 10804
rect 5448 10746 5500 10752
rect 5446 9888 5502 9897
rect 5446 9823 5502 9832
rect 5460 9654 5488 9823
rect 5552 9654 5580 10798
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5368 8430 5396 9114
rect 5552 8974 5580 9318
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5446 8392 5502 8401
rect 5552 8362 5580 8910
rect 5446 8327 5502 8336
rect 5540 8356 5592 8362
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7410 5396 7686
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5460 7002 5488 8327
rect 5540 8298 5592 8304
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5552 6934 5580 7890
rect 5540 6928 5592 6934
rect 5170 6896 5226 6905
rect 4344 6860 4396 6866
rect 5540 6870 5592 6876
rect 5170 6831 5226 6840
rect 5356 6860 5408 6866
rect 4344 6802 4396 6808
rect 5356 6802 5408 6808
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 3516 6248 3568 6254
rect 3514 6216 3516 6225
rect 3608 6248 3660 6254
rect 3568 6216 3570 6225
rect 3608 6190 3660 6196
rect 3514 6151 3570 6160
rect 3620 5914 3648 6190
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2502 5808 2558 5817
rect 2502 5743 2504 5752
rect 2556 5743 2558 5752
rect 2504 5714 2556 5720
rect 2516 5370 2544 5714
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2700 1465 2728 5510
rect 3804 3369 3832 6054
rect 4172 4706 4200 6598
rect 4356 6458 4384 6802
rect 5368 6497 5396 6802
rect 5540 6792 5592 6798
rect 5644 6780 5672 11494
rect 5736 8090 5764 13262
rect 5828 13161 5856 13495
rect 5920 13326 5948 13654
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6012 13258 6040 13874
rect 6288 13870 6316 14436
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6182 13696 6238 13705
rect 6182 13631 6238 13640
rect 6196 13530 6224 13631
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6288 13326 6316 13806
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5814 13152 5870 13161
rect 5814 13087 5870 13096
rect 5828 12238 5856 13087
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6288 12986 6316 13262
rect 6366 13152 6422 13161
rect 6366 13087 6422 13096
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6274 12880 6330 12889
rect 6274 12815 6330 12824
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5920 12084 5948 12242
rect 5828 12056 5948 12084
rect 5828 11626 5856 12056
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 6288 11354 6316 12815
rect 6380 12442 6408 13087
rect 6472 12850 6500 13398
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 10538 5856 11154
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 5816 10532 5868 10538
rect 5816 10474 5868 10480
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5828 8498 5856 10202
rect 6288 9926 6316 11086
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 6288 9382 6316 9862
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6288 8362 6316 8978
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5736 7546 5764 8026
rect 5828 7886 5856 8230
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5920 7732 5948 8298
rect 5828 7704 5948 7732
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5828 7426 5856 7704
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 5592 6752 5672 6780
rect 5736 7398 5856 7426
rect 5540 6734 5592 6740
rect 5354 6488 5410 6497
rect 4344 6452 4396 6458
rect 5552 6458 5580 6734
rect 5354 6423 5410 6432
rect 5540 6452 5592 6458
rect 4344 6394 4396 6400
rect 5540 6394 5592 6400
rect 4080 4678 4200 4706
rect 3790 3360 3846 3369
rect 3790 3295 3846 3304
rect 4080 2145 4108 4678
rect 5736 2310 5764 7398
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5828 6118 5856 6802
rect 6288 6798 6316 8298
rect 6380 7954 6408 12242
rect 6472 12238 6500 12786
rect 6564 12714 6592 14826
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 12102 6500 12174
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6472 6866 6500 11494
rect 6564 7546 6592 12650
rect 6656 12306 6684 17002
rect 6748 16794 6776 19071
rect 7656 18080 7708 18086
rect 7470 18048 7526 18057
rect 7656 18022 7708 18028
rect 7470 17983 7526 17992
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6840 16674 6868 16934
rect 6932 16794 6960 17478
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7484 16726 7512 17983
rect 7668 16998 7696 18022
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7760 17241 7788 17614
rect 7746 17232 7802 17241
rect 7746 17167 7802 17176
rect 7760 17066 7788 17167
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7472 16720 7524 16726
rect 6840 16646 6960 16674
rect 7472 16662 7524 16668
rect 6932 16590 6960 16646
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6840 15706 6868 15982
rect 6932 15706 6960 16526
rect 7484 16046 7512 16662
rect 7668 16590 7696 16934
rect 7746 16688 7802 16697
rect 7746 16623 7802 16632
rect 7760 16590 7788 16623
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7208 15473 7236 15846
rect 7194 15464 7250 15473
rect 7194 15399 7250 15408
rect 7760 15366 7788 16526
rect 6920 15360 6972 15366
rect 6840 15308 6920 15314
rect 6840 15302 6972 15308
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 6840 15286 6960 15302
rect 6840 15162 6868 15286
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14618 6868 14758
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13462 6776 14214
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6840 13138 6868 13942
rect 7208 13870 7236 14554
rect 7286 14240 7342 14249
rect 7286 14175 7342 14184
rect 7300 14074 7328 14175
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7300 13870 7328 14010
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7576 13569 7604 14962
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7562 13560 7618 13569
rect 7562 13495 7618 13504
rect 7668 13433 7696 14758
rect 7654 13424 7710 13433
rect 7654 13359 7710 13368
rect 7288 13184 7340 13190
rect 6840 13110 7052 13138
rect 7288 13126 7340 13132
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6656 11082 6684 12038
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6748 9518 6776 12106
rect 6840 9654 6868 12650
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12238 6960 12582
rect 7024 12374 7052 13110
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 7116 11558 7144 12242
rect 7104 11552 7156 11558
rect 7102 11520 7104 11529
rect 7156 11520 7158 11529
rect 7102 11455 7158 11464
rect 6918 11384 6974 11393
rect 6974 11328 7052 11336
rect 6918 11319 6920 11328
rect 6972 11308 7052 11328
rect 6920 11290 6972 11296
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6932 9178 6960 10474
rect 7024 9586 7052 11308
rect 7300 11286 7328 13126
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7392 12102 7420 12786
rect 7668 12782 7696 13359
rect 7760 13161 7788 15302
rect 7746 13152 7802 13161
rect 7746 13087 7802 13096
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7852 12442 7880 20198
rect 7944 17338 7972 22510
rect 8312 20618 8340 23446
rect 8220 20602 8340 20618
rect 10244 20602 10272 23520
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 8208 20596 8340 20602
rect 8260 20590 8340 20596
rect 10232 20596 10284 20602
rect 8208 20538 8260 20544
rect 10232 20538 10284 20544
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18834 8616 19110
rect 8772 18970 8800 19382
rect 9048 19174 9076 19654
rect 9586 19544 9642 19553
rect 9586 19479 9642 19488
rect 9600 19446 9628 19479
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9036 19168 9088 19174
rect 9034 19136 9036 19145
rect 9088 19136 9090 19145
rect 9034 19071 9090 19080
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8496 18086 8524 18158
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8022 17640 8078 17649
rect 8022 17575 8078 17584
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7944 16454 7972 17070
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 8036 15337 8064 17575
rect 8128 17542 8156 18022
rect 8298 17912 8354 17921
rect 8298 17847 8354 17856
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8312 16794 8340 17847
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8404 17513 8432 17682
rect 8390 17504 8446 17513
rect 8390 17439 8446 17448
rect 8404 17338 8432 17439
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8312 16697 8340 16730
rect 8298 16688 8354 16697
rect 8298 16623 8354 16632
rect 8312 16250 8340 16623
rect 8496 16454 8524 18022
rect 9048 17882 9076 18770
rect 9508 18426 9536 19314
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9600 19122 9628 19178
rect 9600 19094 9812 19122
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9692 17882 9720 18770
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 17542 8616 17614
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 17066 8616 17478
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 16590 8616 17002
rect 9416 16998 9444 17750
rect 9784 17338 9812 19094
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9876 16998 9904 17614
rect 9404 16992 9456 16998
rect 9864 16992 9916 16998
rect 9404 16934 9456 16940
rect 9862 16960 9864 16969
rect 9916 16960 9918 16969
rect 9862 16895 9918 16904
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8496 16046 8524 16390
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8116 15360 8168 15366
rect 8022 15328 8078 15337
rect 8116 15302 8168 15308
rect 8022 15263 8078 15272
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 14074 7972 14214
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8128 13938 8156 15302
rect 8220 15162 8248 15438
rect 8404 15201 8432 15506
rect 8496 15366 8524 15982
rect 8588 15502 8616 16526
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8680 15978 8708 16390
rect 9876 16250 9904 16526
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 8942 16144 8998 16153
rect 8942 16079 8998 16088
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8390 15192 8446 15201
rect 8208 15156 8260 15162
rect 8390 15127 8446 15136
rect 8208 15098 8260 15104
rect 8404 15042 8432 15127
rect 8220 15026 8432 15042
rect 8680 15026 8708 15914
rect 8208 15020 8432 15026
rect 8260 15014 8432 15020
rect 8668 15020 8720 15026
rect 8208 14962 8260 14968
rect 8668 14962 8720 14968
rect 8680 14074 8708 14962
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13530 8524 13806
rect 8864 13530 8892 14350
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8298 13288 8354 13297
rect 8298 13223 8354 13232
rect 8312 12986 8340 13223
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11762 7696 12038
rect 7760 11898 7788 12174
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11354 7512 11494
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 9994 7236 10950
rect 7300 10674 7328 11222
rect 7484 10810 7512 11290
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7470 10704 7526 10713
rect 7288 10668 7340 10674
rect 7470 10639 7526 10648
rect 7656 10668 7708 10674
rect 7288 10610 7340 10616
rect 7484 10606 7512 10639
rect 7656 10610 7708 10616
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 10033 7604 10406
rect 7668 10266 7696 10610
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7286 10024 7342 10033
rect 7196 9988 7248 9994
rect 7286 9959 7342 9968
rect 7562 10024 7618 10033
rect 7562 9959 7618 9968
rect 7196 9930 7248 9936
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7300 9382 7328 9959
rect 7668 9586 7696 10202
rect 7838 10160 7894 10169
rect 7838 10095 7840 10104
rect 7892 10095 7894 10104
rect 7840 10066 7892 10072
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6748 8498 6776 8774
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6748 8294 6776 8434
rect 7196 8424 7248 8430
rect 7194 8392 7196 8401
rect 7248 8392 7250 8401
rect 6840 8362 6960 8378
rect 6840 8356 6972 8362
rect 6840 8350 6920 8356
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6840 7546 6868 8350
rect 7194 8327 7250 8336
rect 6920 8298 6972 8304
rect 7300 7886 7328 9318
rect 7852 8838 7880 10066
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9382 8156 9998
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8312 9081 8340 12582
rect 8496 11694 8524 12854
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 9654 8432 11562
rect 8496 11558 8524 11630
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11218 8524 11494
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8680 10810 8708 12650
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 11694 8800 12038
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8772 11082 8800 11630
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8864 10674 8892 10950
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8956 10606 8984 16079
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9034 14376 9090 14385
rect 9034 14311 9036 14320
rect 9088 14311 9090 14320
rect 9036 14282 9088 14288
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 11626 9076 12038
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 9140 10962 9168 15030
rect 9494 14920 9550 14929
rect 9312 14884 9364 14890
rect 9494 14855 9550 14864
rect 9312 14826 9364 14832
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9232 13530 9260 14486
rect 9324 14385 9352 14826
rect 9404 14816 9456 14822
rect 9402 14784 9404 14793
rect 9456 14784 9458 14793
rect 9402 14719 9458 14728
rect 9508 14482 9536 14855
rect 9600 14550 9628 15370
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9692 14958 9720 15302
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9310 14376 9366 14385
rect 9310 14311 9366 14320
rect 9692 14278 9720 14894
rect 9876 14890 9904 15302
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 9772 14544 9824 14550
rect 9876 14521 9904 14826
rect 9772 14486 9824 14492
rect 9862 14512 9918 14521
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9692 12986 9720 14214
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9218 10976 9274 10985
rect 9140 10934 9218 10962
rect 9218 10911 9274 10920
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10266 9168 10406
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8496 9654 8524 9998
rect 9232 9722 9260 10911
rect 9692 10713 9720 11086
rect 9784 10849 9812 14486
rect 9862 14447 9918 14456
rect 9876 14414 9904 14447
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 12170 9904 14350
rect 9968 14346 9996 20198
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 10322 19952 10378 19961
rect 10322 19887 10378 19896
rect 11612 19916 11664 19922
rect 10336 18970 10364 19887
rect 11612 19858 11664 19864
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 10888 19378 10916 19654
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10138 18864 10194 18873
rect 10704 18834 10732 19110
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 11348 18970 11376 19314
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 10138 18799 10194 18808
rect 10692 18828 10744 18834
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10060 17134 10088 17682
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10152 14550 10180 18799
rect 10692 18770 10744 18776
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10612 18426 10640 18634
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10244 16590 10272 17614
rect 10336 16726 10364 18362
rect 10796 17882 10824 18702
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 11348 17814 11376 18906
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10428 17066 10456 17478
rect 10704 17270 10732 17750
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10980 17202 11008 17546
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10428 16794 10456 17002
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10600 16584 10652 16590
rect 10980 16572 11008 16662
rect 10980 16544 11100 16572
rect 10600 16526 10652 16532
rect 10612 16114 10640 16526
rect 11072 16250 11100 16544
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10336 14822 10364 15506
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9968 12782 9996 13126
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9968 11898 9996 12718
rect 10152 12306 10180 13767
rect 10244 13530 10272 14554
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10244 11898 10272 12174
rect 10336 12102 10364 14758
rect 10612 14414 10640 14758
rect 10888 14482 10916 15438
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10612 14074 10640 14350
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10704 13870 10732 14418
rect 11256 14074 11284 14418
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10704 12442 10732 13806
rect 11348 13802 11376 16934
rect 11440 15609 11468 19654
rect 11624 19174 11652 19858
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11624 18873 11652 19110
rect 11610 18864 11666 18873
rect 11610 18799 11666 18808
rect 11794 18864 11850 18873
rect 11794 18799 11850 18808
rect 11610 16552 11666 16561
rect 11610 16487 11666 16496
rect 11704 16516 11756 16522
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11426 15600 11482 15609
rect 11426 15535 11482 15544
rect 11532 15042 11560 15846
rect 11624 15570 11652 16487
rect 11704 16458 11756 16464
rect 11716 15570 11744 16458
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11624 15162 11652 15506
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11532 15014 11652 15042
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11624 13326 11652 15014
rect 11716 14618 11744 15506
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11072 12986 11100 13126
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10784 12640 10836 12646
rect 10782 12608 10784 12617
rect 10836 12608 10838 12617
rect 10782 12543 10838 12552
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10888 12306 10916 12650
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10138 11520 10194 11529
rect 10138 11455 10194 11464
rect 10152 11354 10180 11455
rect 10520 11354 10548 12242
rect 10782 12200 10838 12209
rect 10600 12164 10652 12170
rect 10782 12135 10838 12144
rect 10600 12106 10652 12112
rect 10612 11830 10640 12106
rect 10796 12102 10824 12135
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 9770 10840 9826 10849
rect 9770 10775 9826 10784
rect 9678 10704 9734 10713
rect 9678 10639 9734 10648
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8574 9616 8630 9625
rect 8574 9551 8630 9560
rect 8588 9382 8616 9551
rect 8772 9450 8800 9658
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8298 9072 8354 9081
rect 8298 9007 8354 9016
rect 8588 8838 8616 9318
rect 8864 9178 8892 9454
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 7852 7954 7880 8774
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 6288 6458 6316 6734
rect 6932 6662 6960 7822
rect 7484 7410 7512 7822
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 7002 7236 7142
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7208 6905 7236 6938
rect 7484 6934 7512 7346
rect 7852 7206 7880 7890
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7472 6928 7524 6934
rect 7194 6896 7250 6905
rect 7472 6870 7524 6876
rect 7194 6831 7250 6840
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5817 5856 6054
rect 5814 5808 5870 5817
rect 5814 5743 5870 5752
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 6932 3097 6960 6598
rect 7484 6458 7512 6870
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7852 4049 7880 7142
rect 8312 6934 8340 7142
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 7838 4040 7894 4049
rect 7838 3975 7894 3984
rect 6918 3088 6974 3097
rect 6918 3023 6974 3032
rect 8312 2650 8340 6870
rect 8588 5273 8616 8774
rect 8574 5264 8630 5273
rect 8574 5199 8630 5208
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7208 2417 7236 2450
rect 7194 2408 7250 2417
rect 7194 2343 7250 2352
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 4066 2136 4122 2145
rect 4066 2071 4122 2080
rect 2686 1456 2742 1465
rect 2686 1391 2742 1400
rect 5000 480 5028 2246
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 10428 1329 10456 10406
rect 10704 9489 10732 12038
rect 10796 10606 10824 12038
rect 11348 11898 11376 12242
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 10888 11354 10916 11834
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 11440 11354 11468 13126
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11532 12850 11560 12922
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12374 11560 12786
rect 11624 12646 11652 13262
rect 11612 12640 11664 12646
rect 11610 12608 11612 12617
rect 11664 12608 11666 12617
rect 11610 12543 11666 12552
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11532 11898 11560 12310
rect 11716 12102 11744 13398
rect 11808 12889 11836 18799
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11992 17882 12020 19654
rect 12176 19553 12204 23520
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12452 19961 12480 20334
rect 13648 19961 13676 22102
rect 14016 20602 14044 23520
rect 15948 23474 15976 23520
rect 15856 23446 15976 23474
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 15580 20466 15608 20742
rect 15856 20602 15884 23446
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 17788 20602 17816 23520
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 19260 20466 19288 20742
rect 19628 20602 19656 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 14924 20392 14976 20398
rect 14554 20360 14610 20369
rect 14924 20334 14976 20340
rect 14554 20295 14556 20304
rect 14608 20295 14610 20304
rect 14556 20266 14608 20272
rect 14936 20262 14964 20334
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 12438 19952 12494 19961
rect 12438 19887 12494 19896
rect 13634 19952 13690 19961
rect 13634 19887 13690 19896
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12162 19544 12218 19553
rect 12162 19479 12218 19488
rect 12544 19378 12572 19790
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12348 19304 12400 19310
rect 12400 19252 12480 19258
rect 12348 19246 12480 19252
rect 12360 19230 12480 19246
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12360 18222 12388 18362
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12452 17882 12480 19230
rect 12544 18970 12572 19314
rect 12820 19310 12848 19654
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12898 19272 12954 19281
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12544 18222 12572 18906
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 11992 17649 12020 17818
rect 12164 17672 12216 17678
rect 11978 17640 12034 17649
rect 12164 17614 12216 17620
rect 11978 17575 12034 17584
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12084 16998 12112 17070
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11992 15366 12020 16050
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11794 12880 11850 12889
rect 11794 12815 11850 12824
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11256 10810 11284 11086
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 11348 10266 11376 11222
rect 11440 10810 11468 11290
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10690 9480 10746 9489
rect 10690 9415 10746 9424
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 11900 7313 11928 15098
rect 11992 15094 12020 15302
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11992 14278 12020 15030
rect 11980 14272 12032 14278
rect 12084 14249 12112 16934
rect 12176 16697 12204 17614
rect 12728 17524 12756 18362
rect 12820 18086 12848 19246
rect 12898 19207 12954 19216
rect 12912 19174 12940 19207
rect 12900 19168 12952 19174
rect 13544 19168 13596 19174
rect 12900 19110 12952 19116
rect 13542 19136 13544 19145
rect 13596 19136 13598 19145
rect 13542 19071 13598 19080
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12808 17536 12860 17542
rect 12728 17496 12808 17524
rect 12808 17478 12860 17484
rect 12820 17270 12848 17478
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12440 16720 12492 16726
rect 12162 16688 12218 16697
rect 12440 16662 12492 16668
rect 12162 16623 12218 16632
rect 12176 16250 12204 16623
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12452 15910 12480 16662
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12162 15600 12218 15609
rect 12162 15535 12218 15544
rect 11980 14214 12032 14220
rect 12070 14240 12126 14249
rect 11992 14074 12020 14214
rect 12070 14175 12126 14184
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12176 13569 12204 15535
rect 12254 15328 12310 15337
rect 12254 15263 12310 15272
rect 12268 13734 12296 15263
rect 12544 14929 12572 16934
rect 12820 16794 12848 17206
rect 12900 16992 12952 16998
rect 12898 16960 12900 16969
rect 12952 16960 12954 16969
rect 12898 16895 12954 16904
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16108 12768 16114
rect 12820 16096 12848 16730
rect 12768 16068 12848 16096
rect 12716 16050 12768 16056
rect 13004 16046 13032 18566
rect 13648 17882 13676 19887
rect 14016 19514 14044 20198
rect 14554 19680 14610 19689
rect 14554 19615 14610 19624
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13924 18154 13952 19110
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17202 13124 17478
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12622 15464 12678 15473
rect 12622 15399 12678 15408
rect 12530 14920 12586 14929
rect 12530 14855 12586 14864
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12452 13841 12480 13942
rect 12438 13832 12494 13841
rect 12438 13767 12494 13776
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12162 13560 12218 13569
rect 12162 13495 12218 13504
rect 12636 12782 12664 15399
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 13530 12756 13806
rect 12806 13560 12862 13569
rect 12716 13524 12768 13530
rect 12806 13495 12862 13504
rect 12716 13466 12768 13472
rect 12820 13190 12848 13495
rect 12808 13184 12860 13190
rect 12912 13161 12940 14758
rect 13096 14482 13124 17138
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 15366 13492 16594
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13174 15192 13230 15201
rect 13174 15127 13176 15136
rect 13228 15127 13230 15136
rect 13176 15098 13228 15104
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13188 14521 13216 14554
rect 13174 14512 13230 14521
rect 13084 14476 13136 14482
rect 13174 14447 13230 14456
rect 13084 14418 13136 14424
rect 13096 13938 13124 14418
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 13190 13032 13670
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12992 13184 13044 13190
rect 12808 13126 12860 13132
rect 12898 13152 12954 13161
rect 12820 12889 12848 13126
rect 12992 13126 13044 13132
rect 12898 13087 12954 13096
rect 12806 12880 12862 12889
rect 12806 12815 12862 12824
rect 12820 12782 12848 12815
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 11286 12480 12582
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12728 11150 12756 12378
rect 13096 12102 13124 13466
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13188 12986 13216 13262
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13280 12442 13308 13874
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12850 13400 13262
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13096 11257 13124 12038
rect 13464 11257 13492 12922
rect 13082 11248 13138 11257
rect 13082 11183 13138 11192
rect 13450 11248 13506 11257
rect 13450 11183 13506 11192
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12254 10976 12310 10985
rect 12254 10911 12310 10920
rect 12268 10810 12296 10911
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 13464 8537 13492 11183
rect 13556 10577 13584 17274
rect 13648 17202 13676 17818
rect 13832 17814 13860 18022
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 14292 17678 14320 18090
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14280 17672 14332 17678
rect 14094 17640 14150 17649
rect 14384 17649 14412 17682
rect 14280 17614 14332 17620
rect 14370 17640 14426 17649
rect 14094 17575 14150 17584
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 14108 16794 14136 17575
rect 14292 16998 14320 17614
rect 14370 17575 14426 17584
rect 14384 17338 14412 17575
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 13832 16590 13860 16730
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13648 15570 13676 16526
rect 13832 15706 13860 16526
rect 14292 16522 14320 16934
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13818 15600 13874 15609
rect 13636 15564 13688 15570
rect 13818 15535 13874 15544
rect 13636 15506 13688 15512
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13648 13462 13676 15302
rect 13728 13524 13780 13530
rect 13832 13512 13860 15535
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13924 14929 13952 14962
rect 13910 14920 13966 14929
rect 13910 14855 13966 14864
rect 13780 13484 13860 13512
rect 13728 13466 13780 13472
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13924 11898 13952 14855
rect 14568 12986 14596 19615
rect 14936 17513 14964 20198
rect 15120 20058 15148 20198
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15212 19258 15240 19858
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 19310 15332 19654
rect 15120 19242 15240 19258
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15108 19236 15240 19242
rect 15160 19230 15240 19236
rect 15108 19178 15160 19184
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 18630 15240 19110
rect 15488 18970 15516 19994
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15028 17746 15056 18158
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 14922 17504 14978 17513
rect 14922 17439 14978 17448
rect 14648 16176 14700 16182
rect 14646 16144 14648 16153
rect 14700 16144 14702 16153
rect 14646 16079 14702 16088
rect 14660 16046 14688 16079
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14936 15745 14964 17439
rect 15028 17338 15056 17682
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15120 17134 15148 17818
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15212 16538 15240 18566
rect 15580 17882 15608 20402
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15856 19174 15884 19790
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 16408 19417 16436 20266
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17512 20058 17540 20198
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16500 19530 16528 19858
rect 17958 19816 18014 19825
rect 17958 19751 18014 19760
rect 16500 19502 16620 19530
rect 16394 19408 16450 19417
rect 16394 19343 16450 19352
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18154 15884 19110
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15304 16697 15332 16730
rect 15290 16688 15346 16697
rect 15290 16623 15346 16632
rect 15212 16510 15332 16538
rect 15014 16416 15070 16425
rect 15014 16351 15070 16360
rect 15028 15910 15056 16351
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 14922 15736 14978 15745
rect 14922 15671 14978 15680
rect 15028 15473 15056 15846
rect 15014 15464 15070 15473
rect 15014 15399 15070 15408
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14844 14822 14872 14962
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14738 14376 14794 14385
rect 14738 14311 14794 14320
rect 14752 14074 14780 14311
rect 14844 14278 14872 14758
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 13530 14964 13670
rect 15120 13530 15148 14758
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14936 13433 14964 13466
rect 14922 13424 14978 13433
rect 14922 13359 14978 13368
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15028 12986 15056 13330
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15028 12442 15056 12718
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15120 12374 15148 13466
rect 15212 12850 15240 15846
rect 15304 13258 15332 16510
rect 15396 15026 15424 17070
rect 15856 16998 15884 18090
rect 16316 17785 16344 18566
rect 16500 18426 16528 19314
rect 16592 19258 16620 19502
rect 16592 19230 16712 19258
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16500 18068 16528 18362
rect 16500 18040 16620 18068
rect 16592 17814 16620 18040
rect 16580 17808 16632 17814
rect 16302 17776 16358 17785
rect 16580 17750 16632 17756
rect 16302 17711 16358 17720
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15568 16448 15620 16454
rect 15672 16425 15700 16594
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15568 16390 15620 16396
rect 15658 16416 15714 16425
rect 15580 16114 15608 16390
rect 15658 16351 15714 16360
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15396 14618 15424 14758
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15396 14074 15424 14554
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15488 13954 15516 15914
rect 15580 15570 15608 16050
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15580 14278 15608 15506
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15396 13926 15516 13954
rect 15580 13938 15608 14214
rect 15568 13932 15620 13938
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12442 15240 12786
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 14844 11121 14872 11494
rect 15304 11393 15332 11494
rect 15290 11384 15346 11393
rect 15290 11319 15346 11328
rect 14830 11112 14886 11121
rect 14830 11047 14886 11056
rect 13542 10568 13598 10577
rect 13542 10503 13598 10512
rect 15396 9625 15424 13926
rect 15568 13874 15620 13880
rect 15476 13864 15528 13870
rect 15474 13832 15476 13841
rect 15528 13832 15530 13841
rect 15474 13767 15530 13776
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15488 12306 15516 13398
rect 15566 12608 15622 12617
rect 15566 12543 15622 12552
rect 15580 12442 15608 12543
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15488 11898 15516 12242
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15488 11354 15516 11698
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15672 10962 15700 15982
rect 15764 15706 15792 16526
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15764 12850 15792 14962
rect 15856 13326 15884 16934
rect 16316 16794 16344 17614
rect 16408 16998 16436 17614
rect 16592 17338 16620 17750
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16684 16658 16712 19230
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 16868 18068 16896 18838
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16960 18426 16988 18702
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17144 18086 17172 18770
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 16948 18080 17000 18086
rect 16868 18040 16948 18068
rect 16948 18022 17000 18028
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 16394 16280 16450 16289
rect 16394 16215 16396 16224
rect 16448 16215 16450 16224
rect 16396 16186 16448 16192
rect 16408 15978 16436 16186
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16304 15360 16356 15366
rect 16580 15360 16632 15366
rect 16304 15302 16356 15308
rect 16500 15308 16580 15314
rect 16500 15302 16632 15308
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16212 14816 16264 14822
rect 16316 14804 16344 15302
rect 16500 15286 16620 15302
rect 16500 15026 16528 15286
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16264 14776 16344 14804
rect 16212 14758 16264 14764
rect 16224 14482 16252 14758
rect 16394 14648 16450 14657
rect 16394 14583 16450 14592
rect 16408 14550 16436 14583
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16486 14512 16542 14521
rect 16212 14476 16264 14482
rect 16264 14436 16344 14464
rect 16212 14418 16264 14424
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16316 13870 16344 14436
rect 16408 14074 16436 14486
rect 16486 14447 16542 14456
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16500 13977 16528 14447
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16486 13968 16542 13977
rect 16486 13903 16542 13912
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16500 13682 16528 13903
rect 16408 13654 16528 13682
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 12986 15884 13262
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 15580 10934 15700 10962
rect 15382 9616 15438 9625
rect 15382 9551 15438 9560
rect 13450 8528 13506 8537
rect 13450 8463 13506 8472
rect 11886 7304 11942 7313
rect 11886 7239 11942 7248
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 15580 5273 15608 10934
rect 15764 10577 15792 12106
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11694 15884 12038
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 16316 11830 16344 12378
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15856 11354 15884 11630
rect 16408 11354 16436 13654
rect 16486 13152 16542 13161
rect 16486 13087 16542 13096
rect 16500 12782 16528 13087
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16500 11626 16528 12582
rect 16684 12424 16712 14010
rect 16960 13190 16988 18022
rect 17144 17649 17172 18022
rect 17788 17882 17816 18362
rect 17880 18086 17908 18702
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17972 17882 18000 19751
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17130 17640 17186 17649
rect 17130 17575 17186 17584
rect 17144 16561 17172 17575
rect 17314 17096 17370 17105
rect 17314 17031 17370 17040
rect 17328 16794 17356 17031
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17130 16552 17186 16561
rect 17130 16487 17186 16496
rect 17236 16250 17264 16730
rect 17328 16425 17356 16730
rect 17788 16640 17816 17818
rect 17958 17776 18014 17785
rect 17958 17711 18014 17720
rect 17972 16794 18000 17711
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17696 16612 17816 16640
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17498 16552 17554 16561
rect 17314 16416 17370 16425
rect 17314 16351 17370 16360
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17328 16182 17356 16351
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 17144 13818 17172 15914
rect 17420 15366 17448 16526
rect 17498 16487 17554 16496
rect 17512 16289 17540 16487
rect 17498 16280 17554 16289
rect 17498 16215 17554 16224
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17052 13802 17172 13818
rect 17040 13796 17172 13802
rect 17092 13790 17172 13796
rect 17040 13738 17092 13744
rect 17144 13410 17172 13790
rect 17512 13462 17540 14214
rect 17696 14074 17724 16612
rect 18064 16538 18092 20334
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18156 19242 18184 19858
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18248 19378 18276 19790
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18156 18426 18184 19178
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 18248 17882 18276 19314
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18156 17377 18184 17818
rect 18142 17368 18198 17377
rect 18142 17303 18198 17312
rect 18156 16658 18184 17303
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 17788 16510 18092 16538
rect 17788 14634 17816 16510
rect 18156 16250 18184 16594
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 18234 15464 18290 15473
rect 17868 14816 17920 14822
rect 17972 14804 18000 15438
rect 18234 15399 18290 15408
rect 17920 14776 18000 14804
rect 17868 14758 17920 14764
rect 17788 14606 17908 14634
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17052 13394 17172 13410
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17040 13388 17172 13394
rect 17092 13382 17172 13388
rect 17040 13330 17092 13336
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 17144 12986 17172 13382
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16592 12396 16712 12424
rect 16592 11778 16620 12396
rect 17052 12306 17080 12786
rect 17144 12306 17172 12922
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16592 11762 16712 11778
rect 16580 11756 16712 11762
rect 16632 11750 16712 11756
rect 16580 11698 16632 11704
rect 16592 11667 16620 11698
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15856 10810 15884 11154
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16408 10810 16436 11290
rect 16592 10810 16620 11494
rect 16684 11150 16712 11750
rect 16960 11354 16988 12174
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 15750 10568 15806 10577
rect 15750 10503 15806 10512
rect 16868 10470 16896 10950
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 16868 9518 16896 10406
rect 17038 10024 17094 10033
rect 17038 9959 17094 9968
rect 17052 9586 17080 9959
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 17328 5817 17356 13126
rect 17512 12986 17540 13398
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17512 11762 17540 12922
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17512 11558 17540 11698
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10169 17448 11154
rect 17406 10160 17462 10169
rect 17406 10095 17462 10104
rect 17512 9654 17540 11494
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17696 9466 17724 13670
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17788 12442 17816 12650
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17880 11354 17908 14606
rect 17972 12986 18000 14776
rect 18248 14074 18276 15399
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 11830 18000 12242
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 11098 18000 11154
rect 17880 11070 18000 11098
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17880 10810 17908 11070
rect 18064 10810 18092 11086
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 18064 10266 18092 10746
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18156 9654 18184 11562
rect 18340 11234 18368 19654
rect 18616 19242 18644 19790
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18616 18630 18644 19178
rect 18984 19174 19012 19246
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18432 15706 18460 17614
rect 18524 17270 18552 17682
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18524 16794 18552 17206
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18512 16448 18564 16454
rect 18616 16436 18644 18566
rect 18984 18086 19012 19110
rect 19168 18970 19196 20198
rect 19536 19961 19564 20198
rect 19522 19952 19578 19961
rect 19522 19887 19578 19896
rect 19628 19825 19656 20198
rect 19614 19816 19670 19825
rect 19614 19751 19670 19760
rect 19628 19718 19656 19751
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19720 19242 19748 20402
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20732 19700 20760 20334
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 20640 19672 20760 19700
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 20260 19236 20312 19242
rect 20260 19178 20312 19184
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19168 18290 19196 18906
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19444 18290 19472 18770
rect 20272 18630 20300 19178
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20534 19136 20590 19145
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18290 20300 18566
rect 20456 18426 20484 19110
rect 20534 19071 20590 19080
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20548 18329 20576 19071
rect 20534 18320 20590 18329
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 20260 18284 20312 18290
rect 20534 18255 20590 18264
rect 20260 18226 20312 18232
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18800 17134 18828 17750
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18984 16998 19012 18022
rect 19444 17678 19472 18226
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17882 20208 18022
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 18564 16408 18644 16436
rect 18512 16390 18564 16396
rect 18524 16046 18552 16390
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18602 16008 18658 16017
rect 18984 15978 19012 16934
rect 19076 16590 19104 16934
rect 19444 16794 19472 17614
rect 20272 16998 20300 18226
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20364 17882 20392 18158
rect 20548 18154 20576 18255
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20534 17776 20590 17785
rect 20534 17711 20590 17720
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20456 17338 20484 17546
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18602 15943 18658 15952
rect 18972 15972 19024 15978
rect 18510 15736 18566 15745
rect 18420 15700 18472 15706
rect 18510 15671 18566 15680
rect 18420 15642 18472 15648
rect 18524 15473 18552 15671
rect 18510 15464 18566 15473
rect 18510 15399 18566 15408
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18432 15162 18460 15302
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18510 15056 18566 15065
rect 18510 14991 18566 15000
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18432 12374 18460 13126
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18432 11898 18460 12310
rect 18524 12073 18552 14991
rect 18616 14249 18644 15943
rect 18972 15914 19024 15920
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18800 14618 18828 15506
rect 18984 15042 19012 15914
rect 19076 15502 19104 16526
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19062 15056 19118 15065
rect 18984 15014 19062 15042
rect 19062 14991 19064 15000
rect 19116 14991 19118 15000
rect 19064 14962 19116 14968
rect 19352 14890 19380 15846
rect 19614 14920 19670 14929
rect 19340 14884 19392 14890
rect 19614 14855 19670 14864
rect 20352 14884 20404 14890
rect 19340 14826 19392 14832
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18696 14272 18748 14278
rect 18602 14240 18658 14249
rect 18696 14214 18748 14220
rect 18602 14175 18658 14184
rect 18510 12064 18566 12073
rect 18510 11999 18566 12008
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18248 11206 18368 11234
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 17696 9438 18000 9466
rect 17972 9382 18000 9438
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 9110 18000 9318
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18248 6225 18276 11206
rect 18432 11150 18460 11834
rect 18420 11144 18472 11150
rect 18326 11112 18382 11121
rect 18420 11086 18472 11092
rect 18326 11047 18382 11056
rect 18340 10266 18368 11047
rect 18432 10742 18460 11086
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18340 9178 18368 10066
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18524 9722 18552 9998
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18418 9616 18474 9625
rect 18418 9551 18420 9560
rect 18472 9551 18474 9560
rect 18420 9522 18472 9528
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18616 9042 18644 14175
rect 18708 13734 18736 14214
rect 18800 14074 18828 14554
rect 19352 14346 19380 14826
rect 19628 14482 19656 14855
rect 20352 14826 20404 14832
rect 20364 14618 20392 14826
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14657 20484 14758
rect 20442 14648 20498 14657
rect 20352 14612 20404 14618
rect 20442 14583 20498 14592
rect 20352 14554 20404 14560
rect 19708 14544 19760 14550
rect 19708 14486 19760 14492
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 14113 19288 14214
rect 19246 14104 19302 14113
rect 18788 14068 18840 14074
rect 19628 14074 19656 14418
rect 19246 14039 19302 14048
rect 19616 14068 19668 14074
rect 18788 14010 18840 14016
rect 19616 14010 19668 14016
rect 18880 14000 18932 14006
rect 18800 13948 18880 13954
rect 18800 13942 18932 13948
rect 18800 13926 18920 13942
rect 19156 13932 19208 13938
rect 18800 13870 18828 13926
rect 19156 13874 19208 13880
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 18708 12753 18736 12951
rect 18694 12744 18750 12753
rect 18694 12679 18750 12688
rect 18800 11257 18828 13806
rect 18878 13560 18934 13569
rect 18878 13495 18934 13504
rect 18892 13297 18920 13495
rect 18878 13288 18934 13297
rect 18878 13223 18934 13232
rect 18786 11248 18842 11257
rect 18786 11183 18842 11192
rect 18892 9178 18920 13223
rect 19168 12850 19196 13874
rect 19616 13864 19668 13870
rect 19614 13832 19616 13841
rect 19668 13832 19670 13841
rect 19614 13767 19670 13776
rect 19248 13728 19300 13734
rect 19300 13688 19380 13716
rect 19248 13670 19300 13676
rect 19352 12889 19380 13688
rect 19720 13462 19748 14486
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19708 13456 19760 13462
rect 19708 13398 19760 13404
rect 19338 12880 19394 12889
rect 19156 12844 19208 12850
rect 19338 12815 19394 12824
rect 19156 12786 19208 12792
rect 19062 12744 19118 12753
rect 19062 12679 19064 12688
rect 19116 12679 19118 12688
rect 19064 12650 19116 12656
rect 19352 12209 19380 12815
rect 19338 12200 19394 12209
rect 19394 12158 19472 12186
rect 19338 12135 19394 12144
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11626 19196 12038
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19168 11286 19196 11562
rect 19246 11520 19302 11529
rect 19246 11455 19302 11464
rect 19260 11354 19288 11455
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19352 11098 19380 11290
rect 19444 11286 19472 12158
rect 19614 12064 19670 12073
rect 19614 11999 19670 12008
rect 19628 11354 19656 11999
rect 19706 11384 19762 11393
rect 19616 11348 19668 11354
rect 19706 11319 19762 11328
rect 19616 11290 19668 11296
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19260 11070 19380 11098
rect 19260 10810 19288 11070
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19444 10266 19472 11222
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19168 9722 19196 10202
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19720 9654 19748 11319
rect 19812 10266 19840 14214
rect 19904 13841 19932 14350
rect 20364 13938 20392 14554
rect 20548 14550 20576 17711
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20260 13864 20312 13870
rect 19890 13832 19946 13841
rect 20260 13806 20312 13812
rect 19890 13767 19946 13776
rect 19904 13530 19932 13767
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19890 11248 19946 11257
rect 19890 11183 19946 11192
rect 19904 10538 19932 11183
rect 20180 11150 20208 11494
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20180 10674 20208 11086
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 19984 10600 20036 10606
rect 19982 10568 19984 10577
rect 20036 10568 20038 10577
rect 19892 10532 19944 10538
rect 19982 10503 20038 10512
rect 19892 10474 19944 10480
rect 19996 10266 20024 10503
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19812 9586 19840 10202
rect 20272 9704 20300 13806
rect 20444 13796 20496 13802
rect 20444 13738 20496 13744
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20364 13433 20392 13466
rect 20350 13424 20406 13433
rect 20350 13359 20406 13368
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20364 10849 20392 13262
rect 20456 12850 20484 13738
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20548 13530 20576 13670
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20548 12730 20576 13466
rect 20640 12986 20668 19672
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20916 18222 20944 18702
rect 20904 18216 20956 18222
rect 20810 18184 20866 18193
rect 20904 18158 20956 18164
rect 20810 18119 20812 18128
rect 20864 18119 20866 18128
rect 20812 18090 20864 18096
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 21284 17105 21312 20742
rect 21560 20602 21588 23520
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21362 19952 21418 19961
rect 21362 19887 21418 19896
rect 21376 18306 21404 19887
rect 23400 19553 23428 23520
rect 24950 21584 25006 21593
rect 24950 21519 25006 21528
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23860 20262 23888 20946
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 22006 19544 22062 19553
rect 22006 19479 22062 19488
rect 23386 19544 23442 19553
rect 23386 19479 23442 19488
rect 21824 19304 21876 19310
rect 21454 19272 21510 19281
rect 21824 19246 21876 19252
rect 21454 19207 21510 19216
rect 21468 18970 21496 19207
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21468 18426 21496 18906
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21376 18278 21496 18306
rect 21560 18290 21588 18566
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21376 17338 21404 17682
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21270 17096 21326 17105
rect 21270 17031 21326 17040
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16250 21220 16390
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20456 12702 20576 12730
rect 20350 10840 20406 10849
rect 20350 10775 20406 10784
rect 20180 9676 20300 9704
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18616 8634 18644 8978
rect 18892 8634 18920 9114
rect 19260 8974 19288 9522
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20088 9178 20116 9454
rect 20180 9382 20208 9676
rect 20352 9648 20404 9654
rect 20456 9636 20484 12702
rect 20732 12646 20760 13126
rect 20824 12986 20852 13942
rect 21100 13802 21128 14418
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 21284 13716 21312 17031
rect 21376 16182 21404 17274
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 21376 15706 21404 16118
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21468 15450 21496 18278
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21560 17542 21588 18226
rect 21638 17776 21694 17785
rect 21638 17711 21694 17720
rect 21548 17536 21600 17542
rect 21652 17513 21680 17711
rect 21548 17478 21600 17484
rect 21638 17504 21694 17513
rect 21560 16590 21588 17478
rect 21638 17439 21694 17448
rect 21836 17338 21864 19246
rect 22020 19174 22048 19479
rect 22466 19408 22522 19417
rect 22466 19343 22522 19352
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22480 18970 22508 19343
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 23110 18864 23166 18873
rect 22008 18828 22060 18834
rect 23110 18799 23166 18808
rect 22008 18770 22060 18776
rect 22020 18222 22048 18770
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 21916 18080 21968 18086
rect 22100 18080 22152 18086
rect 21916 18022 21968 18028
rect 22020 18040 22100 18068
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21560 15910 21588 16526
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21560 15638 21588 15846
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21468 15422 21588 15450
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21468 15094 21496 15302
rect 21456 15088 21508 15094
rect 21454 15056 21456 15065
rect 21508 15056 21510 15065
rect 21454 14991 21510 15000
rect 21468 14414 21496 14991
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 14074 21404 14214
rect 21468 14074 21496 14350
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21284 13688 21404 13716
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 21008 12850 21036 13126
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20548 11898 20576 12038
rect 20824 11898 20852 12718
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20916 11830 20944 12242
rect 21192 11830 21220 12242
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 20720 11688 20772 11694
rect 20640 11636 20720 11642
rect 20640 11630 20772 11636
rect 20640 11614 20760 11630
rect 20812 11620 20864 11626
rect 20640 10810 20668 11614
rect 20812 11562 20864 11568
rect 20824 11529 20852 11562
rect 20810 11520 20866 11529
rect 20810 11455 20866 11464
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 21180 11212 21232 11218
rect 21180 11154 21232 11160
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 21192 10742 21220 11154
rect 21284 10810 21312 12582
rect 21376 11778 21404 13688
rect 21468 13462 21496 14010
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21468 12374 21496 13398
rect 21456 12368 21508 12374
rect 21560 12345 21588 15422
rect 21652 15162 21680 17002
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21836 16250 21864 16730
rect 21928 16708 21956 18022
rect 22020 17882 22048 18040
rect 22100 18022 22152 18028
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22296 17270 22324 17478
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 16794 22232 16934
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22008 16720 22060 16726
rect 21928 16680 22008 16708
rect 22008 16662 22060 16668
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21822 16144 21878 16153
rect 21822 16079 21878 16088
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 15502 21772 15846
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21744 14074 21772 14894
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 21456 12310 21508 12316
rect 21546 12336 21602 12345
rect 21546 12271 21602 12280
rect 21376 11750 21496 11778
rect 21362 11656 21418 11665
rect 21362 11591 21418 11600
rect 21376 11354 21404 11591
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21180 10736 21232 10742
rect 21180 10678 21232 10684
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20404 9608 20484 9636
rect 20352 9590 20404 9596
rect 20824 9586 20852 10406
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 21376 10266 21404 10610
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21468 10198 21496 11750
rect 21560 11218 21588 12271
rect 21652 11558 21680 12650
rect 21744 12481 21772 13466
rect 21836 13025 21864 16079
rect 21928 15910 21956 16390
rect 22112 15910 22140 16662
rect 22296 16454 22324 17206
rect 22388 16454 22416 17682
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22388 16114 22416 16390
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22020 14958 22048 15506
rect 22388 15026 22416 16050
rect 22480 16046 22508 18634
rect 23124 18426 23152 18799
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23124 18222 23152 18362
rect 23492 18290 23520 18566
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 22652 18148 22704 18154
rect 22652 18090 22704 18096
rect 22744 18148 22796 18154
rect 22744 18090 22796 18096
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22572 14822 22600 15506
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22572 14278 22600 14758
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13530 22140 13670
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21822 13016 21878 13025
rect 21822 12951 21878 12960
rect 21730 12472 21786 12481
rect 21730 12407 21786 12416
rect 21836 11914 21864 12951
rect 21928 12442 21956 13330
rect 22112 12986 22140 13466
rect 22190 13424 22246 13433
rect 22190 13359 22246 13368
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22204 12782 22232 13359
rect 22572 12850 22600 14214
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22204 12646 22232 12718
rect 22192 12640 22244 12646
rect 22468 12640 22520 12646
rect 22192 12582 22244 12588
rect 22466 12608 22468 12617
rect 22520 12608 22522 12617
rect 22466 12543 22522 12552
rect 22572 12442 22600 12786
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 21744 11886 21864 11914
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21640 10532 21692 10538
rect 21640 10474 21692 10480
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 21560 9722 21588 10406
rect 21652 9994 21680 10474
rect 21744 10282 21772 11886
rect 21928 11778 21956 12378
rect 21836 11762 21956 11778
rect 21824 11756 21956 11762
rect 21876 11750 21956 11756
rect 21824 11698 21876 11704
rect 21836 11014 21864 11698
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 22112 11354 22140 11562
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 21824 11008 21876 11014
rect 21824 10950 21876 10956
rect 21836 10674 21864 10950
rect 22006 10840 22062 10849
rect 22006 10775 22062 10784
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21744 10254 21864 10282
rect 22020 10266 22048 10775
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 21454 9480 21510 9489
rect 21454 9415 21456 9424
rect 21508 9415 21510 9424
rect 21456 9386 21508 9392
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19248 8968 19300 8974
rect 20180 8945 20208 9318
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 21744 9178 21772 10134
rect 21836 9518 21864 10254
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22020 10010 22048 10202
rect 22284 10056 22336 10062
rect 22020 9982 22140 10010
rect 22284 9998 22336 10004
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 22112 9178 22140 9982
rect 22296 9586 22324 9998
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 19248 8910 19300 8916
rect 20166 8936 20222 8945
rect 19260 8634 19288 8910
rect 20166 8871 20222 8880
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 22664 7993 22692 18090
rect 22756 13870 22784 18090
rect 23110 17776 23166 17785
rect 23110 17711 23166 17720
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22848 14074 22876 15574
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 23020 13456 23072 13462
rect 23020 13398 23072 13404
rect 23032 12986 23060 13398
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23124 11898 23152 17711
rect 23768 16454 23796 19110
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23768 16046 23796 16390
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23754 15464 23810 15473
rect 23754 15399 23810 15408
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23492 14822 23520 14962
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23492 13161 23520 14758
rect 23664 14544 23716 14550
rect 23662 14512 23664 14521
rect 23716 14512 23718 14521
rect 23662 14447 23718 14456
rect 23676 14074 23704 14447
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23768 13818 23796 15399
rect 23584 13790 23796 13818
rect 23478 13152 23534 13161
rect 23478 13087 23534 13096
rect 23584 12306 23612 13790
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23768 12918 23796 13262
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23664 12708 23716 12714
rect 23664 12650 23716 12656
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23584 11898 23612 12242
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 22756 11354 22784 11494
rect 23676 11354 23704 12650
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 22756 10266 22784 11290
rect 23480 11280 23532 11286
rect 23400 11228 23480 11234
rect 23400 11222 23532 11228
rect 23400 11206 23520 11222
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22940 10470 22968 11086
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 23308 9466 23336 11018
rect 23400 10810 23428 11206
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23676 10674 23704 11290
rect 23768 11121 23796 12038
rect 23754 11112 23810 11121
rect 23754 11047 23810 11056
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23400 10266 23428 10474
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23676 10198 23704 10610
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23664 10192 23716 10198
rect 23664 10134 23716 10140
rect 23768 10130 23796 10406
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 23400 9654 23428 10066
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23308 9450 23520 9466
rect 23308 9444 23532 9450
rect 23308 9438 23480 9444
rect 23480 9386 23532 9392
rect 23768 8974 23796 10066
rect 23860 9654 23888 20198
rect 24136 19514 24164 20198
rect 24400 19916 24452 19922
rect 24400 19858 24452 19864
rect 24124 19508 24176 19514
rect 24124 19450 24176 19456
rect 24216 19304 24268 19310
rect 24216 19246 24268 19252
rect 24228 18902 24256 19246
rect 24216 18896 24268 18902
rect 24216 18838 24268 18844
rect 24412 18329 24440 19858
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24780 19394 24808 19654
rect 24780 19366 24900 19394
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24398 18320 24454 18329
rect 24398 18255 24454 18264
rect 23940 18080 23992 18086
rect 23938 18048 23940 18057
rect 24032 18080 24084 18086
rect 23992 18048 23994 18057
rect 24032 18022 24084 18028
rect 23938 17983 23994 17992
rect 24044 17542 24072 18022
rect 24124 17604 24176 17610
rect 24124 17546 24176 17552
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 24044 14498 24072 17478
rect 24136 17066 24164 17546
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24136 16794 24164 17002
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24136 15026 24164 15302
rect 24228 15026 24256 15574
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24136 14618 24164 14962
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24044 14470 24164 14498
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 24044 14249 24072 14350
rect 24030 14240 24086 14249
rect 24030 14175 24086 14184
rect 24044 14074 24072 14175
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23938 13832 23994 13841
rect 23938 13767 23940 13776
rect 23992 13767 23994 13776
rect 23940 13738 23992 13744
rect 23952 13530 23980 13738
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 24044 12918 24072 14010
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 24136 12481 24164 14470
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24320 13870 24348 14214
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24320 13462 24348 13806
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 24306 13152 24362 13161
rect 24306 13087 24362 13096
rect 24122 12472 24178 12481
rect 24122 12407 24178 12416
rect 24122 12336 24178 12345
rect 24122 12271 24124 12280
rect 24176 12271 24178 12280
rect 24124 12242 24176 12248
rect 24136 11694 24164 12242
rect 24320 12186 24348 13087
rect 24228 12158 24348 12186
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 24228 9738 24256 12158
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24320 11830 24348 12038
rect 24308 11824 24360 11830
rect 24308 11766 24360 11772
rect 24320 11150 24348 11766
rect 24412 11354 24440 18255
rect 24688 18086 24716 18770
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24688 17338 24716 18022
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24780 16232 24808 18226
rect 24872 16794 24900 19366
rect 24964 18873 24992 21519
rect 25056 19922 25084 23559
rect 25226 23520 25282 24000
rect 27158 23520 27214 24000
rect 28998 23520 29054 24000
rect 25240 20602 25268 23520
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25134 20496 25190 20505
rect 25134 20431 25190 20440
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 25056 19378 25084 19722
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 24950 18864 25006 18873
rect 24950 18799 25006 18808
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24964 16425 24992 18294
rect 25042 17232 25098 17241
rect 25042 17167 25098 17176
rect 24950 16416 25006 16425
rect 24950 16351 25006 16360
rect 24860 16244 24912 16250
rect 24780 16204 24860 16232
rect 24860 16186 24912 16192
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24596 14822 24624 15506
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24596 11626 24624 14758
rect 24872 14618 24900 16186
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24674 14376 24730 14385
rect 24674 14311 24730 14320
rect 24688 12442 24716 14311
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24964 12345 24992 15914
rect 25056 15094 25084 17167
rect 25148 16538 25176 20431
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25240 19922 25268 20198
rect 25424 19938 25452 23015
rect 25686 22400 25742 22409
rect 25686 22335 25742 22344
rect 25502 21312 25558 21321
rect 25502 21247 25558 21256
rect 25516 20806 25544 21247
rect 25504 20800 25556 20806
rect 25504 20742 25556 20748
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25516 19990 25544 20198
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25332 19910 25452 19938
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 25240 19009 25268 19858
rect 25332 19292 25360 19910
rect 25412 19848 25464 19854
rect 25412 19790 25464 19796
rect 25424 19514 25452 19790
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25516 19446 25544 19926
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25332 19264 25452 19292
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25226 19000 25282 19009
rect 25332 18970 25360 19110
rect 25226 18935 25282 18944
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25226 18864 25282 18873
rect 25226 18799 25282 18808
rect 25240 17785 25268 18799
rect 25424 18358 25452 19264
rect 25700 19174 25728 22335
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 27172 21146 27200 23520
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 29012 21078 29040 23520
rect 29000 21072 29052 21078
rect 29000 21014 29052 21020
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 25792 20330 25820 20742
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 18465 25728 19110
rect 25792 18970 25820 20266
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25884 19718 25912 20198
rect 26160 19854 26188 20402
rect 26148 19848 26200 19854
rect 26516 19848 26568 19854
rect 26200 19796 26372 19802
rect 26148 19790 26372 19796
rect 26516 19790 26568 19796
rect 26160 19774 26372 19790
rect 26160 19725 26188 19774
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25884 19514 25912 19654
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25872 19508 25924 19514
rect 25872 19450 25924 19456
rect 26344 19258 26372 19774
rect 26528 19310 26556 19790
rect 26516 19304 26568 19310
rect 26344 19230 26464 19258
rect 26516 19246 26568 19252
rect 25780 18964 25832 18970
rect 25780 18906 25832 18912
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25686 18456 25742 18465
rect 25956 18448 26252 18468
rect 26436 18426 26464 19230
rect 26514 19000 26570 19009
rect 26514 18935 26570 18944
rect 25686 18391 25742 18400
rect 26424 18420 26476 18426
rect 26424 18362 26476 18368
rect 25412 18352 25464 18358
rect 25412 18294 25464 18300
rect 25412 18148 25464 18154
rect 25412 18090 25464 18096
rect 25226 17776 25282 17785
rect 25226 17711 25282 17720
rect 25424 17542 25452 18090
rect 25688 17808 25740 17814
rect 25688 17750 25740 17756
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25240 16726 25268 17478
rect 25318 17368 25374 17377
rect 25318 17303 25320 17312
rect 25372 17303 25374 17312
rect 25320 17274 25372 17280
rect 25424 17202 25452 17478
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 25424 16590 25452 17138
rect 25516 16998 25544 17614
rect 25596 17604 25648 17610
rect 25596 17546 25648 17552
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25516 16794 25544 16934
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25320 16584 25372 16590
rect 25148 16510 25268 16538
rect 25320 16526 25372 16532
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 25134 15872 25190 15881
rect 25134 15807 25190 15816
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 25042 14648 25098 14657
rect 25042 14583 25098 14592
rect 24766 12336 24822 12345
rect 24766 12271 24822 12280
rect 24950 12336 25006 12345
rect 24950 12271 25006 12280
rect 24780 12073 24808 12271
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24766 12064 24822 12073
rect 24766 11999 24822 12008
rect 24584 11620 24636 11626
rect 24584 11562 24636 11568
rect 24964 11354 24992 12174
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24308 11144 24360 11150
rect 24308 11086 24360 11092
rect 24320 10538 24348 11086
rect 24412 10810 24440 11290
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 24228 9710 24348 9738
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 24216 9444 24268 9450
rect 24216 9386 24268 9392
rect 24228 9110 24256 9386
rect 24216 9104 24268 9110
rect 24216 9046 24268 9052
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 22650 7984 22706 7993
rect 22650 7919 22706 7928
rect 24320 7449 24348 9710
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24504 9178 24532 9318
rect 24872 9178 24900 10678
rect 25056 10033 25084 14583
rect 25148 14550 25176 15807
rect 25136 14544 25188 14550
rect 25136 14486 25188 14492
rect 25134 14104 25190 14113
rect 25134 14039 25190 14048
rect 25148 12238 25176 14039
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25134 10432 25190 10441
rect 25134 10367 25190 10376
rect 25042 10024 25098 10033
rect 25042 9959 25098 9968
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9586 24992 9862
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24872 8106 24900 9114
rect 24780 8090 24900 8106
rect 24768 8084 24900 8090
rect 24820 8078 24900 8084
rect 24768 8026 24820 8032
rect 24306 7440 24362 7449
rect 24306 7375 24362 7384
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 18234 6216 18290 6225
rect 18234 6151 18290 6160
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 17314 5808 17370 5817
rect 17314 5743 17370 5752
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 15566 5264 15622 5273
rect 15566 5199 15622 5208
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 14922 2408 14978 2417
rect 14922 2343 14978 2352
rect 10414 1320 10470 1329
rect 10414 1255 10470 1264
rect 14936 480 14964 2343
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 24964 480 24992 9522
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25056 8634 25084 9114
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 25148 8566 25176 10367
rect 25240 9625 25268 16510
rect 25332 15706 25360 16526
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25424 15638 25452 16526
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25516 16182 25544 16458
rect 25504 16176 25556 16182
rect 25502 16144 25504 16153
rect 25556 16144 25558 16153
rect 25502 16079 25558 16088
rect 25412 15632 25464 15638
rect 25412 15574 25464 15580
rect 25504 15496 25556 15502
rect 25318 15464 25374 15473
rect 25504 15438 25556 15444
rect 25318 15399 25374 15408
rect 25412 15428 25464 15434
rect 25332 15162 25360 15399
rect 25412 15370 25464 15376
rect 25320 15156 25372 15162
rect 25320 15098 25372 15104
rect 25424 14890 25452 15370
rect 25412 14884 25464 14890
rect 25412 14826 25464 14832
rect 25424 14362 25452 14826
rect 25516 14550 25544 15438
rect 25504 14544 25556 14550
rect 25504 14486 25556 14492
rect 25424 14334 25544 14362
rect 25412 13524 25464 13530
rect 25412 13466 25464 13472
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25226 9616 25282 9625
rect 25332 9602 25360 12922
rect 25424 12782 25452 13466
rect 25412 12776 25464 12782
rect 25516 12753 25544 14334
rect 25412 12718 25464 12724
rect 25502 12744 25558 12753
rect 25424 12442 25452 12718
rect 25502 12679 25558 12688
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25516 12238 25544 12679
rect 25608 12374 25636 17546
rect 25700 13977 25728 17750
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 25792 16658 25820 17682
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 26344 17134 26372 17478
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26344 16794 26372 17070
rect 26436 16998 26464 17682
rect 26528 17338 26556 18935
rect 26516 17332 26568 17338
rect 26516 17274 26568 17280
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25686 13968 25742 13977
rect 25686 13903 25742 13912
rect 25688 12708 25740 12714
rect 25688 12650 25740 12656
rect 25596 12368 25648 12374
rect 25596 12310 25648 12316
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25410 12064 25466 12073
rect 25410 11999 25466 12008
rect 25424 9738 25452 11999
rect 25516 11830 25544 12174
rect 25504 11824 25556 11830
rect 25504 11766 25556 11772
rect 25608 11354 25636 12310
rect 25700 11762 25728 12650
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25700 11354 25728 11698
rect 25792 11393 25820 16594
rect 25872 16516 25924 16522
rect 25872 16458 25924 16464
rect 25884 15978 25912 16458
rect 26252 16436 26280 16730
rect 26436 16697 26464 16934
rect 26422 16688 26478 16697
rect 26478 16646 26556 16674
rect 26422 16623 26478 16632
rect 26332 16448 26384 16454
rect 26252 16408 26332 16436
rect 26332 16390 26384 16396
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 26160 15348 26188 15982
rect 26344 15978 26372 16390
rect 26332 15972 26384 15978
rect 26332 15914 26384 15920
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26252 15473 26280 15506
rect 26344 15502 26372 15914
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26332 15496 26384 15502
rect 26238 15464 26294 15473
rect 26332 15438 26384 15444
rect 26238 15399 26294 15408
rect 26332 15360 26384 15366
rect 26160 15320 26332 15348
rect 26332 15302 26384 15308
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 26344 15144 26372 15302
rect 26436 15162 26464 15574
rect 26252 15116 26372 15144
rect 26424 15156 26476 15162
rect 26148 14952 26200 14958
rect 26252 14940 26280 15116
rect 26424 15098 26476 15104
rect 26200 14912 26280 14940
rect 26148 14894 26200 14900
rect 26160 14414 26188 14894
rect 26332 14884 26384 14890
rect 26332 14826 26384 14832
rect 26344 14618 26372 14826
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 25884 13530 25912 14010
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 25976 13326 26004 13670
rect 25964 13320 26016 13326
rect 25884 13280 25964 13308
rect 25884 12306 25912 13280
rect 25964 13262 26016 13268
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26528 13002 26556 16646
rect 26620 14618 26648 20742
rect 26974 20088 27030 20097
rect 26974 20023 27030 20032
rect 26988 19825 27016 20023
rect 26974 19816 27030 19825
rect 26974 19751 27030 19760
rect 26988 18970 27016 19751
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27356 19174 27384 19314
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 26976 18964 27028 18970
rect 26976 18906 27028 18912
rect 26700 18828 26752 18834
rect 26700 18770 26752 18776
rect 26712 18154 26740 18770
rect 26988 18426 27016 18906
rect 27356 18766 27384 19110
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 28172 18760 28224 18766
rect 28172 18702 28224 18708
rect 26976 18420 27028 18426
rect 26976 18362 27028 18368
rect 26974 18320 27030 18329
rect 26974 18255 27030 18264
rect 26700 18148 26752 18154
rect 26700 18090 26752 18096
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26608 14408 26660 14414
rect 26606 14376 26608 14385
rect 26660 14376 26662 14385
rect 26606 14311 26662 14320
rect 26620 14006 26648 14311
rect 26608 14000 26660 14006
rect 26608 13942 26660 13948
rect 26344 12974 26556 13002
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 25884 11898 25912 12242
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 25872 11892 25924 11898
rect 25872 11834 25924 11840
rect 25778 11384 25834 11393
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25688 11348 25740 11354
rect 25778 11319 25834 11328
rect 25688 11290 25740 11296
rect 26344 11234 26372 12974
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26436 12170 26464 12582
rect 26712 12374 26740 18090
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26896 16425 26924 16594
rect 26882 16416 26938 16425
rect 26882 16351 26938 16360
rect 26790 16144 26846 16153
rect 26790 16079 26846 16088
rect 26804 13938 26832 16079
rect 26988 15638 27016 18255
rect 28184 18086 28212 18702
rect 28172 18080 28224 18086
rect 28172 18022 28224 18028
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27448 17066 27476 17614
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 27436 17060 27488 17066
rect 27436 17002 27488 17008
rect 26976 15632 27028 15638
rect 26976 15574 27028 15580
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26792 13728 26844 13734
rect 26792 13670 26844 13676
rect 26804 13376 26832 13670
rect 26896 13530 26924 14418
rect 26988 13530 27016 15302
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27172 14074 27200 14350
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 26884 13524 26936 13530
rect 26884 13466 26936 13472
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26884 13388 26936 13394
rect 26804 13348 26884 13376
rect 26884 13330 26936 13336
rect 26896 12986 26924 13330
rect 26884 12980 26936 12986
rect 26884 12922 26936 12928
rect 26988 12918 27016 13466
rect 27068 13320 27120 13326
rect 27068 13262 27120 13268
rect 26976 12912 27028 12918
rect 26882 12880 26938 12889
rect 26976 12854 27028 12860
rect 27080 12850 27108 13262
rect 26882 12815 26938 12824
rect 27068 12844 27120 12850
rect 26700 12368 26752 12374
rect 26700 12310 26752 12316
rect 26896 12306 26924 12815
rect 27068 12786 27120 12792
rect 27066 12608 27122 12617
rect 27066 12543 27122 12552
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26698 12200 26754 12209
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26436 11694 26464 12106
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26528 11354 26556 12038
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26344 11206 26464 11234
rect 26332 11076 26384 11082
rect 26332 11018 26384 11024
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 25962 10704 26018 10713
rect 25962 10639 26018 10648
rect 25976 10606 26004 10639
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 25594 10024 25650 10033
rect 25594 9959 25650 9968
rect 25424 9710 25544 9738
rect 25516 9625 25544 9710
rect 25502 9616 25558 9625
rect 25332 9574 25452 9602
rect 25226 9551 25282 9560
rect 25318 9480 25374 9489
rect 25318 9415 25374 9424
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25240 8634 25268 8910
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25332 8430 25360 9415
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 25318 7984 25374 7993
rect 25318 7919 25320 7928
rect 25372 7919 25374 7928
rect 25320 7890 25372 7896
rect 25332 7546 25360 7890
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25424 3913 25452 9574
rect 25502 9551 25558 9560
rect 25502 9344 25558 9353
rect 25502 9279 25558 9288
rect 25516 8634 25544 9279
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25608 8090 25636 9959
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26344 9194 26372 11018
rect 26160 9178 26372 9194
rect 26148 9172 26372 9178
rect 26200 9166 26372 9172
rect 26148 9114 26200 9120
rect 25686 9072 25742 9081
rect 26436 9058 26464 11206
rect 26620 10130 26648 12174
rect 26698 12135 26754 12144
rect 26712 10538 26740 12135
rect 26896 11626 26924 12242
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26976 11552 27028 11558
rect 26976 11494 27028 11500
rect 26882 11384 26938 11393
rect 26882 11319 26938 11328
rect 26896 11286 26924 11319
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 26896 10810 26924 11222
rect 26988 11150 27016 11494
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 26700 10532 26752 10538
rect 26700 10474 26752 10480
rect 26712 10266 26740 10474
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26608 10124 26660 10130
rect 26608 10066 26660 10072
rect 26620 9722 26648 10066
rect 26608 9716 26660 9722
rect 26608 9658 26660 9664
rect 26896 9654 26924 10746
rect 26988 10674 27016 11086
rect 26976 10668 27028 10674
rect 26976 10610 27028 10616
rect 26988 10266 27016 10610
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 26976 9920 27028 9926
rect 26976 9862 27028 9868
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 25686 9007 25742 9016
rect 26344 9030 26464 9058
rect 26516 9036 26568 9042
rect 25700 8498 25728 9007
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 25778 8256 25834 8265
rect 25778 8191 25834 8200
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25410 3904 25466 3913
rect 25410 3839 25466 3848
rect 25792 3505 25820 8191
rect 26344 8090 26372 9030
rect 26516 8978 26568 8984
rect 26422 8936 26478 8945
rect 26422 8871 26478 8880
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 26344 5250 26372 7686
rect 26436 7342 26464 8871
rect 26528 8634 26556 8978
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26528 8537 26556 8570
rect 26608 8560 26660 8566
rect 26514 8528 26570 8537
rect 26608 8502 26660 8508
rect 26514 8463 26570 8472
rect 26620 8401 26648 8502
rect 26606 8392 26662 8401
rect 26606 8327 26662 8336
rect 26712 8265 26740 8774
rect 26698 8256 26754 8265
rect 26698 8191 26754 8200
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26528 6866 26556 8026
rect 26606 6896 26662 6905
rect 26516 6860 26568 6866
rect 26606 6831 26662 6840
rect 26516 6802 26568 6808
rect 26528 6390 26556 6802
rect 26620 6458 26648 6831
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26516 6384 26568 6390
rect 26712 6361 26740 6598
rect 26516 6326 26568 6332
rect 26698 6352 26754 6361
rect 26698 6287 26754 6296
rect 26514 5808 26570 5817
rect 26514 5743 26516 5752
rect 26568 5743 26570 5752
rect 26516 5714 26568 5720
rect 26528 5370 26556 5714
rect 26698 5672 26754 5681
rect 26698 5607 26700 5616
rect 26752 5607 26754 5616
rect 26700 5578 26752 5584
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 25884 5222 26372 5250
rect 26422 5264 26478 5273
rect 25778 3496 25834 3505
rect 25778 3431 25834 3440
rect 25884 1465 25912 5222
rect 26422 5199 26478 5208
rect 26436 5166 26464 5199
rect 26424 5160 26476 5166
rect 26424 5102 26476 5108
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26620 5030 26648 5063
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26804 4185 26832 9318
rect 26884 7200 26936 7206
rect 26884 7142 26936 7148
rect 26790 4176 26846 4185
rect 26790 4111 26846 4120
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26422 3088 26478 3097
rect 26422 3023 26478 3032
rect 26436 2990 26464 3023
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26608 2848 26660 2854
rect 26606 2816 26608 2825
rect 26660 2816 26662 2825
rect 26606 2751 26662 2760
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 25870 1456 25926 1465
rect 25870 1391 25926 1400
rect 2226 368 2282 377
rect 2226 303 2282 312
rect 4986 0 5042 480
rect 14922 0 14978 480
rect 24950 0 25006 480
rect 26896 377 26924 7142
rect 26988 6338 27016 9862
rect 27080 7954 27108 12543
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27172 11898 27200 12174
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 27080 7546 27108 7890
rect 27068 7540 27120 7546
rect 27068 7482 27120 7488
rect 26988 6310 27108 6338
rect 27172 6322 27200 10542
rect 27264 8566 27292 17002
rect 27448 15484 27476 17002
rect 27540 16250 27568 17138
rect 27816 16998 27844 17682
rect 28184 17202 28212 18022
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27528 15496 27580 15502
rect 27448 15456 27528 15484
rect 27528 15438 27580 15444
rect 27540 14822 27568 15438
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27342 14104 27398 14113
rect 27342 14039 27398 14048
rect 27356 12209 27384 14039
rect 27540 13938 27568 14758
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27540 13841 27568 13874
rect 27526 13832 27582 13841
rect 27526 13767 27582 13776
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 27632 12850 27660 13738
rect 27724 13530 27752 13874
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27816 13433 27844 16934
rect 27802 13424 27858 13433
rect 27802 13359 27858 13368
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27436 12368 27488 12374
rect 27436 12310 27488 12316
rect 27342 12200 27398 12209
rect 27342 12135 27398 12144
rect 27448 9738 27476 12310
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27632 10810 27660 11290
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27526 10160 27582 10169
rect 27526 10095 27582 10104
rect 27356 9710 27476 9738
rect 27356 9081 27384 9710
rect 27434 9616 27490 9625
rect 27434 9551 27490 9560
rect 27448 9518 27476 9551
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27342 9072 27398 9081
rect 27342 9007 27398 9016
rect 27252 8560 27304 8566
rect 27252 8502 27304 8508
rect 27540 8430 27568 10095
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27710 8664 27766 8673
rect 27710 8599 27712 8608
rect 27764 8599 27766 8608
rect 27712 8570 27764 8576
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27712 7472 27764 7478
rect 27526 7440 27582 7449
rect 27526 7375 27582 7384
rect 27710 7440 27712 7449
rect 27764 7440 27766 7449
rect 27710 7375 27766 7384
rect 27540 7342 27568 7375
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 26974 4176 27030 4185
rect 26974 4111 27030 4120
rect 26988 2145 27016 4111
rect 26974 2136 27030 2145
rect 26974 2071 27030 2080
rect 27080 921 27108 6310
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27816 4457 27844 9318
rect 27802 4448 27858 4457
rect 27802 4383 27858 4392
rect 27066 912 27122 921
rect 27066 847 27122 856
rect 26882 368 26938 377
rect 26882 303 26938 312
<< via2 >>
rect 2962 23568 3018 23624
rect 1398 20440 1454 20496
rect 1122 15272 1178 15328
rect 1766 16768 1822 16824
rect 2226 14048 2282 14104
rect 1582 13368 1638 13424
rect 1214 12280 1270 12336
rect 1674 10260 1730 10296
rect 1674 10240 1676 10260
rect 1676 10240 1728 10260
rect 1728 10240 1730 10260
rect 1582 7420 1584 7440
rect 1584 7420 1636 7440
rect 1636 7420 1638 7440
rect 1582 7384 1638 7420
rect 1582 6840 1638 6896
rect 1582 6332 1584 6352
rect 1584 6332 1636 6352
rect 1636 6332 1638 6352
rect 1582 6296 1638 6332
rect 1582 5636 1638 5672
rect 1582 5616 1584 5636
rect 1584 5616 1636 5636
rect 1636 5616 1638 5636
rect 1582 5072 1638 5128
rect 1766 7248 1822 7304
rect 2042 13504 2098 13560
rect 2134 12552 2190 12608
rect 2134 10532 2190 10568
rect 2134 10512 2136 10532
rect 2136 10512 2188 10532
rect 2188 10512 2190 10532
rect 25042 23568 25098 23624
rect 3330 23024 3386 23080
rect 3146 22344 3202 22400
rect 2962 19488 3018 19544
rect 2778 16652 2834 16688
rect 2778 16632 2780 16652
rect 2780 16632 2832 16652
rect 2832 16632 2834 16652
rect 2594 15952 2650 16008
rect 2870 13912 2926 13968
rect 2594 13640 2650 13696
rect 2594 11212 2650 11248
rect 2594 11192 2596 11212
rect 2596 11192 2648 11212
rect 2648 11192 2650 11212
rect 2594 9696 2650 9752
rect 2502 8064 2558 8120
rect 2042 6432 2098 6488
rect 2042 5228 2098 5264
rect 2042 5208 2044 5228
rect 2044 5208 2096 5228
rect 2096 5208 2098 5228
rect 1674 4392 1730 4448
rect 2042 3984 2098 4040
rect 1490 3848 1546 3904
rect 1582 2624 1638 2680
rect 2870 12300 2926 12336
rect 2870 12280 2872 12300
rect 2872 12280 2924 12300
rect 2924 12280 2926 12300
rect 4066 21800 4122 21856
rect 4434 21256 4490 21312
rect 3606 20576 3662 20632
rect 3330 15816 3386 15872
rect 3330 14048 3386 14104
rect 3790 17040 3846 17096
rect 3882 16904 3938 16960
rect 3790 16088 3846 16144
rect 3514 14456 3570 14512
rect 2870 10804 2926 10840
rect 2870 10784 2872 10804
rect 2872 10784 2924 10804
rect 2924 10784 2926 10804
rect 2778 9036 2834 9072
rect 2778 9016 2780 9036
rect 2780 9016 2832 9036
rect 2832 9016 2834 9036
rect 3330 10240 3386 10296
rect 3882 14220 3884 14240
rect 3884 14220 3936 14240
rect 3936 14220 3938 14240
rect 3882 14184 3938 14220
rect 4066 18264 4122 18320
rect 4158 14320 4214 14376
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 4986 20476 4988 20496
rect 4988 20476 5040 20496
rect 5040 20476 5042 20496
rect 4986 20440 5042 20476
rect 4618 19488 4674 19544
rect 4802 19216 4858 19272
rect 4618 17856 4674 17912
rect 4434 16788 4490 16824
rect 4434 16768 4436 16788
rect 4436 16768 4488 16788
rect 4488 16768 4490 16788
rect 4434 15544 4490 15600
rect 4342 14728 4398 14784
rect 4250 12552 4306 12608
rect 4986 18028 4988 18048
rect 4988 18028 5040 18048
rect 5040 18028 5042 18048
rect 4986 17992 5042 18028
rect 5078 16360 5134 16416
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 6550 20440 6606 20496
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 6734 19080 6790 19136
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5722 18128 5778 18184
rect 4066 11600 4122 11656
rect 3698 10512 3754 10568
rect 3514 9968 3570 10024
rect 3606 9696 3662 9752
rect 3146 6840 3202 6896
rect 4250 11056 4306 11112
rect 4066 10376 4122 10432
rect 4066 9288 4122 9344
rect 3790 8880 3846 8936
rect 4250 8608 4306 8664
rect 4434 12280 4490 12336
rect 4526 12144 4582 12200
rect 5630 15544 5686 15600
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 6550 15852 6552 15872
rect 6552 15852 6604 15872
rect 6604 15852 6606 15872
rect 6550 15816 6606 15852
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5814 15000 5870 15056
rect 5722 14184 5778 14240
rect 5630 13504 5686 13560
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5262 13268 5264 13288
rect 5264 13268 5316 13288
rect 5316 13268 5318 13288
rect 5262 13232 5318 13268
rect 5170 11328 5226 11384
rect 5814 13504 5870 13560
rect 5630 12688 5686 12744
rect 5446 9832 5502 9888
rect 5446 8336 5502 8392
rect 5170 6840 5226 6896
rect 3514 6196 3516 6216
rect 3516 6196 3568 6216
rect 3568 6196 3570 6216
rect 3514 6160 3570 6196
rect 2502 5772 2558 5808
rect 2502 5752 2504 5772
rect 2504 5752 2556 5772
rect 2556 5752 2558 5772
rect 6182 13640 6238 13696
rect 5814 13096 5870 13152
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 6366 13096 6422 13152
rect 6274 12824 6330 12880
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 5354 6432 5410 6488
rect 3790 3304 3846 3360
rect 7470 17992 7526 18048
rect 7746 17176 7802 17232
rect 7746 16632 7802 16688
rect 7194 15408 7250 15464
rect 7286 14184 7342 14240
rect 7562 13504 7618 13560
rect 7654 13368 7710 13424
rect 7102 11500 7104 11520
rect 7104 11500 7156 11520
rect 7156 11500 7158 11520
rect 7102 11464 7158 11500
rect 6918 11348 6974 11384
rect 6918 11328 6920 11348
rect 6920 11328 6972 11348
rect 6972 11328 6974 11348
rect 7746 13096 7802 13152
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 9586 19488 9642 19544
rect 9034 19116 9036 19136
rect 9036 19116 9088 19136
rect 9088 19116 9090 19136
rect 9034 19080 9090 19116
rect 8022 17584 8078 17640
rect 8298 17856 8354 17912
rect 8390 17448 8446 17504
rect 8298 16632 8354 16688
rect 9862 16940 9864 16960
rect 9864 16940 9916 16960
rect 9916 16940 9918 16960
rect 9862 16904 9918 16940
rect 8022 15272 8078 15328
rect 8942 16088 8998 16144
rect 8390 15136 8446 15192
rect 8298 13232 8354 13288
rect 7470 10648 7526 10704
rect 7286 9968 7342 10024
rect 7562 9968 7618 10024
rect 7838 10124 7894 10160
rect 7838 10104 7840 10124
rect 7840 10104 7892 10124
rect 7892 10104 7894 10124
rect 7194 8372 7196 8392
rect 7196 8372 7248 8392
rect 7248 8372 7250 8392
rect 7194 8336 7250 8372
rect 9034 14340 9090 14376
rect 9034 14320 9036 14340
rect 9036 14320 9088 14340
rect 9088 14320 9090 14340
rect 9494 14864 9550 14920
rect 9402 14764 9404 14784
rect 9404 14764 9456 14784
rect 9456 14764 9458 14784
rect 9402 14728 9458 14764
rect 9310 14320 9366 14376
rect 9218 10920 9274 10976
rect 9862 14456 9918 14512
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10322 19896 10378 19952
rect 10138 18808 10194 18864
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10138 13776 10194 13832
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 11610 18808 11666 18864
rect 11794 18808 11850 18864
rect 11610 16496 11666 16552
rect 11426 15544 11482 15600
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 10782 12588 10784 12608
rect 10784 12588 10836 12608
rect 10836 12588 10838 12608
rect 10782 12552 10838 12588
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10138 11464 10194 11520
rect 10782 12144 10838 12200
rect 9770 10784 9826 10840
rect 9678 10648 9734 10704
rect 8574 9560 8630 9616
rect 8298 9016 8354 9072
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 7194 6840 7250 6896
rect 5814 5752 5870 5808
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 7838 3984 7894 4040
rect 6918 3032 6974 3088
rect 8574 5208 8630 5264
rect 7194 2352 7250 2408
rect 4066 2080 4122 2136
rect 2686 1400 2742 1456
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 11610 12588 11612 12608
rect 11612 12588 11664 12608
rect 11664 12588 11666 12608
rect 11610 12552 11666 12588
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 14554 20324 14610 20360
rect 14554 20304 14556 20324
rect 14556 20304 14608 20324
rect 14608 20304 14610 20324
rect 12438 19896 12494 19952
rect 13634 19896 13690 19952
rect 12162 19488 12218 19544
rect 11978 17584 12034 17640
rect 11794 12824 11850 12880
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10690 9424 10746 9480
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 12898 19216 12954 19272
rect 13542 19116 13544 19136
rect 13544 19116 13596 19136
rect 13596 19116 13598 19136
rect 13542 19080 13598 19116
rect 12162 16632 12218 16688
rect 12162 15544 12218 15600
rect 12070 14184 12126 14240
rect 12254 15272 12310 15328
rect 12898 16940 12900 16960
rect 12900 16940 12952 16960
rect 12952 16940 12954 16960
rect 12898 16904 12954 16940
rect 14554 19624 14610 19680
rect 12622 15408 12678 15464
rect 12530 14864 12586 14920
rect 12438 13776 12494 13832
rect 12162 13504 12218 13560
rect 12806 13504 12862 13560
rect 13174 15156 13230 15192
rect 13174 15136 13176 15156
rect 13176 15136 13228 15156
rect 13228 15136 13230 15156
rect 13174 14456 13230 14512
rect 12898 13096 12954 13152
rect 12806 12824 12862 12880
rect 13082 11192 13138 11248
rect 13450 11192 13506 11248
rect 12254 10920 12310 10976
rect 14094 17584 14150 17640
rect 14370 17584 14426 17640
rect 13818 15544 13874 15600
rect 13910 14864 13966 14920
rect 14922 17448 14978 17504
rect 14646 16124 14648 16144
rect 14648 16124 14700 16144
rect 14700 16124 14702 16144
rect 14646 16088 14702 16124
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 17958 19760 18014 19816
rect 16394 19352 16450 19408
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15290 16632 15346 16688
rect 15014 16360 15070 16416
rect 14922 15680 14978 15736
rect 15014 15408 15070 15464
rect 14738 14320 14794 14376
rect 14922 13368 14978 13424
rect 16302 17720 16358 17776
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 15658 16360 15714 16416
rect 15290 11328 15346 11384
rect 14830 11056 14886 11112
rect 13542 10512 13598 10568
rect 15474 13812 15476 13832
rect 15476 13812 15528 13832
rect 15528 13812 15530 13832
rect 15474 13776 15530 13812
rect 15566 12552 15622 12608
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 16394 16244 16450 16280
rect 16394 16224 16396 16244
rect 16396 16224 16448 16244
rect 16448 16224 16450 16244
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 16394 14592 16450 14648
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 16486 14456 16542 14512
rect 16486 13912 16542 13968
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15382 9560 15438 9616
rect 13450 8472 13506 8528
rect 11886 7248 11942 7304
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 16486 13096 16542 13152
rect 17130 17584 17186 17640
rect 17314 17040 17370 17096
rect 17130 16496 17186 16552
rect 17958 17720 18014 17776
rect 17314 16360 17370 16416
rect 17498 16496 17554 16552
rect 17498 16224 17554 16280
rect 18142 17312 18198 17368
rect 18234 15408 18290 15464
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15750 10512 15806 10568
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 17038 9968 17094 10024
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 17406 10104 17462 10160
rect 19522 19896 19578 19952
rect 19614 19760 19670 19816
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 20534 19080 20590 19136
rect 20534 18264 20590 18320
rect 18602 15952 18658 16008
rect 20534 17720 20590 17776
rect 18510 15680 18566 15736
rect 18510 15408 18566 15464
rect 18510 15000 18566 15056
rect 19062 15020 19118 15056
rect 19062 15000 19064 15020
rect 19064 15000 19116 15020
rect 19116 15000 19118 15020
rect 19614 14864 19670 14920
rect 18602 14184 18658 14240
rect 18510 12008 18566 12064
rect 18326 11056 18382 11112
rect 18418 9580 18474 9616
rect 18418 9560 18420 9580
rect 18420 9560 18472 9580
rect 18472 9560 18474 9580
rect 20442 14592 20498 14648
rect 19246 14048 19302 14104
rect 18694 12960 18750 13016
rect 18694 12688 18750 12744
rect 18878 13504 18934 13560
rect 18878 13232 18934 13288
rect 18786 11192 18842 11248
rect 19614 13812 19616 13832
rect 19616 13812 19668 13832
rect 19668 13812 19670 13832
rect 19614 13776 19670 13812
rect 19338 12824 19394 12880
rect 19062 12708 19118 12744
rect 19062 12688 19064 12708
rect 19064 12688 19116 12708
rect 19116 12688 19118 12708
rect 19338 12144 19394 12200
rect 19246 11464 19302 11520
rect 19614 12008 19670 12064
rect 19706 11328 19762 11384
rect 19890 13776 19946 13832
rect 19890 11192 19946 11248
rect 19982 10548 19984 10568
rect 19984 10548 20036 10568
rect 20036 10548 20038 10568
rect 19982 10512 20038 10548
rect 20350 13368 20406 13424
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 20810 18148 20866 18184
rect 20810 18128 20812 18148
rect 20812 18128 20864 18148
rect 20864 18128 20866 18148
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 21362 19896 21418 19952
rect 24950 21528 25006 21584
rect 22006 19488 22062 19544
rect 23386 19488 23442 19544
rect 21454 19216 21510 19272
rect 21270 17040 21326 17096
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20350 10784 20406 10840
rect 21638 17720 21694 17776
rect 21638 17448 21694 17504
rect 22466 19352 22522 19408
rect 23110 18808 23166 18864
rect 21454 15036 21456 15056
rect 21456 15036 21508 15056
rect 21508 15036 21510 15056
rect 21454 15000 21510 15036
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20810 11464 20866 11520
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 21822 16088 21878 16144
rect 21546 12280 21602 12336
rect 21362 11600 21418 11656
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 21822 12960 21878 13016
rect 21730 12416 21786 12472
rect 22190 13368 22246 13424
rect 22466 12588 22468 12608
rect 22468 12588 22520 12608
rect 22520 12588 22522 12608
rect 22466 12552 22522 12588
rect 22006 10784 22062 10840
rect 21454 9444 21510 9480
rect 21454 9424 21456 9444
rect 21456 9424 21508 9444
rect 21508 9424 21510 9444
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 20166 8880 20222 8936
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 23110 17720 23166 17776
rect 23754 15408 23810 15464
rect 23662 14492 23664 14512
rect 23664 14492 23716 14512
rect 23716 14492 23718 14512
rect 23662 14456 23718 14492
rect 23478 13096 23534 13152
rect 23754 11056 23810 11112
rect 24398 18264 24454 18320
rect 23938 18028 23940 18048
rect 23940 18028 23992 18048
rect 23992 18028 23994 18048
rect 23938 17992 23994 18028
rect 24030 14184 24086 14240
rect 23938 13796 23994 13832
rect 23938 13776 23940 13796
rect 23940 13776 23992 13796
rect 23992 13776 23994 13796
rect 24306 13096 24362 13152
rect 24122 12416 24178 12472
rect 24122 12300 24178 12336
rect 24122 12280 24124 12300
rect 24124 12280 24176 12300
rect 24176 12280 24178 12300
rect 25410 23024 25466 23080
rect 25134 20440 25190 20496
rect 24950 18808 25006 18864
rect 25042 17176 25098 17232
rect 24950 16360 25006 16416
rect 24674 14320 24730 14376
rect 25686 22344 25742 22400
rect 25502 21256 25558 21312
rect 25226 18944 25282 19000
rect 25226 18808 25282 18864
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25686 18400 25742 18456
rect 26514 18944 26570 19000
rect 25226 17720 25282 17776
rect 25318 17332 25374 17368
rect 25318 17312 25320 17332
rect 25320 17312 25372 17332
rect 25372 17312 25374 17332
rect 25134 15816 25190 15872
rect 25042 14592 25098 14648
rect 24766 12280 24822 12336
rect 24950 12280 25006 12336
rect 24766 12008 24822 12064
rect 22650 7928 22706 7984
rect 25134 14048 25190 14104
rect 25134 10376 25190 10432
rect 25042 9968 25098 10024
rect 24306 7384 24362 7440
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 18234 6160 18290 6216
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 17314 5752 17370 5808
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 15566 5208 15622 5264
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 14922 2352 14978 2408
rect 10414 1264 10470 1320
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 25502 16124 25504 16144
rect 25504 16124 25556 16144
rect 25556 16124 25558 16144
rect 25502 16088 25558 16124
rect 25318 15408 25374 15464
rect 25226 9560 25282 9616
rect 25502 12688 25558 12744
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25686 13912 25742 13968
rect 25410 12008 25466 12064
rect 26422 16632 26478 16688
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 26238 15408 26294 15464
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 26974 20032 27030 20088
rect 26974 19760 27030 19816
rect 26974 18264 27030 18320
rect 26606 14356 26608 14376
rect 26608 14356 26660 14376
rect 26660 14356 26662 14376
rect 26606 14320 26662 14356
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 25778 11328 25834 11384
rect 26882 16360 26938 16416
rect 26790 16088 26846 16144
rect 26882 12824 26938 12880
rect 27066 12552 27122 12608
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 25962 10648 26018 10704
rect 25594 9968 25650 10024
rect 25318 9424 25374 9480
rect 25318 7948 25374 7984
rect 25318 7928 25320 7948
rect 25320 7928 25372 7948
rect 25372 7928 25374 7948
rect 25502 9560 25558 9616
rect 25502 9288 25558 9344
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 25686 9016 25742 9072
rect 26698 12144 26754 12200
rect 26882 11328 26938 11384
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25778 8200 25834 8256
rect 25410 3848 25466 3904
rect 26422 8880 26478 8936
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 26514 8472 26570 8528
rect 26606 8336 26662 8392
rect 26698 8200 26754 8256
rect 26606 6840 26662 6896
rect 26698 6296 26754 6352
rect 26514 5772 26570 5808
rect 26514 5752 26516 5772
rect 26516 5752 26568 5772
rect 26568 5752 26570 5772
rect 26698 5636 26754 5672
rect 26698 5616 26700 5636
rect 26700 5616 26752 5636
rect 26752 5616 26754 5636
rect 25778 3440 25834 3496
rect 26422 5208 26478 5264
rect 26606 5072 26662 5128
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26790 4120 26846 4176
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 26422 3032 26478 3088
rect 26606 2796 26608 2816
rect 26608 2796 26660 2816
rect 26660 2796 26662 2816
rect 26606 2760 26662 2796
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 1400 25926 1456
rect 2226 312 2282 368
rect 27342 14048 27398 14104
rect 27526 13776 27582 13832
rect 27802 13368 27858 13424
rect 27342 12144 27398 12200
rect 27526 10104 27582 10160
rect 27434 9560 27490 9616
rect 27342 9016 27398 9072
rect 27710 8628 27766 8664
rect 27710 8608 27712 8628
rect 27712 8608 27764 8628
rect 27764 8608 27766 8628
rect 27526 7384 27582 7440
rect 27710 7420 27712 7440
rect 27712 7420 27764 7440
rect 27764 7420 27766 7440
rect 27710 7384 27766 7420
rect 26974 4120 27030 4176
rect 26974 2080 27030 2136
rect 27802 4392 27858 4448
rect 27066 856 27122 912
rect 26882 312 26938 368
<< metal3 >>
rect 0 23626 480 23656
rect 2957 23626 3023 23629
rect 0 23624 3023 23626
rect 0 23568 2962 23624
rect 3018 23568 3023 23624
rect 0 23566 3023 23568
rect 0 23536 480 23566
rect 2957 23563 3023 23566
rect 25037 23626 25103 23629
rect 29520 23626 30000 23656
rect 25037 23624 30000 23626
rect 25037 23568 25042 23624
rect 25098 23568 30000 23624
rect 25037 23566 30000 23568
rect 25037 23563 25103 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3325 23082 3391 23085
rect 0 23080 3391 23082
rect 0 23024 3330 23080
rect 3386 23024 3391 23080
rect 0 23022 3391 23024
rect 0 22992 480 23022
rect 3325 23019 3391 23022
rect 25405 23082 25471 23085
rect 29520 23082 30000 23112
rect 25405 23080 30000 23082
rect 25405 23024 25410 23080
rect 25466 23024 30000 23080
rect 25405 23022 30000 23024
rect 25405 23019 25471 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 3141 22402 3207 22405
rect 0 22400 3207 22402
rect 0 22344 3146 22400
rect 3202 22344 3207 22400
rect 0 22342 3207 22344
rect 0 22312 480 22342
rect 3141 22339 3207 22342
rect 25681 22402 25747 22405
rect 29520 22402 30000 22432
rect 25681 22400 30000 22402
rect 25681 22344 25686 22400
rect 25742 22344 30000 22400
rect 25681 22342 30000 22344
rect 25681 22339 25747 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 4061 21858 4127 21861
rect 29520 21858 30000 21888
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 480 21798
rect 4061 21795 4127 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 24945 21586 25011 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 24945 21584 26434 21586
rect 24945 21528 24950 21584
rect 25006 21528 26434 21584
rect 24945 21526 26434 21528
rect 24945 21523 25011 21526
rect 0 21314 480 21344
rect 4429 21314 4495 21317
rect 0 21312 4495 21314
rect 0 21256 4434 21312
rect 4490 21256 4495 21312
rect 0 21254 4495 21256
rect 0 21224 480 21254
rect 4429 21251 4495 21254
rect 25497 21314 25563 21317
rect 29520 21314 30000 21344
rect 25497 21312 30000 21314
rect 25497 21256 25502 21312
rect 25558 21256 30000 21312
rect 25497 21254 30000 21256
rect 25497 21251 25563 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3601 20634 3667 20637
rect 29520 20634 30000 20664
rect 0 20632 3667 20634
rect 0 20576 3606 20632
rect 3662 20576 3667 20632
rect 0 20574 3667 20576
rect 0 20544 480 20574
rect 3601 20571 3667 20574
rect 26374 20574 30000 20634
rect 1393 20498 1459 20501
rect 4981 20498 5047 20501
rect 6545 20498 6611 20501
rect 1393 20496 2882 20498
rect 1393 20440 1398 20496
rect 1454 20440 2882 20496
rect 1393 20438 2882 20440
rect 1393 20435 1459 20438
rect 2822 20362 2882 20438
rect 4981 20496 6611 20498
rect 4981 20440 4986 20496
rect 5042 20440 6550 20496
rect 6606 20440 6611 20496
rect 4981 20438 6611 20440
rect 4981 20435 5047 20438
rect 6545 20435 6611 20438
rect 25129 20498 25195 20501
rect 26374 20498 26434 20574
rect 29520 20544 30000 20574
rect 25129 20496 26434 20498
rect 25129 20440 25134 20496
rect 25190 20440 26434 20496
rect 25129 20438 26434 20440
rect 25129 20435 25195 20438
rect 14549 20362 14615 20365
rect 2822 20360 14615 20362
rect 2822 20304 14554 20360
rect 14610 20304 14615 20360
rect 2822 20302 14615 20304
rect 14549 20299 14615 20302
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 26969 20090 27035 20093
rect 29520 20090 30000 20120
rect 0 20030 2698 20090
rect 0 20000 480 20030
rect 2638 19954 2698 20030
rect 26969 20088 30000 20090
rect 26969 20032 26974 20088
rect 27030 20032 30000 20088
rect 26969 20030 30000 20032
rect 26969 20027 27035 20030
rect 29520 20000 30000 20030
rect 10317 19954 10383 19957
rect 12433 19954 12499 19957
rect 2638 19894 2882 19954
rect 2822 19818 2882 19894
rect 10317 19952 12499 19954
rect 10317 19896 10322 19952
rect 10378 19896 12438 19952
rect 12494 19896 12499 19952
rect 10317 19894 12499 19896
rect 10317 19891 10383 19894
rect 12433 19891 12499 19894
rect 13629 19954 13695 19957
rect 19517 19954 19583 19957
rect 21357 19954 21423 19957
rect 13629 19952 21423 19954
rect 13629 19896 13634 19952
rect 13690 19896 19522 19952
rect 19578 19896 21362 19952
rect 21418 19896 21423 19952
rect 13629 19894 21423 19896
rect 13629 19891 13695 19894
rect 19517 19891 19583 19894
rect 21357 19891 21423 19894
rect 17953 19818 18019 19821
rect 2822 19816 18019 19818
rect 2822 19760 17958 19816
rect 18014 19760 18019 19816
rect 2822 19758 18019 19760
rect 17953 19755 18019 19758
rect 19609 19818 19675 19821
rect 26969 19818 27035 19821
rect 19609 19816 27035 19818
rect 19609 19760 19614 19816
rect 19670 19760 26974 19816
rect 27030 19760 27035 19816
rect 19609 19758 27035 19760
rect 19609 19755 19675 19758
rect 26969 19755 27035 19758
rect 9622 19620 9628 19684
rect 9692 19682 9698 19684
rect 14549 19682 14615 19685
rect 9692 19680 14615 19682
rect 9692 19624 14554 19680
rect 14610 19624 14615 19680
rect 9692 19622 14615 19624
rect 9692 19620 9698 19622
rect 14549 19619 14615 19622
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 2957 19546 3023 19549
rect 4613 19546 4679 19549
rect 2957 19544 4679 19546
rect 2957 19488 2962 19544
rect 3018 19488 4618 19544
rect 4674 19488 4679 19544
rect 2957 19486 4679 19488
rect 2957 19483 3023 19486
rect 4613 19483 4679 19486
rect 9581 19546 9647 19549
rect 12157 19546 12223 19549
rect 9581 19544 12223 19546
rect 9581 19488 9586 19544
rect 9642 19488 12162 19544
rect 12218 19488 12223 19544
rect 9581 19486 12223 19488
rect 9581 19483 9647 19486
rect 12157 19483 12223 19486
rect 22001 19546 22067 19549
rect 23381 19546 23447 19549
rect 22001 19544 23447 19546
rect 22001 19488 22006 19544
rect 22062 19488 23386 19544
rect 23442 19488 23447 19544
rect 22001 19486 23447 19488
rect 22001 19483 22067 19486
rect 23381 19483 23447 19486
rect 0 19410 480 19440
rect 9622 19410 9628 19412
rect 0 19350 9628 19410
rect 0 19320 480 19350
rect 9622 19348 9628 19350
rect 9692 19348 9698 19412
rect 16389 19410 16455 19413
rect 22461 19410 22527 19413
rect 29520 19410 30000 19440
rect 16389 19408 21466 19410
rect 16389 19352 16394 19408
rect 16450 19352 21466 19408
rect 16389 19350 21466 19352
rect 16389 19347 16455 19350
rect 21406 19277 21466 19350
rect 22461 19408 30000 19410
rect 22461 19352 22466 19408
rect 22522 19352 30000 19408
rect 22461 19350 30000 19352
rect 22461 19347 22527 19350
rect 29520 19320 30000 19350
rect 4797 19274 4863 19277
rect 12893 19274 12959 19277
rect 4797 19272 12959 19274
rect 4797 19216 4802 19272
rect 4858 19216 12898 19272
rect 12954 19216 12959 19272
rect 4797 19214 12959 19216
rect 21406 19272 21515 19277
rect 21406 19216 21454 19272
rect 21510 19216 21515 19272
rect 21406 19214 21515 19216
rect 4797 19211 4863 19214
rect 12893 19211 12959 19214
rect 21449 19211 21515 19214
rect 6729 19138 6795 19141
rect 9029 19138 9095 19141
rect 6729 19136 9095 19138
rect 6729 19080 6734 19136
rect 6790 19080 9034 19136
rect 9090 19080 9095 19136
rect 6729 19078 9095 19080
rect 6729 19075 6795 19078
rect 9029 19075 9095 19078
rect 13537 19138 13603 19141
rect 20529 19138 20595 19141
rect 13537 19136 20595 19138
rect 13537 19080 13542 19136
rect 13598 19080 20534 19136
rect 20590 19080 20595 19136
rect 13537 19078 20595 19080
rect 13537 19075 13603 19078
rect 20529 19075 20595 19078
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 25221 19002 25287 19005
rect 26509 19002 26575 19005
rect 25221 19000 26575 19002
rect 25221 18944 25226 19000
rect 25282 18944 26514 19000
rect 26570 18944 26575 19000
rect 25221 18942 26575 18944
rect 25221 18939 25287 18942
rect 26509 18939 26575 18942
rect 0 18866 480 18896
rect 10133 18866 10199 18869
rect 11605 18866 11671 18869
rect 0 18864 11671 18866
rect 0 18808 10138 18864
rect 10194 18808 11610 18864
rect 11666 18808 11671 18864
rect 0 18806 11671 18808
rect 0 18776 480 18806
rect 10133 18803 10199 18806
rect 11605 18803 11671 18806
rect 11789 18866 11855 18869
rect 23105 18866 23171 18869
rect 24945 18866 25011 18869
rect 11789 18864 25011 18866
rect 11789 18808 11794 18864
rect 11850 18808 23110 18864
rect 23166 18808 24950 18864
rect 25006 18808 25011 18864
rect 11789 18806 25011 18808
rect 11789 18803 11855 18806
rect 23105 18803 23171 18806
rect 24945 18803 25011 18806
rect 25221 18866 25287 18869
rect 29520 18866 30000 18896
rect 25221 18864 30000 18866
rect 25221 18808 25226 18864
rect 25282 18808 30000 18864
rect 25221 18806 30000 18808
rect 25221 18803 25287 18806
rect 29520 18776 30000 18806
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 25681 18458 25747 18461
rect 17174 18456 25747 18458
rect 17174 18400 25686 18456
rect 25742 18400 25747 18456
rect 17174 18398 25747 18400
rect 0 18322 480 18352
rect 4061 18322 4127 18325
rect 17174 18322 17234 18398
rect 25681 18395 25747 18398
rect 0 18262 2698 18322
rect 0 18232 480 18262
rect 2638 17914 2698 18262
rect 4061 18320 17234 18322
rect 4061 18264 4066 18320
rect 4122 18264 17234 18320
rect 4061 18262 17234 18264
rect 20529 18322 20595 18325
rect 24393 18322 24459 18325
rect 20529 18320 24459 18322
rect 20529 18264 20534 18320
rect 20590 18264 24398 18320
rect 24454 18264 24459 18320
rect 20529 18262 24459 18264
rect 4061 18259 4127 18262
rect 20529 18259 20595 18262
rect 24393 18259 24459 18262
rect 26969 18322 27035 18325
rect 29520 18322 30000 18352
rect 26969 18320 30000 18322
rect 26969 18264 26974 18320
rect 27030 18264 30000 18320
rect 26969 18262 30000 18264
rect 26969 18259 27035 18262
rect 29520 18232 30000 18262
rect 5717 18186 5783 18189
rect 20805 18186 20871 18189
rect 5717 18184 20871 18186
rect 5717 18128 5722 18184
rect 5778 18128 20810 18184
rect 20866 18128 20871 18184
rect 5717 18126 20871 18128
rect 5717 18123 5783 18126
rect 20805 18123 20871 18126
rect 4981 18050 5047 18053
rect 7465 18050 7531 18053
rect 23933 18050 23999 18053
rect 4981 18048 7531 18050
rect 4981 17992 4986 18048
rect 5042 17992 7470 18048
rect 7526 17992 7531 18048
rect 4981 17990 7531 17992
rect 4981 17987 5047 17990
rect 7465 17987 7531 17990
rect 21406 18048 23999 18050
rect 21406 17992 23938 18048
rect 23994 17992 23999 18048
rect 21406 17990 23999 17992
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 4613 17914 4679 17917
rect 8293 17914 8359 17917
rect 2638 17912 8359 17914
rect 2638 17856 4618 17912
rect 4674 17856 8298 17912
rect 8354 17856 8359 17912
rect 2638 17854 8359 17856
rect 4613 17851 4679 17854
rect 8293 17851 8359 17854
rect 16297 17778 16363 17781
rect 17953 17778 18019 17781
rect 16297 17776 18019 17778
rect 16297 17720 16302 17776
rect 16358 17720 17958 17776
rect 18014 17720 18019 17776
rect 16297 17718 18019 17720
rect 16297 17715 16363 17718
rect 17953 17715 18019 17718
rect 20529 17778 20595 17781
rect 21406 17778 21466 17990
rect 23933 17987 23999 17990
rect 20529 17776 21466 17778
rect 20529 17720 20534 17776
rect 20590 17720 21466 17776
rect 20529 17718 21466 17720
rect 21633 17778 21699 17781
rect 23105 17778 23171 17781
rect 25221 17778 25287 17781
rect 21633 17776 25287 17778
rect 21633 17720 21638 17776
rect 21694 17720 23110 17776
rect 23166 17720 25226 17776
rect 25282 17720 25287 17776
rect 21633 17718 25287 17720
rect 20529 17715 20595 17718
rect 21633 17715 21699 17718
rect 23105 17715 23171 17718
rect 25221 17715 25287 17718
rect 0 17642 480 17672
rect 8017 17642 8083 17645
rect 0 17640 8083 17642
rect 0 17584 8022 17640
rect 8078 17584 8083 17640
rect 0 17582 8083 17584
rect 0 17552 480 17582
rect 8017 17579 8083 17582
rect 11973 17642 12039 17645
rect 14089 17642 14155 17645
rect 11973 17640 14155 17642
rect 11973 17584 11978 17640
rect 12034 17584 14094 17640
rect 14150 17584 14155 17640
rect 11973 17582 14155 17584
rect 11973 17579 12039 17582
rect 14089 17579 14155 17582
rect 14365 17642 14431 17645
rect 17125 17642 17191 17645
rect 29520 17642 30000 17672
rect 14365 17640 16498 17642
rect 14365 17584 14370 17640
rect 14426 17584 16498 17640
rect 14365 17582 16498 17584
rect 14365 17579 14431 17582
rect 8385 17506 8451 17509
rect 14917 17506 14983 17509
rect 8385 17504 14983 17506
rect 8385 17448 8390 17504
rect 8446 17448 14922 17504
rect 14978 17448 14983 17504
rect 8385 17446 14983 17448
rect 16438 17506 16498 17582
rect 17125 17640 30000 17642
rect 17125 17584 17130 17640
rect 17186 17584 30000 17640
rect 17125 17582 30000 17584
rect 17125 17579 17191 17582
rect 29520 17552 30000 17582
rect 21633 17506 21699 17509
rect 16438 17504 21699 17506
rect 16438 17448 21638 17504
rect 21694 17448 21699 17504
rect 16438 17446 21699 17448
rect 8385 17443 8451 17446
rect 14917 17443 14983 17446
rect 21633 17443 21699 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 18137 17370 18203 17373
rect 25313 17370 25379 17373
rect 18137 17368 25379 17370
rect 18137 17312 18142 17368
rect 18198 17312 25318 17368
rect 25374 17312 25379 17368
rect 18137 17310 25379 17312
rect 18137 17307 18203 17310
rect 25313 17307 25379 17310
rect 7741 17234 7807 17237
rect 25037 17234 25103 17237
rect 7741 17232 25103 17234
rect 7741 17176 7746 17232
rect 7802 17176 25042 17232
rect 25098 17176 25103 17232
rect 7741 17174 25103 17176
rect 7741 17171 7807 17174
rect 25037 17171 25103 17174
rect 0 17098 480 17128
rect 3785 17098 3851 17101
rect 17309 17098 17375 17101
rect 21265 17098 21331 17101
rect 29520 17098 30000 17128
rect 0 17096 3851 17098
rect 0 17040 3790 17096
rect 3846 17040 3851 17096
rect 0 17038 3851 17040
rect 0 17008 480 17038
rect 3785 17035 3851 17038
rect 9998 17096 17375 17098
rect 9998 17040 17314 17096
rect 17370 17040 17375 17096
rect 9998 17038 17375 17040
rect 3877 16962 3943 16965
rect 9857 16962 9923 16965
rect 9998 16962 10058 17038
rect 17309 17035 17375 17038
rect 17542 17096 21331 17098
rect 17542 17040 21270 17096
rect 21326 17040 21331 17096
rect 17542 17038 21331 17040
rect 3877 16960 10058 16962
rect 3877 16904 3882 16960
rect 3938 16904 9862 16960
rect 9918 16904 10058 16960
rect 3877 16902 10058 16904
rect 12893 16962 12959 16965
rect 17542 16962 17602 17038
rect 21265 17035 21331 17038
rect 25822 17038 30000 17098
rect 12893 16960 17602 16962
rect 12893 16904 12898 16960
rect 12954 16904 17602 16960
rect 12893 16902 17602 16904
rect 3877 16899 3943 16902
rect 9857 16899 9923 16902
rect 12893 16899 12959 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 1761 16826 1827 16829
rect 4429 16826 4495 16829
rect 1761 16824 4495 16826
rect 1761 16768 1766 16824
rect 1822 16768 4434 16824
rect 4490 16768 4495 16824
rect 1761 16766 4495 16768
rect 1761 16763 1827 16766
rect 4429 16763 4495 16766
rect 2773 16690 2839 16693
rect 7741 16690 7807 16693
rect 2773 16688 7807 16690
rect 2773 16632 2778 16688
rect 2834 16632 7746 16688
rect 7802 16632 7807 16688
rect 2773 16630 7807 16632
rect 2773 16627 2839 16630
rect 7741 16627 7807 16630
rect 8293 16692 8359 16693
rect 8293 16688 8340 16692
rect 8404 16690 8410 16692
rect 12157 16690 12223 16693
rect 15285 16690 15351 16693
rect 8293 16632 8298 16688
rect 8293 16628 8340 16632
rect 8404 16630 8450 16690
rect 12157 16688 15351 16690
rect 12157 16632 12162 16688
rect 12218 16632 15290 16688
rect 15346 16632 15351 16688
rect 12157 16630 15351 16632
rect 8404 16628 8410 16630
rect 8293 16627 8359 16628
rect 12157 16627 12223 16630
rect 15285 16627 15351 16630
rect 11605 16554 11671 16557
rect 17125 16554 17191 16557
rect 11605 16552 17191 16554
rect 11605 16496 11610 16552
rect 11666 16496 17130 16552
rect 17186 16496 17191 16552
rect 11605 16494 17191 16496
rect 11605 16491 11671 16494
rect 17125 16491 17191 16494
rect 17493 16554 17559 16557
rect 25822 16554 25882 17038
rect 29520 17008 30000 17038
rect 26417 16690 26483 16693
rect 26550 16690 26556 16692
rect 26417 16688 26556 16690
rect 26417 16632 26422 16688
rect 26478 16632 26556 16688
rect 26417 16630 26556 16632
rect 26417 16627 26483 16630
rect 26550 16628 26556 16630
rect 26620 16628 26626 16692
rect 17493 16552 25882 16554
rect 17493 16496 17498 16552
rect 17554 16496 25882 16552
rect 17493 16494 25882 16496
rect 17493 16491 17559 16494
rect 0 16418 480 16448
rect 5073 16418 5139 16421
rect 0 16416 5139 16418
rect 0 16360 5078 16416
rect 5134 16360 5139 16416
rect 0 16358 5139 16360
rect 0 16328 480 16358
rect 5073 16355 5139 16358
rect 15009 16418 15075 16421
rect 15653 16418 15719 16421
rect 15009 16416 15719 16418
rect 15009 16360 15014 16416
rect 15070 16360 15658 16416
rect 15714 16360 15719 16416
rect 15009 16358 15719 16360
rect 15009 16355 15075 16358
rect 15653 16355 15719 16358
rect 17309 16418 17375 16421
rect 24945 16418 25011 16421
rect 26877 16418 26943 16421
rect 29520 16418 30000 16448
rect 17309 16416 25882 16418
rect 17309 16360 17314 16416
rect 17370 16360 24950 16416
rect 25006 16360 25882 16416
rect 17309 16358 25882 16360
rect 17309 16355 17375 16358
rect 24945 16355 25011 16358
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 16389 16282 16455 16285
rect 17493 16282 17559 16285
rect 16389 16280 17559 16282
rect 16389 16224 16394 16280
rect 16450 16224 17498 16280
rect 17554 16224 17559 16280
rect 16389 16222 17559 16224
rect 16389 16219 16455 16222
rect 17493 16219 17559 16222
rect 3785 16146 3851 16149
rect 8937 16146 9003 16149
rect 14641 16146 14707 16149
rect 3785 16144 14707 16146
rect 3785 16088 3790 16144
rect 3846 16088 8942 16144
rect 8998 16088 14646 16144
rect 14702 16088 14707 16144
rect 3785 16086 14707 16088
rect 3785 16083 3851 16086
rect 8937 16083 9003 16086
rect 14641 16083 14707 16086
rect 21817 16146 21883 16149
rect 25497 16146 25563 16149
rect 21817 16144 25563 16146
rect 21817 16088 21822 16144
rect 21878 16088 25502 16144
rect 25558 16088 25563 16144
rect 21817 16086 25563 16088
rect 25822 16146 25882 16358
rect 26877 16416 30000 16418
rect 26877 16360 26882 16416
rect 26938 16360 30000 16416
rect 26877 16358 30000 16360
rect 26877 16355 26943 16358
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 29520 16328 30000 16358
rect 25944 16287 26264 16288
rect 26785 16146 26851 16149
rect 25822 16144 26851 16146
rect 25822 16088 26790 16144
rect 26846 16088 26851 16144
rect 25822 16086 26851 16088
rect 21817 16083 21883 16086
rect 25497 16083 25563 16086
rect 26785 16083 26851 16086
rect 2589 16010 2655 16013
rect 18597 16010 18663 16013
rect 2454 16008 18663 16010
rect 2454 15952 2594 16008
rect 2650 15952 18602 16008
rect 18658 15952 18663 16008
rect 2454 15950 18663 15952
rect 0 15874 480 15904
rect 2454 15874 2514 15950
rect 2589 15947 2655 15950
rect 18597 15947 18663 15950
rect 0 15814 2514 15874
rect 3325 15874 3391 15877
rect 6545 15874 6611 15877
rect 3325 15872 6611 15874
rect 3325 15816 3330 15872
rect 3386 15816 6550 15872
rect 6606 15816 6611 15872
rect 3325 15814 6611 15816
rect 0 15784 480 15814
rect 3325 15811 3391 15814
rect 6545 15811 6611 15814
rect 25129 15874 25195 15877
rect 29520 15874 30000 15904
rect 25129 15872 30000 15874
rect 25129 15816 25134 15872
rect 25190 15816 30000 15872
rect 25129 15814 30000 15816
rect 25129 15811 25195 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 14917 15738 14983 15741
rect 18505 15738 18571 15741
rect 14917 15736 18571 15738
rect 14917 15680 14922 15736
rect 14978 15680 18510 15736
rect 18566 15680 18571 15736
rect 14917 15678 18571 15680
rect 14917 15675 14983 15678
rect 18505 15675 18571 15678
rect 4429 15602 4495 15605
rect 5625 15602 5691 15605
rect 11421 15602 11487 15605
rect 12157 15602 12223 15605
rect 4429 15600 12223 15602
rect 4429 15544 4434 15600
rect 4490 15544 5630 15600
rect 5686 15544 11426 15600
rect 11482 15544 12162 15600
rect 12218 15544 12223 15600
rect 4429 15542 12223 15544
rect 4429 15539 4495 15542
rect 5625 15539 5691 15542
rect 11421 15539 11487 15542
rect 12157 15539 12223 15542
rect 13813 15602 13879 15605
rect 13813 15600 26434 15602
rect 13813 15544 13818 15600
rect 13874 15544 26434 15600
rect 13813 15542 26434 15544
rect 13813 15539 13879 15542
rect 7189 15466 7255 15469
rect 12617 15466 12683 15469
rect 15009 15466 15075 15469
rect 18229 15466 18295 15469
rect 7189 15464 18295 15466
rect 7189 15408 7194 15464
rect 7250 15408 12622 15464
rect 12678 15408 15014 15464
rect 15070 15408 18234 15464
rect 18290 15408 18295 15464
rect 7189 15406 18295 15408
rect 7189 15403 7255 15406
rect 12617 15403 12683 15406
rect 15009 15403 15075 15406
rect 18229 15403 18295 15406
rect 18505 15466 18571 15469
rect 23749 15466 23815 15469
rect 25313 15466 25379 15469
rect 26233 15466 26299 15469
rect 18505 15464 26299 15466
rect 18505 15408 18510 15464
rect 18566 15408 23754 15464
rect 23810 15408 25318 15464
rect 25374 15408 26238 15464
rect 26294 15408 26299 15464
rect 18505 15406 26299 15408
rect 18505 15403 18571 15406
rect 23749 15403 23815 15406
rect 25313 15403 25379 15406
rect 26233 15403 26299 15406
rect 0 15330 480 15360
rect 1117 15330 1183 15333
rect 0 15328 1183 15330
rect 0 15272 1122 15328
rect 1178 15272 1183 15328
rect 0 15270 1183 15272
rect 0 15240 480 15270
rect 1117 15267 1183 15270
rect 8017 15330 8083 15333
rect 12249 15330 12315 15333
rect 8017 15328 12315 15330
rect 8017 15272 8022 15328
rect 8078 15272 12254 15328
rect 12310 15272 12315 15328
rect 8017 15270 12315 15272
rect 26374 15330 26434 15542
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 8017 15267 8083 15270
rect 12249 15267 12315 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 8385 15194 8451 15197
rect 13169 15194 13235 15197
rect 8385 15192 13235 15194
rect 8385 15136 8390 15192
rect 8446 15136 13174 15192
rect 13230 15136 13235 15192
rect 8385 15134 13235 15136
rect 8385 15131 8451 15134
rect 13169 15131 13235 15134
rect 5809 15058 5875 15061
rect 18505 15058 18571 15061
rect 5809 15056 18571 15058
rect 5809 15000 5814 15056
rect 5870 15000 18510 15056
rect 18566 15000 18571 15056
rect 5809 14998 18571 15000
rect 5809 14995 5875 14998
rect 18505 14995 18571 14998
rect 19057 15058 19123 15061
rect 21449 15058 21515 15061
rect 19057 15056 21515 15058
rect 19057 15000 19062 15056
rect 19118 15000 21454 15056
rect 21510 15000 21515 15056
rect 19057 14998 21515 15000
rect 19057 14995 19123 14998
rect 21449 14995 21515 14998
rect 9489 14922 9555 14925
rect 12525 14922 12591 14925
rect 9489 14920 12591 14922
rect 9489 14864 9494 14920
rect 9550 14864 12530 14920
rect 12586 14864 12591 14920
rect 9489 14862 12591 14864
rect 9489 14859 9555 14862
rect 12525 14859 12591 14862
rect 13905 14922 13971 14925
rect 19609 14922 19675 14925
rect 13905 14920 19675 14922
rect 13905 14864 13910 14920
rect 13966 14864 19614 14920
rect 19670 14864 19675 14920
rect 13905 14862 19675 14864
rect 13905 14859 13971 14862
rect 19609 14859 19675 14862
rect 4337 14786 4403 14789
rect 9397 14786 9463 14789
rect 4337 14784 9463 14786
rect 4337 14728 4342 14784
rect 4398 14728 9402 14784
rect 9458 14728 9463 14784
rect 4337 14726 9463 14728
rect 4337 14723 4403 14726
rect 9397 14723 9463 14726
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 16389 14650 16455 14653
rect 20437 14650 20503 14653
rect 0 14590 2698 14650
rect 0 14560 480 14590
rect 2638 14514 2698 14590
rect 16389 14648 20503 14650
rect 16389 14592 16394 14648
rect 16450 14592 20442 14648
rect 20498 14592 20503 14648
rect 16389 14590 20503 14592
rect 16389 14587 16455 14590
rect 20437 14587 20503 14590
rect 25037 14650 25103 14653
rect 29520 14650 30000 14680
rect 25037 14648 30000 14650
rect 25037 14592 25042 14648
rect 25098 14592 30000 14648
rect 25037 14590 30000 14592
rect 25037 14587 25103 14590
rect 29520 14560 30000 14590
rect 3509 14514 3575 14517
rect 2638 14512 3575 14514
rect 2638 14456 3514 14512
rect 3570 14456 3575 14512
rect 2638 14454 3575 14456
rect 3509 14451 3575 14454
rect 9857 14514 9923 14517
rect 13169 14514 13235 14517
rect 9857 14512 13235 14514
rect 9857 14456 9862 14512
rect 9918 14456 13174 14512
rect 13230 14456 13235 14512
rect 9857 14454 13235 14456
rect 9857 14451 9923 14454
rect 13169 14451 13235 14454
rect 16481 14514 16547 14517
rect 23657 14514 23723 14517
rect 16481 14512 23723 14514
rect 16481 14456 16486 14512
rect 16542 14456 23662 14512
rect 23718 14456 23723 14512
rect 16481 14454 23723 14456
rect 16481 14451 16547 14454
rect 23657 14451 23723 14454
rect 4153 14378 4219 14381
rect 9029 14378 9095 14381
rect 4153 14376 9095 14378
rect 4153 14320 4158 14376
rect 4214 14320 9034 14376
rect 9090 14320 9095 14376
rect 4153 14318 9095 14320
rect 4153 14315 4219 14318
rect 9029 14315 9095 14318
rect 9305 14378 9371 14381
rect 14733 14378 14799 14381
rect 9305 14376 14799 14378
rect 9305 14320 9310 14376
rect 9366 14320 14738 14376
rect 14794 14320 14799 14376
rect 9305 14318 14799 14320
rect 9305 14315 9371 14318
rect 14733 14315 14799 14318
rect 24669 14378 24735 14381
rect 26601 14378 26667 14381
rect 24669 14376 26667 14378
rect 24669 14320 24674 14376
rect 24730 14320 26606 14376
rect 26662 14320 26667 14376
rect 24669 14318 26667 14320
rect 24669 14315 24735 14318
rect 26601 14315 26667 14318
rect 3877 14242 3943 14245
rect 5717 14242 5783 14245
rect 3877 14240 5783 14242
rect 3877 14184 3882 14240
rect 3938 14184 5722 14240
rect 5778 14184 5783 14240
rect 3877 14182 5783 14184
rect 3877 14179 3943 14182
rect 5717 14179 5783 14182
rect 7281 14242 7347 14245
rect 12065 14242 12131 14245
rect 7281 14240 12131 14242
rect 7281 14184 7286 14240
rect 7342 14184 12070 14240
rect 12126 14184 12131 14240
rect 7281 14182 12131 14184
rect 7281 14179 7347 14182
rect 12065 14179 12131 14182
rect 18597 14242 18663 14245
rect 24025 14242 24091 14245
rect 18597 14240 24091 14242
rect 18597 14184 18602 14240
rect 18658 14184 24030 14240
rect 24086 14184 24091 14240
rect 18597 14182 24091 14184
rect 18597 14179 18663 14182
rect 24025 14179 24091 14182
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 2221 14106 2287 14109
rect 3325 14106 3391 14109
rect 0 14104 3391 14106
rect 0 14048 2226 14104
rect 2282 14048 3330 14104
rect 3386 14048 3391 14104
rect 0 14046 3391 14048
rect 0 14016 480 14046
rect 2221 14043 2287 14046
rect 3325 14043 3391 14046
rect 19241 14106 19307 14109
rect 25129 14106 25195 14109
rect 19241 14104 25195 14106
rect 19241 14048 19246 14104
rect 19302 14048 25134 14104
rect 25190 14048 25195 14104
rect 19241 14046 25195 14048
rect 19241 14043 19307 14046
rect 25129 14043 25195 14046
rect 27337 14106 27403 14109
rect 29520 14106 30000 14136
rect 27337 14104 30000 14106
rect 27337 14048 27342 14104
rect 27398 14048 30000 14104
rect 27337 14046 30000 14048
rect 27337 14043 27403 14046
rect 2865 13970 2931 13973
rect 16481 13970 16547 13973
rect 2865 13968 16547 13970
rect 2865 13912 2870 13968
rect 2926 13912 16486 13968
rect 16542 13912 16547 13968
rect 2865 13910 16547 13912
rect 2865 13907 2931 13910
rect 16481 13907 16547 13910
rect 25681 13970 25747 13973
rect 27340 13970 27400 14043
rect 29520 14016 30000 14046
rect 25681 13968 27400 13970
rect 25681 13912 25686 13968
rect 25742 13912 27400 13968
rect 25681 13910 27400 13912
rect 25681 13907 25747 13910
rect 10133 13834 10199 13837
rect 12433 13834 12499 13837
rect 10133 13832 12499 13834
rect 10133 13776 10138 13832
rect 10194 13776 12438 13832
rect 12494 13776 12499 13832
rect 10133 13774 12499 13776
rect 10133 13771 10199 13774
rect 12433 13771 12499 13774
rect 15469 13834 15535 13837
rect 19609 13834 19675 13837
rect 15469 13832 19675 13834
rect 15469 13776 15474 13832
rect 15530 13776 19614 13832
rect 19670 13776 19675 13832
rect 15469 13774 19675 13776
rect 15469 13771 15535 13774
rect 19609 13771 19675 13774
rect 19885 13834 19951 13837
rect 23933 13834 23999 13837
rect 27521 13834 27587 13837
rect 19885 13832 27587 13834
rect 19885 13776 19890 13832
rect 19946 13776 23938 13832
rect 23994 13776 27526 13832
rect 27582 13776 27587 13832
rect 19885 13774 27587 13776
rect 19885 13771 19951 13774
rect 23933 13771 23999 13774
rect 27521 13771 27587 13774
rect 2589 13698 2655 13701
rect 6177 13698 6243 13701
rect 2589 13696 6243 13698
rect 2589 13640 2594 13696
rect 2650 13640 6182 13696
rect 6238 13640 6243 13696
rect 2589 13638 6243 13640
rect 2589 13635 2655 13638
rect 6177 13635 6243 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 2037 13562 2103 13565
rect 5625 13562 5691 13565
rect 2037 13560 5691 13562
rect 2037 13504 2042 13560
rect 2098 13504 5630 13560
rect 5686 13504 5691 13560
rect 2037 13502 5691 13504
rect 2037 13499 2103 13502
rect 5625 13499 5691 13502
rect 5809 13562 5875 13565
rect 7557 13562 7623 13565
rect 5809 13560 7623 13562
rect 5809 13504 5814 13560
rect 5870 13504 7562 13560
rect 7618 13504 7623 13560
rect 5809 13502 7623 13504
rect 5809 13499 5875 13502
rect 7557 13499 7623 13502
rect 12157 13562 12223 13565
rect 12801 13562 12867 13565
rect 12157 13560 12867 13562
rect 12157 13504 12162 13560
rect 12218 13504 12806 13560
rect 12862 13504 12867 13560
rect 12157 13502 12867 13504
rect 12157 13499 12223 13502
rect 12801 13499 12867 13502
rect 18873 13562 18939 13565
rect 18873 13560 20546 13562
rect 18873 13504 18878 13560
rect 18934 13504 20546 13560
rect 18873 13502 20546 13504
rect 18873 13499 18939 13502
rect 0 13426 480 13456
rect 1577 13426 1643 13429
rect 7649 13426 7715 13429
rect 14917 13426 14983 13429
rect 20345 13426 20411 13429
rect 0 13424 1962 13426
rect 0 13368 1582 13424
rect 1638 13368 1962 13424
rect 0 13366 1962 13368
rect 0 13336 480 13366
rect 1577 13363 1643 13366
rect 1902 13154 1962 13366
rect 7649 13424 20411 13426
rect 7649 13368 7654 13424
rect 7710 13368 14922 13424
rect 14978 13368 20350 13424
rect 20406 13368 20411 13424
rect 7649 13366 20411 13368
rect 20486 13426 20546 13502
rect 22185 13426 22251 13429
rect 27797 13426 27863 13429
rect 29520 13426 30000 13456
rect 20486 13424 30000 13426
rect 20486 13368 22190 13424
rect 22246 13368 27802 13424
rect 27858 13368 30000 13424
rect 20486 13366 30000 13368
rect 7649 13363 7715 13366
rect 14917 13363 14983 13366
rect 20345 13363 20411 13366
rect 22185 13363 22251 13366
rect 27797 13363 27863 13366
rect 29520 13336 30000 13366
rect 5257 13290 5323 13293
rect 8293 13290 8359 13293
rect 18873 13290 18939 13293
rect 5257 13288 8359 13290
rect 5257 13232 5262 13288
rect 5318 13232 8298 13288
rect 8354 13232 8359 13288
rect 5257 13230 8359 13232
rect 5257 13227 5323 13230
rect 8293 13227 8359 13230
rect 15702 13288 18939 13290
rect 15702 13232 18878 13288
rect 18934 13232 18939 13288
rect 15702 13230 18939 13232
rect 5809 13154 5875 13157
rect 1902 13152 5875 13154
rect 1902 13096 5814 13152
rect 5870 13096 5875 13152
rect 1902 13094 5875 13096
rect 5809 13091 5875 13094
rect 6361 13154 6427 13157
rect 7741 13154 7807 13157
rect 12893 13154 12959 13157
rect 15702 13154 15762 13230
rect 18873 13227 18939 13230
rect 6361 13152 15762 13154
rect 6361 13096 6366 13152
rect 6422 13096 7746 13152
rect 7802 13096 12898 13152
rect 12954 13096 15762 13152
rect 6361 13094 15762 13096
rect 16481 13154 16547 13157
rect 23473 13154 23539 13157
rect 24301 13154 24367 13157
rect 16481 13152 24367 13154
rect 16481 13096 16486 13152
rect 16542 13096 23478 13152
rect 23534 13096 24306 13152
rect 24362 13096 24367 13152
rect 16481 13094 24367 13096
rect 6361 13091 6427 13094
rect 7741 13091 7807 13094
rect 12893 13091 12959 13094
rect 16481 13091 16547 13094
rect 23473 13091 23539 13094
rect 24301 13091 24367 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 18689 13018 18755 13021
rect 21817 13018 21883 13021
rect 18689 13016 21883 13018
rect 18689 12960 18694 13016
rect 18750 12960 21822 13016
rect 21878 12960 21883 13016
rect 18689 12958 21883 12960
rect 18689 12955 18755 12958
rect 21817 12955 21883 12958
rect 0 12882 480 12912
rect 6269 12882 6335 12885
rect 11789 12882 11855 12885
rect 0 12822 2146 12882
rect 0 12792 480 12822
rect 2086 12613 2146 12822
rect 6269 12880 11855 12882
rect 6269 12824 6274 12880
rect 6330 12824 11794 12880
rect 11850 12824 11855 12880
rect 6269 12822 11855 12824
rect 6269 12819 6335 12822
rect 11789 12819 11855 12822
rect 12801 12882 12867 12885
rect 19333 12882 19399 12885
rect 12801 12880 19399 12882
rect 12801 12824 12806 12880
rect 12862 12824 19338 12880
rect 19394 12824 19399 12880
rect 12801 12822 19399 12824
rect 12801 12819 12867 12822
rect 19333 12819 19399 12822
rect 26877 12882 26943 12885
rect 29520 12882 30000 12912
rect 26877 12880 30000 12882
rect 26877 12824 26882 12880
rect 26938 12824 30000 12880
rect 26877 12822 30000 12824
rect 26877 12819 26943 12822
rect 29520 12792 30000 12822
rect 5625 12746 5691 12749
rect 18689 12746 18755 12749
rect 5625 12744 18755 12746
rect 5625 12688 5630 12744
rect 5686 12688 18694 12744
rect 18750 12688 18755 12744
rect 5625 12686 18755 12688
rect 5625 12683 5691 12686
rect 18689 12683 18755 12686
rect 19057 12746 19123 12749
rect 25497 12746 25563 12749
rect 19057 12744 25563 12746
rect 19057 12688 19062 12744
rect 19118 12688 25502 12744
rect 25558 12688 25563 12744
rect 19057 12686 25563 12688
rect 19057 12683 19123 12686
rect 25497 12683 25563 12686
rect 2086 12610 2195 12613
rect 4245 12610 4311 12613
rect 10777 12610 10843 12613
rect 2086 12608 10843 12610
rect 2086 12552 2134 12608
rect 2190 12552 4250 12608
rect 4306 12552 10782 12608
rect 10838 12552 10843 12608
rect 2086 12550 10843 12552
rect 2129 12547 2195 12550
rect 4245 12547 4311 12550
rect 10777 12547 10843 12550
rect 11605 12610 11671 12613
rect 15561 12610 15627 12613
rect 11605 12608 15627 12610
rect 11605 12552 11610 12608
rect 11666 12552 15566 12608
rect 15622 12552 15627 12608
rect 11605 12550 15627 12552
rect 11605 12547 11671 12550
rect 15561 12547 15627 12550
rect 22461 12610 22527 12613
rect 27061 12610 27127 12613
rect 22461 12608 27127 12610
rect 22461 12552 22466 12608
rect 22522 12552 27066 12608
rect 27122 12552 27127 12608
rect 22461 12550 27127 12552
rect 22461 12547 22527 12550
rect 27061 12547 27127 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 21725 12474 21791 12477
rect 24117 12474 24183 12477
rect 21725 12472 25146 12474
rect 21725 12416 21730 12472
rect 21786 12416 24122 12472
rect 24178 12416 25146 12472
rect 21725 12414 25146 12416
rect 21725 12411 21791 12414
rect 24117 12411 24183 12414
rect 0 12338 480 12368
rect 1209 12338 1275 12341
rect 0 12336 1275 12338
rect 0 12280 1214 12336
rect 1270 12280 1275 12336
rect 0 12278 1275 12280
rect 0 12248 480 12278
rect 1209 12275 1275 12278
rect 2865 12338 2931 12341
rect 4429 12338 4495 12341
rect 2865 12336 4495 12338
rect 2865 12280 2870 12336
rect 2926 12280 4434 12336
rect 4490 12280 4495 12336
rect 2865 12278 4495 12280
rect 2865 12275 2931 12278
rect 4429 12275 4495 12278
rect 21541 12338 21607 12341
rect 24117 12338 24183 12341
rect 21541 12336 24183 12338
rect 21541 12280 21546 12336
rect 21602 12280 24122 12336
rect 24178 12280 24183 12336
rect 21541 12278 24183 12280
rect 21541 12275 21607 12278
rect 24117 12275 24183 12278
rect 24761 12338 24827 12341
rect 24945 12338 25011 12341
rect 24761 12336 25011 12338
rect 24761 12280 24766 12336
rect 24822 12280 24950 12336
rect 25006 12280 25011 12336
rect 24761 12278 25011 12280
rect 25086 12338 25146 12414
rect 29520 12338 30000 12368
rect 25086 12278 30000 12338
rect 24761 12275 24827 12278
rect 24945 12275 25011 12278
rect 29520 12248 30000 12278
rect 4521 12202 4587 12205
rect 10777 12202 10843 12205
rect 4521 12200 10843 12202
rect 4521 12144 4526 12200
rect 4582 12144 10782 12200
rect 10838 12144 10843 12200
rect 4521 12142 10843 12144
rect 4521 12139 4587 12142
rect 10777 12139 10843 12142
rect 19333 12202 19399 12205
rect 26693 12202 26759 12205
rect 27337 12202 27403 12205
rect 19333 12200 27403 12202
rect 19333 12144 19338 12200
rect 19394 12144 26698 12200
rect 26754 12144 27342 12200
rect 27398 12144 27403 12200
rect 19333 12142 27403 12144
rect 19333 12139 19399 12142
rect 26693 12139 26759 12142
rect 27337 12139 27403 12142
rect 18505 12066 18571 12069
rect 19609 12066 19675 12069
rect 24761 12066 24827 12069
rect 25405 12066 25471 12069
rect 18505 12064 25471 12066
rect 18505 12008 18510 12064
rect 18566 12008 19614 12064
rect 19670 12008 24766 12064
rect 24822 12008 25410 12064
rect 25466 12008 25471 12064
rect 18505 12006 25471 12008
rect 18505 12003 18571 12006
rect 19609 12003 19675 12006
rect 24761 12003 24827 12006
rect 25405 12003 25471 12006
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 0 11658 480 11688
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11568 480 11598
rect 4061 11595 4127 11598
rect 21357 11658 21423 11661
rect 29520 11658 30000 11688
rect 21357 11656 30000 11658
rect 21357 11600 21362 11656
rect 21418 11600 30000 11656
rect 21357 11598 30000 11600
rect 21357 11595 21423 11598
rect 29520 11568 30000 11598
rect 7097 11522 7163 11525
rect 10133 11522 10199 11525
rect 7097 11520 10199 11522
rect 7097 11464 7102 11520
rect 7158 11464 10138 11520
rect 10194 11464 10199 11520
rect 7097 11462 10199 11464
rect 7097 11459 7163 11462
rect 10133 11459 10199 11462
rect 19241 11522 19307 11525
rect 20805 11522 20871 11525
rect 19241 11520 20871 11522
rect 19241 11464 19246 11520
rect 19302 11464 20810 11520
rect 20866 11464 20871 11520
rect 19241 11462 20871 11464
rect 19241 11459 19307 11462
rect 20805 11459 20871 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 5165 11386 5231 11389
rect 6913 11386 6979 11389
rect 5165 11384 6979 11386
rect 5165 11328 5170 11384
rect 5226 11328 6918 11384
rect 6974 11328 6979 11384
rect 5165 11326 6979 11328
rect 5165 11323 5231 11326
rect 6913 11323 6979 11326
rect 15285 11386 15351 11389
rect 19701 11386 19767 11389
rect 25773 11386 25839 11389
rect 26877 11386 26943 11389
rect 15285 11384 19767 11386
rect 15285 11328 15290 11384
rect 15346 11328 19706 11384
rect 19762 11328 19767 11384
rect 15285 11326 19767 11328
rect 15285 11323 15351 11326
rect 19701 11323 19767 11326
rect 21406 11384 26943 11386
rect 21406 11328 25778 11384
rect 25834 11328 26882 11384
rect 26938 11328 26943 11384
rect 21406 11326 26943 11328
rect 2589 11250 2655 11253
rect 13077 11250 13143 11253
rect 2589 11248 13143 11250
rect 2589 11192 2594 11248
rect 2650 11192 13082 11248
rect 13138 11192 13143 11248
rect 2589 11190 13143 11192
rect 2589 11187 2655 11190
rect 13077 11187 13143 11190
rect 13302 11188 13308 11252
rect 13372 11250 13378 11252
rect 13445 11250 13511 11253
rect 13372 11248 13511 11250
rect 13372 11192 13450 11248
rect 13506 11192 13511 11248
rect 13372 11190 13511 11192
rect 13372 11188 13378 11190
rect 13445 11187 13511 11190
rect 18781 11250 18847 11253
rect 19885 11250 19951 11253
rect 21406 11250 21466 11326
rect 25773 11323 25839 11326
rect 26877 11323 26943 11326
rect 18781 11248 21466 11250
rect 18781 11192 18786 11248
rect 18842 11192 19890 11248
rect 19946 11192 21466 11248
rect 18781 11190 21466 11192
rect 18781 11187 18847 11190
rect 19885 11187 19951 11190
rect 0 11114 480 11144
rect 4245 11114 4311 11117
rect 0 11112 4311 11114
rect 0 11056 4250 11112
rect 4306 11056 4311 11112
rect 0 11054 4311 11056
rect 0 11024 480 11054
rect 4245 11051 4311 11054
rect 14825 11114 14891 11117
rect 18321 11114 18387 11117
rect 14825 11112 18387 11114
rect 14825 11056 14830 11112
rect 14886 11056 18326 11112
rect 18382 11056 18387 11112
rect 14825 11054 18387 11056
rect 14825 11051 14891 11054
rect 18321 11051 18387 11054
rect 23749 11114 23815 11117
rect 29520 11114 30000 11144
rect 23749 11112 30000 11114
rect 23749 11056 23754 11112
rect 23810 11056 30000 11112
rect 23749 11054 30000 11056
rect 23749 11051 23815 11054
rect 29520 11024 30000 11054
rect 9213 10978 9279 10981
rect 12249 10978 12315 10981
rect 9213 10976 12315 10978
rect 9213 10920 9218 10976
rect 9274 10920 12254 10976
rect 12310 10920 12315 10976
rect 9213 10918 12315 10920
rect 9213 10915 9279 10918
rect 12249 10915 12315 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 2865 10842 2931 10845
rect 2998 10842 3004 10844
rect 2865 10840 3004 10842
rect 2865 10784 2870 10840
rect 2926 10784 3004 10840
rect 2865 10782 3004 10784
rect 2865 10779 2931 10782
rect 2998 10780 3004 10782
rect 3068 10780 3074 10844
rect 9765 10842 9831 10845
rect 20345 10842 20411 10845
rect 22001 10842 22067 10845
rect 7238 10840 9874 10842
rect 7238 10784 9770 10840
rect 9826 10784 9874 10840
rect 7238 10782 9874 10784
rect 7238 10706 7298 10782
rect 9765 10779 9874 10782
rect 20345 10840 22067 10842
rect 20345 10784 20350 10840
rect 20406 10784 22006 10840
rect 22062 10784 22067 10840
rect 20345 10782 22067 10784
rect 20345 10779 20411 10782
rect 22001 10779 22067 10782
rect 3558 10646 7298 10706
rect 7465 10706 7531 10709
rect 9673 10706 9739 10709
rect 7465 10704 9739 10706
rect 7465 10648 7470 10704
rect 7526 10648 9678 10704
rect 9734 10648 9739 10704
rect 7465 10646 9739 10648
rect 9814 10706 9874 10779
rect 25957 10706 26023 10709
rect 9814 10704 26023 10706
rect 9814 10648 25962 10704
rect 26018 10648 26023 10704
rect 9814 10646 26023 10648
rect 2129 10570 2195 10573
rect 3558 10570 3618 10646
rect 7465 10643 7531 10646
rect 9673 10643 9739 10646
rect 25957 10643 26023 10646
rect 2129 10568 3618 10570
rect 2129 10512 2134 10568
rect 2190 10512 3618 10568
rect 2129 10510 3618 10512
rect 3693 10570 3759 10573
rect 13537 10570 13603 10573
rect 3693 10568 13603 10570
rect 3693 10512 3698 10568
rect 3754 10512 13542 10568
rect 13598 10512 13603 10568
rect 3693 10510 13603 10512
rect 2129 10507 2195 10510
rect 3693 10507 3759 10510
rect 13537 10507 13603 10510
rect 15745 10570 15811 10573
rect 19977 10570 20043 10573
rect 15745 10568 20043 10570
rect 15745 10512 15750 10568
rect 15806 10512 19982 10568
rect 20038 10512 20043 10568
rect 15745 10510 20043 10512
rect 15745 10507 15811 10510
rect 19977 10507 20043 10510
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 25129 10434 25195 10437
rect 29520 10434 30000 10464
rect 25129 10432 30000 10434
rect 25129 10376 25134 10432
rect 25190 10376 30000 10432
rect 25129 10374 30000 10376
rect 25129 10371 25195 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 1669 10298 1735 10301
rect 3325 10298 3391 10301
rect 1669 10296 3391 10298
rect 1669 10240 1674 10296
rect 1730 10240 3330 10296
rect 3386 10240 3391 10296
rect 1669 10238 3391 10240
rect 1669 10235 1735 10238
rect 3325 10235 3391 10238
rect 7833 10162 7899 10165
rect 17401 10162 17467 10165
rect 27521 10162 27587 10165
rect 7833 10160 17234 10162
rect 7833 10104 7838 10160
rect 7894 10104 17234 10160
rect 7833 10102 17234 10104
rect 7833 10099 7899 10102
rect 3509 10026 3575 10029
rect 7281 10026 7347 10029
rect 3509 10024 7347 10026
rect 3509 9968 3514 10024
rect 3570 9968 7286 10024
rect 7342 9968 7347 10024
rect 3509 9966 7347 9968
rect 3509 9963 3575 9966
rect 7281 9963 7347 9966
rect 7557 10026 7623 10029
rect 17033 10026 17099 10029
rect 7557 10024 17099 10026
rect 7557 9968 7562 10024
rect 7618 9968 17038 10024
rect 17094 9968 17099 10024
rect 7557 9966 17099 9968
rect 17174 10026 17234 10102
rect 17401 10160 27587 10162
rect 17401 10104 17406 10160
rect 17462 10104 27526 10160
rect 27582 10104 27587 10160
rect 17401 10102 27587 10104
rect 17401 10099 17467 10102
rect 27521 10099 27587 10102
rect 25037 10026 25103 10029
rect 17174 10024 25103 10026
rect 17174 9968 25042 10024
rect 25098 9968 25103 10024
rect 17174 9966 25103 9968
rect 7557 9963 7623 9966
rect 17033 9963 17099 9966
rect 25037 9963 25103 9966
rect 25589 10026 25655 10029
rect 25589 10024 26434 10026
rect 25589 9968 25594 10024
rect 25650 9968 26434 10024
rect 25589 9966 26434 9968
rect 25589 9963 25655 9966
rect 0 9890 480 9920
rect 5441 9890 5507 9893
rect 0 9888 5507 9890
rect 0 9832 5446 9888
rect 5502 9832 5507 9888
rect 0 9830 5507 9832
rect 26374 9890 26434 9966
rect 29520 9890 30000 9920
rect 26374 9830 30000 9890
rect 0 9800 480 9830
rect 5441 9827 5507 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 2589 9754 2655 9757
rect 3601 9754 3667 9757
rect 2589 9752 3667 9754
rect 2589 9696 2594 9752
rect 2650 9696 3606 9752
rect 3662 9696 3667 9752
rect 2589 9694 3667 9696
rect 2589 9691 2655 9694
rect 3601 9691 3667 9694
rect 8569 9618 8635 9621
rect 15377 9618 15443 9621
rect 8569 9616 15443 9618
rect 8569 9560 8574 9616
rect 8630 9560 15382 9616
rect 15438 9560 15443 9616
rect 8569 9558 15443 9560
rect 8569 9555 8635 9558
rect 15377 9555 15443 9558
rect 18413 9618 18479 9621
rect 25221 9618 25287 9621
rect 18413 9616 25287 9618
rect 18413 9560 18418 9616
rect 18474 9560 25226 9616
rect 25282 9560 25287 9616
rect 18413 9558 25287 9560
rect 18413 9555 18479 9558
rect 25221 9555 25287 9558
rect 25497 9618 25563 9621
rect 27429 9618 27495 9621
rect 25497 9616 27495 9618
rect 25497 9560 25502 9616
rect 25558 9560 27434 9616
rect 27490 9560 27495 9616
rect 25497 9558 27495 9560
rect 25497 9555 25563 9558
rect 27429 9555 27495 9558
rect 10685 9482 10751 9485
rect 21449 9482 21515 9485
rect 25313 9482 25379 9485
rect 10685 9480 25379 9482
rect 10685 9424 10690 9480
rect 10746 9424 21454 9480
rect 21510 9424 25318 9480
rect 25374 9424 25379 9480
rect 10685 9422 25379 9424
rect 10685 9419 10751 9422
rect 21449 9419 21515 9422
rect 25313 9419 25379 9422
rect 0 9346 480 9376
rect 4061 9346 4127 9349
rect 0 9344 4127 9346
rect 0 9288 4066 9344
rect 4122 9288 4127 9344
rect 0 9286 4127 9288
rect 0 9256 480 9286
rect 4061 9283 4127 9286
rect 25497 9346 25563 9349
rect 29520 9346 30000 9376
rect 25497 9344 30000 9346
rect 25497 9288 25502 9344
rect 25558 9288 30000 9344
rect 25497 9286 30000 9288
rect 25497 9283 25563 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 2773 9074 2839 9077
rect 8293 9074 8359 9077
rect 25681 9074 25747 9077
rect 27337 9074 27403 9077
rect 2773 9072 8359 9074
rect 2773 9016 2778 9072
rect 2834 9016 8298 9072
rect 8354 9016 8359 9072
rect 2773 9014 8359 9016
rect 2773 9011 2839 9014
rect 8293 9011 8359 9014
rect 8526 9072 27403 9074
rect 8526 9016 25686 9072
rect 25742 9016 27342 9072
rect 27398 9016 27403 9072
rect 8526 9014 27403 9016
rect 3785 8938 3851 8941
rect 8526 8938 8586 9014
rect 25681 9011 25747 9014
rect 27337 9011 27403 9014
rect 3785 8936 8586 8938
rect 3785 8880 3790 8936
rect 3846 8880 8586 8936
rect 3785 8878 8586 8880
rect 20161 8938 20227 8941
rect 26417 8938 26483 8941
rect 20161 8936 26483 8938
rect 20161 8880 20166 8936
rect 20222 8880 26422 8936
rect 26478 8880 26483 8936
rect 20161 8878 26483 8880
rect 3785 8875 3851 8878
rect 20161 8875 20227 8878
rect 26417 8875 26483 8878
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 4245 8666 4311 8669
rect 0 8664 4311 8666
rect 0 8608 4250 8664
rect 4306 8608 4311 8664
rect 0 8606 4311 8608
rect 0 8576 480 8606
rect 4245 8603 4311 8606
rect 27705 8666 27771 8669
rect 29520 8666 30000 8696
rect 27705 8664 30000 8666
rect 27705 8608 27710 8664
rect 27766 8608 30000 8664
rect 27705 8606 30000 8608
rect 27705 8603 27771 8606
rect 29520 8576 30000 8606
rect 13445 8530 13511 8533
rect 26509 8530 26575 8533
rect 13445 8528 26575 8530
rect 13445 8472 13450 8528
rect 13506 8472 26514 8528
rect 26570 8472 26575 8528
rect 13445 8470 26575 8472
rect 13445 8467 13511 8470
rect 26509 8467 26575 8470
rect 5441 8394 5507 8397
rect 7189 8394 7255 8397
rect 5441 8392 7255 8394
rect 5441 8336 5446 8392
rect 5502 8336 7194 8392
rect 7250 8336 7255 8392
rect 5441 8334 7255 8336
rect 5441 8331 5507 8334
rect 7189 8331 7255 8334
rect 26601 8394 26667 8397
rect 26601 8392 27538 8394
rect 26601 8336 26606 8392
rect 26662 8336 27538 8392
rect 26601 8334 27538 8336
rect 26601 8331 26667 8334
rect 25773 8258 25839 8261
rect 26693 8258 26759 8261
rect 25773 8256 26759 8258
rect 25773 8200 25778 8256
rect 25834 8200 26698 8256
rect 26754 8200 26759 8256
rect 25773 8198 26759 8200
rect 25773 8195 25839 8198
rect 26693 8195 26759 8198
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 2497 8122 2563 8125
rect 0 8120 2563 8122
rect 0 8064 2502 8120
rect 2558 8064 2563 8120
rect 0 8062 2563 8064
rect 27478 8122 27538 8334
rect 29520 8122 30000 8152
rect 27478 8062 30000 8122
rect 0 8032 480 8062
rect 2497 8059 2563 8062
rect 29520 8032 30000 8062
rect 22645 7986 22711 7989
rect 25313 7986 25379 7989
rect 22645 7984 25379 7986
rect 22645 7928 22650 7984
rect 22706 7928 25318 7984
rect 25374 7928 25379 7984
rect 22645 7926 25379 7928
rect 22645 7923 22711 7926
rect 25313 7923 25379 7926
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 24301 7442 24367 7445
rect 27521 7442 27587 7445
rect 24301 7440 27587 7442
rect 24301 7384 24306 7440
rect 24362 7384 27526 7440
rect 27582 7384 27587 7440
rect 24301 7382 27587 7384
rect 24301 7379 24367 7382
rect 27521 7379 27587 7382
rect 27705 7442 27771 7445
rect 29520 7442 30000 7472
rect 27705 7440 30000 7442
rect 27705 7384 27710 7440
rect 27766 7384 30000 7440
rect 27705 7382 30000 7384
rect 27705 7379 27771 7382
rect 29520 7352 30000 7382
rect 1761 7306 1827 7309
rect 11881 7306 11947 7309
rect 1761 7304 11947 7306
rect 1761 7248 1766 7304
rect 1822 7248 11886 7304
rect 11942 7248 11947 7304
rect 1761 7246 11947 7248
rect 1761 7243 1827 7246
rect 11881 7243 11947 7246
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 3141 6898 3207 6901
rect 5165 6898 5231 6901
rect 7189 6898 7255 6901
rect 3141 6896 7255 6898
rect 3141 6840 3146 6896
rect 3202 6840 5170 6896
rect 5226 6840 7194 6896
rect 7250 6840 7255 6896
rect 3141 6838 7255 6840
rect 3141 6835 3207 6838
rect 5165 6835 5231 6838
rect 7189 6835 7255 6838
rect 26601 6898 26667 6901
rect 29520 6898 30000 6928
rect 26601 6896 30000 6898
rect 26601 6840 26606 6896
rect 26662 6840 30000 6896
rect 26601 6838 30000 6840
rect 26601 6835 26667 6838
rect 29520 6808 30000 6838
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 2037 6490 2103 6493
rect 5349 6490 5415 6493
rect 2037 6488 5415 6490
rect 2037 6432 2042 6488
rect 2098 6432 5354 6488
rect 5410 6432 5415 6488
rect 2037 6430 5415 6432
rect 2037 6427 2103 6430
rect 5349 6427 5415 6430
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 26693 6354 26759 6357
rect 29520 6354 30000 6384
rect 26693 6352 30000 6354
rect 26693 6296 26698 6352
rect 26754 6296 30000 6352
rect 26693 6294 30000 6296
rect 26693 6291 26759 6294
rect 29520 6264 30000 6294
rect 3509 6218 3575 6221
rect 18229 6218 18295 6221
rect 3509 6216 18295 6218
rect 3509 6160 3514 6216
rect 3570 6160 18234 6216
rect 18290 6160 18295 6216
rect 3509 6158 18295 6160
rect 3509 6155 3575 6158
rect 18229 6155 18295 6158
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 2497 5810 2563 5813
rect 5809 5810 5875 5813
rect 2497 5808 5875 5810
rect 2497 5752 2502 5808
rect 2558 5752 5814 5808
rect 5870 5752 5875 5808
rect 2497 5750 5875 5752
rect 2497 5747 2563 5750
rect 5809 5747 5875 5750
rect 17309 5810 17375 5813
rect 26509 5810 26575 5813
rect 17309 5808 26575 5810
rect 17309 5752 17314 5808
rect 17370 5752 26514 5808
rect 26570 5752 26575 5808
rect 17309 5750 26575 5752
rect 17309 5747 17375 5750
rect 26509 5747 26575 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 26693 5674 26759 5677
rect 29520 5674 30000 5704
rect 26693 5672 30000 5674
rect 26693 5616 26698 5672
rect 26754 5616 30000 5672
rect 26693 5614 30000 5616
rect 26693 5611 26759 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 2037 5266 2103 5269
rect 8569 5266 8635 5269
rect 2037 5264 8635 5266
rect 2037 5208 2042 5264
rect 2098 5208 8574 5264
rect 8630 5208 8635 5264
rect 2037 5206 8635 5208
rect 2037 5203 2103 5206
rect 8569 5203 8635 5206
rect 15561 5266 15627 5269
rect 26417 5266 26483 5269
rect 15561 5264 26483 5266
rect 15561 5208 15566 5264
rect 15622 5208 26422 5264
rect 26478 5208 26483 5264
rect 15561 5206 26483 5208
rect 15561 5203 15627 5206
rect 26417 5203 26483 5206
rect 0 5130 480 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 480 5070
rect 1577 5067 1643 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 0 4450 480 4480
rect 1669 4450 1735 4453
rect 0 4448 1735 4450
rect 0 4392 1674 4448
rect 1730 4392 1735 4448
rect 0 4390 1735 4392
rect 0 4360 480 4390
rect 1669 4387 1735 4390
rect 27797 4450 27863 4453
rect 29520 4450 30000 4480
rect 27797 4448 30000 4450
rect 27797 4392 27802 4448
rect 27858 4392 30000 4448
rect 27797 4390 30000 4392
rect 27797 4387 27863 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 26785 4178 26851 4181
rect 26969 4178 27035 4181
rect 26785 4176 27035 4178
rect 26785 4120 26790 4176
rect 26846 4120 26974 4176
rect 27030 4120 27035 4176
rect 26785 4118 27035 4120
rect 26785 4115 26851 4118
rect 26969 4115 27035 4118
rect 2037 4042 2103 4045
rect 7833 4042 7899 4045
rect 2037 4040 7899 4042
rect 2037 3984 2042 4040
rect 2098 3984 7838 4040
rect 7894 3984 7899 4040
rect 2037 3982 7899 3984
rect 2037 3979 2103 3982
rect 7833 3979 7899 3982
rect 0 3906 480 3936
rect 1485 3906 1551 3909
rect 0 3904 1551 3906
rect 0 3848 1490 3904
rect 1546 3848 1551 3904
rect 0 3846 1551 3848
rect 0 3816 480 3846
rect 1485 3843 1551 3846
rect 25405 3906 25471 3909
rect 29520 3906 30000 3936
rect 25405 3904 30000 3906
rect 25405 3848 25410 3904
rect 25466 3848 30000 3904
rect 25405 3846 30000 3848
rect 25405 3843 25471 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 25773 3498 25839 3501
rect 25773 3496 26434 3498
rect 25773 3440 25778 3496
rect 25834 3440 26434 3496
rect 25773 3438 26434 3440
rect 25773 3435 25839 3438
rect 0 3362 480 3392
rect 3785 3362 3851 3365
rect 0 3360 3851 3362
rect 0 3304 3790 3360
rect 3846 3304 3851 3360
rect 0 3302 3851 3304
rect 26374 3362 26434 3438
rect 29520 3362 30000 3392
rect 26374 3302 30000 3362
rect 0 3272 480 3302
rect 3785 3299 3851 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 6913 3090 6979 3093
rect 26417 3090 26483 3093
rect 6913 3088 26483 3090
rect 6913 3032 6918 3088
rect 6974 3032 26422 3088
rect 26478 3032 26483 3088
rect 6913 3030 26483 3032
rect 6913 3027 6979 3030
rect 26417 3027 26483 3030
rect 26601 2818 26667 2821
rect 26601 2816 26802 2818
rect 26601 2760 26606 2816
rect 26662 2760 26802 2816
rect 26601 2758 26802 2760
rect 26601 2755 26667 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 26742 2682 26802 2758
rect 29520 2682 30000 2712
rect 26742 2622 30000 2682
rect 0 2592 480 2622
rect 1577 2619 1643 2622
rect 29520 2592 30000 2622
rect 7189 2410 7255 2413
rect 14917 2410 14983 2413
rect 7189 2408 14983 2410
rect 7189 2352 7194 2408
rect 7250 2352 14922 2408
rect 14978 2352 14983 2408
rect 7189 2350 14983 2352
rect 7189 2347 7255 2350
rect 14917 2347 14983 2350
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 4061 2138 4127 2141
rect 0 2136 4127 2138
rect 0 2080 4066 2136
rect 4122 2080 4127 2136
rect 0 2078 4127 2080
rect 0 2048 480 2078
rect 4061 2075 4127 2078
rect 26969 2138 27035 2141
rect 29520 2138 30000 2168
rect 26969 2136 30000 2138
rect 26969 2080 26974 2136
rect 27030 2080 30000 2136
rect 26969 2078 30000 2080
rect 26969 2075 27035 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 2681 1458 2747 1461
rect 0 1456 2747 1458
rect 0 1400 2686 1456
rect 2742 1400 2747 1456
rect 0 1398 2747 1400
rect 0 1368 480 1398
rect 2681 1395 2747 1398
rect 25865 1458 25931 1461
rect 29520 1458 30000 1488
rect 25865 1456 30000 1458
rect 25865 1400 25870 1456
rect 25926 1400 30000 1456
rect 25865 1398 30000 1400
rect 25865 1395 25931 1398
rect 29520 1368 30000 1398
rect 10409 1322 10475 1325
rect 614 1320 10475 1322
rect 614 1264 10414 1320
rect 10470 1264 10475 1320
rect 614 1262 10475 1264
rect 0 914 480 944
rect 614 914 674 1262
rect 10409 1259 10475 1262
rect 0 854 674 914
rect 27061 914 27127 917
rect 29520 914 30000 944
rect 27061 912 30000 914
rect 27061 856 27066 912
rect 27122 856 30000 912
rect 27061 854 30000 856
rect 0 824 480 854
rect 27061 851 27127 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 2221 370 2287 373
rect 0 368 2287 370
rect 0 312 2226 368
rect 2282 312 2287 368
rect 0 310 2287 312
rect 0 280 480 310
rect 2221 307 2287 310
rect 26877 370 26943 373
rect 29520 370 30000 400
rect 26877 368 30000 370
rect 26877 312 26882 368
rect 26938 312 30000 368
rect 26877 310 30000 312
rect 26877 307 26943 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 9628 19620 9692 19684
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 9628 19348 9692 19412
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 8340 16688 8404 16692
rect 8340 16632 8354 16688
rect 8354 16632 8404 16688
rect 8340 16628 8404 16632
rect 26556 16628 26620 16692
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 13308 11188 13372 11252
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 3004 10780 3068 10844
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 9627 19684 9693 19685
rect 9627 19620 9628 19684
rect 9692 19620 9693 19684
rect 9627 19619 9693 19620
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 9630 19413 9690 19619
rect 9627 19412 9693 19413
rect 9627 19348 9628 19412
rect 9692 19348 9693 19412
rect 9627 19347 9693 19348
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 3006 10845 3066 11102
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 3003 10844 3069 10845
rect 3003 10780 3004 10844
rect 3068 10780 3069 10844
rect 3003 10779 3069 10780
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
<< via4 >>
rect 8254 16692 8490 16778
rect 8254 16628 8340 16692
rect 8340 16628 8404 16692
rect 8404 16628 8490 16692
rect 8254 16542 8490 16628
rect 2918 11102 3154 11338
rect 13222 11252 13458 11338
rect 13222 11188 13308 11252
rect 13308 11188 13372 11252
rect 13372 11188 13458 11252
rect 13222 11102 13458 11188
rect 26470 16692 26706 16778
rect 26470 16628 26556 16692
rect 26556 16628 26620 16692
rect 26620 16628 26706 16692
rect 26470 16542 26706 16628
<< metal5 >>
rect 8212 16778 26748 16820
rect 8212 16542 8254 16778
rect 8490 16542 26470 16778
rect 26706 16542 26748 16778
rect 8212 16500 26748 16542
rect 2876 11338 13500 11380
rect 2876 11102 2918 11338
rect 3154 11102 13222 11338
rect 13458 11102 13500 11338
rect 2876 11060 13500 11102
use scs8hd_buf_2  _47_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__47__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_11
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_82 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_279
timestamp 1586364061
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_283
timestamp 1586364061
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_295
timestamp 1586364061
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_298 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 28520 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_296
timestamp 1586364061
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_296
timestamp 1586364061
transform 1 0 28336 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_29
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_41
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_279
timestamp 1586364061
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_283
timestamp 1586364061
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_287
timestamp 1586364061
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_280
timestamp 1586364061
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_6_292
timestamp 1586364061
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_279
timestamp 1586364061
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_283
timestamp 1586364061
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_295
timestamp 1586364061
transform 1 0 28244 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_298
timestamp 1586364061
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_280
timestamp 1586364061
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_292
timestamp 1586364061
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_298
timestamp 1586364061
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_54
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 590 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 27508 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_279
timestamp 1586364061
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_283
timestamp 1586364061
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_291
timestamp 1586364061
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_295
timestamp 1586364061
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2668 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_256
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 590 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_262
timestamp 1586364061
transform 1 0 25208 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_280
timestamp 1586364061
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_292
timestamp 1586364061
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_298
timestamp 1586364061
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1472 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_211
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_223
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 774 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_255
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_259
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_271
timestamp 1586364061
transform 1 0 26036 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 27508 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_279
timestamp 1586364061
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_283
timestamp 1586364061
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_291
timestamp 1586364061
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_295
timestamp 1586364061
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _19_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_183
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_225
timestamp 1586364061
transform 1 0 21804 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_229
timestamp 1586364061
transform 1 0 22172 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_241
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_245
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_249
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_280
timestamp 1586364061
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_292
timestamp 1586364061
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_298
timestamp 1586364061
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_1.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_37
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_41
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_109
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18124 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_194
timestamp 1586364061
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_215
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_211
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_221
timestamp 1586364061
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_219
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_3_
timestamp 1586364061
transform 1 0 21620 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_2_
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l4_in_0_
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_256
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_240
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_262
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_270
timestamp 1586364061
transform 1 0 25944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_272
timestamp 1586364061
transform 1 0 26128 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_268
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 26128 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 406 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_280
timestamp 1586364061
transform 1 0 26864 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_283
timestamp 1586364061
transform 1 0 27140 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_279
timestamp 1586364061
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 27048 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 27508 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_296
timestamp 1586364061
transform 1 0 28336 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_295
timestamp 1586364061
transform 1 0 28244 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_291
timestamp 1586364061
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_284
timestamp 1586364061
transform 1 0 27232 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_43
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_48
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_78
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_177
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_181
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_192
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_209
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_228
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_264
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 27508 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_285
timestamp 1586364061
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_289
timestamp 1586364061
transform 1 0 27692 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 590 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_8
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_100
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_140
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_2_
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_175
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l4_in_0_
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_196
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l3_in_1_
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_222
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_226
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_3_
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_243
timestamp 1586364061
transform 1 0 23460 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_256
timestamp 1586364061
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_260
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_285
timestamp 1586364061
transform 1 0 27324 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_297
timestamp 1586364061
transform 1 0 28428 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_9
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_10.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_230
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 26128 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_261
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_265
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_268
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_291
timestamp 1586364061
transform 1 0 27876 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_295
timestamp 1586364061
transform 1 0 28244 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_57
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_78
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9752 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_103
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_146
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_162
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_201
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_209
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_212
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_234
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_238
timestamp 1586364061
transform 1 0 23000 0 -1 12512
box -38 -48 590 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_248
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_252
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_265
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_269
timestamp 1586364061
transform 1 0 25852 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_285
timestamp 1586364061
transform 1 0 27324 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_297
timestamp 1586364061
transform 1 0 28428 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1786 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_22
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_26
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_76
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_76
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 314 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_85
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_91
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_101
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_164
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_171
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_196
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 130 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_11.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_219
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_238
timestamp 1586364061
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23184 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23736 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l3_in_1_
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_267
timestamp 1586364061
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_285
timestamp 1586364061
transform 1 0 27324 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_284
timestamp 1586364061
transform 1 0 27232 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_280
timestamp 1586364061
transform 1 0 26864 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 27416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 27048 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_289
timestamp 1586364061
transform 1 0 27692 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_295
timestamp 1586364061
transform 1 0 28244 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_291
timestamp 1586364061
transform 1 0 27876 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 27508 0 -1 13600
box -38 -48 222 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 27600 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_297
timestamp 1586364061
transform 1 0 28428 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_140
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_148
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 130 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_199
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_203
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_216
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_233
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_237
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_241
timestamp 1586364061
transform 1 0 23276 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_251
timestamp 1586364061
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_272
timestamp 1586364061
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_3_
timestamp 1586364061
transform 1 0 26864 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 26680 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 27876 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 28244 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_289
timestamp 1586364061
transform 1 0 27692 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_293
timestamp 1586364061
transform 1 0 28060 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_297
timestamp 1586364061
transform 1 0 28428 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 14688
box -38 -48 1786 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_42
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_135
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_139
timestamp 1586364061
transform 1 0 13892 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_182
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_188
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_192
timestamp 1586364061
transform 1 0 18768 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21528 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21344 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_219
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_22_266
timestamp 1586364061
transform 1 0 25576 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_262
timestamp 1586364061
transform 1 0 25208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_258
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25392 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 25024 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25760 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l4_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_285
timestamp 1586364061
transform 1 0 27324 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_297
timestamp 1586364061
transform 1 0 28428 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 1786 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_26
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_84
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_88
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_115
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_119
timestamp 1586364061
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_129
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_142
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_23_190
timestamp 1586364061
transform 1 0 18584 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_233
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 26128 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_260
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_264
timestamp 1586364061
transform 1 0 25392 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_268
timestamp 1586364061
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 28060 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_291
timestamp 1586364061
transform 1 0 27876 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_295
timestamp 1586364061
transform 1 0 28244 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_16
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_20
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_24
timestamp 1586364061
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_139
timestamp 1586364061
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_173
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_177
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_185
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_209
timestamp 1586364061
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 21344 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_222
timestamp 1586364061
transform 1 0 21528 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_245
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_249
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_253
timestamp 1586364061
transform 1 0 24380 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 15776
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_2_
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 26128 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_267
timestamp 1586364061
transform 1 0 25668 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 27508 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_285
timestamp 1586364061
transform 1 0 27324 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_289
timestamp 1586364061
transform 1 0 27692 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_297
timestamp 1586364061
transform 1 0 28428 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_170
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_238
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 26128 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_264
timestamp 1586364061
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_268
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 28060 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_291
timestamp 1586364061
transform 1 0 27876 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_295
timestamp 1586364061
transform 1 0 28244 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_54
timestamp 1586364061
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_50
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_67
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_122
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_144
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_139
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_168
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_172
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_176
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_185
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_212
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_221
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l4_in_0_
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_238
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21620 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_242
timestamp 1586364061
transform 1 0 23368 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_255
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 -1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24012 0 1 16864
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_26_267
timestamp 1586364061
transform 1 0 25668 0 -1 16864
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25944 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_271
timestamp 1586364061
transform 1 0 26036 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_268
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_272
timestamp 1586364061
transform 1 0 26128 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 26312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l1_in_2_
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_285
timestamp 1586364061
transform 1 0 27324 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_285
timestamp 1586364061
transform 1 0 27324 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_293
timestamp 1586364061
transform 1 0 28060 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_289
timestamp 1586364061
transform 1 0 27692 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_289
timestamp 1586364061
transform 1 0 27692 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 27508 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 28244 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 27876 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 27508 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_297
timestamp 1586364061
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_297
timestamp 1586364061
transform 1 0 28428 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1472 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_2_
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_185
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 21528 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_220
timestamp 1586364061
transform 1 0 21344 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_247
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_255
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24840 0 -1 17952
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_285
timestamp 1586364061
transform 1 0 27324 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_297
timestamp 1586364061
transform 1 0 28428 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1472 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_13
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_30
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 1786 592
use scs8hd_conb_1  _16_
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_100
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_104
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_188
timestamp 1586364061
transform 1 0 18400 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_200
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_3_
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_223
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23920 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 25484 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_261
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 27416 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 27784 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 28152 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_284
timestamp 1586364061
transform 1 0 27232 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_288
timestamp 1586364061
transform 1 0 27600 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_292
timestamp 1586364061
transform 1 0 27968 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_296
timestamp 1586364061
transform 1 0 28336 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_14
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_22
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_26
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_50
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_74
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 590 592
use scs8hd_buf_1  mux_bottom_ipin_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_4  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_109
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_136
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_148
timestamp 1586364061
transform 1 0 14720 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_164
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_174
timestamp 1586364061
transform 1 0 17112 0 -1 19040
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 17848 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_201
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_6  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_12.mux_l2_in_2_
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 21804 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_236
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23920 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23736 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23368 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_244
timestamp 1586364061
transform 1 0 23552 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_2_
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_285
timestamp 1586364061
transform 1 0 27324 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_297
timestamp 1586364061
transform 1 0 28428 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_14
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_25
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_41
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_6.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_120
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_146
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_191
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_ipin_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_222
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_228
timestamp 1586364061
transform 1 0 22080 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l4_in_0_
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 24012 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_251
timestamp 1586364061
transform 1 0 24196 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l2_in_3_
timestamp 1586364061
transform 1 0 26312 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_264
timestamp 1586364061
transform 1 0 25392 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_270
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 27324 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_283
timestamp 1586364061
transform 1 0 27140 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_287
timestamp 1586364061
transform 1 0 27508 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 11960 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_107
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_175
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_198
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 23920 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_247
timestamp 1586364061
transform 1 0 23828 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_250
timestamp 1586364061
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_254
timestamp 1586364061
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 25852 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_271
timestamp 1586364061
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_279
timestamp 1586364061
transform 1 0 26772 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_291
timestamp 1586364061
transform 1 0 27876 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 590 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_43
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6900 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_66
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_70
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_82
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_88
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_92
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_126
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_130
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_148
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_ipin_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_34_158
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_161
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_169
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_170
timestamp 1586364061
transform 1 0 16744 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_ipin_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_194
timestamp 1586364061
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_191
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 19136 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_ipin_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_34_198
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_182
timestamp 1586364061
transform 1 0 17848 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_205
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_216
timestamp 1586364061
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_210
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_253
timestamp 1586364061
transform 1 0 24380 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_247
timestamp 1586364061
transform 1 0 23828 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24012 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_ipin_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24104 0 -1 21216
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_ipin_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24196 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_264
timestamp 1586364061
transform 1 0 25392 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_260
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 25576 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_ipin_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25116 0 -1 21216
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_13.mux_l3_in_1_
timestamp 1586364061
transform 1 0 25484 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_272
timestamp 1586364061
transform 1 0 26128 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_268
timestamp 1586364061
transform 1 0 25760 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_274
timestamp 1586364061
transform 1 0 26312 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_286
timestamp 1586364061
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_288
timestamp 1586364061
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_296
timestamp 1586364061
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_298
timestamp 1586364061
transform 1 0 28520 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_242
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_249
timestamp 1586364061
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_261
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_273
timestamp 1586364061
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_280
timestamp 1586364061
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_292
timestamp 1586364061
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_298
timestamp 1586364061
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 14922 0 14978 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 24950 0 25006 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 prog_clk
port 82 nsew default input
rlabel metal2 s 938 23520 994 24000 6 top_grid_pin_16_
port 83 nsew default tristate
rlabel metal2 s 2778 23520 2834 24000 6 top_grid_pin_17_
port 84 nsew default tristate
rlabel metal2 s 4618 23520 4674 24000 6 top_grid_pin_18_
port 85 nsew default tristate
rlabel metal2 s 6550 23520 6606 24000 6 top_grid_pin_19_
port 86 nsew default tristate
rlabel metal2 s 8390 23520 8446 24000 6 top_grid_pin_20_
port 87 nsew default tristate
rlabel metal2 s 10230 23520 10286 24000 6 top_grid_pin_21_
port 88 nsew default tristate
rlabel metal2 s 12162 23520 12218 24000 6 top_grid_pin_22_
port 89 nsew default tristate
rlabel metal2 s 14002 23520 14058 24000 6 top_grid_pin_23_
port 90 nsew default tristate
rlabel metal2 s 15934 23520 15990 24000 6 top_grid_pin_24_
port 91 nsew default tristate
rlabel metal2 s 17774 23520 17830 24000 6 top_grid_pin_25_
port 92 nsew default tristate
rlabel metal2 s 19614 23520 19670 24000 6 top_grid_pin_26_
port 93 nsew default tristate
rlabel metal2 s 21546 23520 21602 24000 6 top_grid_pin_27_
port 94 nsew default tristate
rlabel metal2 s 23386 23520 23442 24000 6 top_grid_pin_28_
port 95 nsew default tristate
rlabel metal2 s 25226 23520 25282 24000 6 top_grid_pin_29_
port 96 nsew default tristate
rlabel metal2 s 27158 23520 27214 24000 6 top_grid_pin_30_
port 97 nsew default tristate
rlabel metal2 s 28998 23520 29054 24000 6 top_grid_pin_31_
port 98 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 vpwr
port 99 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 vgnd
port 100 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
