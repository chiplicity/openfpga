magic
tech sky130A
magscale 1 2
timestamp 1605129599
<< locali >>
rect 14933 33303 14967 33405
rect 12909 30651 12943 30821
rect 17509 30583 17543 30753
rect 3341 28407 3375 28713
rect 16313 27931 16347 28033
rect 31953 27931 31987 28033
rect 34529 22015 34563 22185
rect 31585 20247 31619 20553
rect 24225 15963 24259 16201
rect 34529 14943 34563 15113
<< viali >>
rect 7021 36873 7055 36907
rect 6837 36669 6871 36703
rect 7481 36533 7515 36567
rect 22661 36261 22695 36295
rect 6837 36193 6871 36227
rect 15669 36193 15703 36227
rect 23857 36193 23891 36227
rect 15761 36125 15795 36159
rect 15945 36125 15979 36159
rect 22753 36125 22787 36159
rect 22937 36125 22971 36159
rect 7021 35989 7055 36023
rect 14013 35989 14047 36023
rect 15301 35989 15335 36023
rect 21465 35989 21499 36023
rect 22293 35989 22327 36023
rect 24041 35989 24075 36023
rect 24961 35989 24995 36023
rect 26709 35989 26743 36023
rect 5641 35785 5675 35819
rect 7757 35785 7791 35819
rect 8401 35785 8435 35819
rect 15945 35785 15979 35819
rect 22477 35785 22511 35819
rect 22845 35785 22879 35819
rect 24685 35785 24719 35819
rect 35633 35785 35667 35819
rect 15669 35717 15703 35751
rect 21373 35717 21407 35751
rect 23121 35717 23155 35751
rect 22017 35649 22051 35683
rect 26893 35649 26927 35683
rect 5457 35581 5491 35615
rect 7113 35581 7147 35615
rect 8217 35581 8251 35615
rect 13921 35581 13955 35615
rect 16313 35581 16347 35615
rect 21741 35581 21775 35615
rect 23673 35581 23707 35615
rect 24225 35581 24259 35615
rect 24961 35581 24995 35615
rect 25881 35581 25915 35615
rect 26709 35581 26743 35615
rect 35449 35581 35483 35615
rect 36001 35581 36035 35615
rect 8861 35513 8895 35547
rect 13829 35513 13863 35547
rect 14166 35513 14200 35547
rect 21833 35513 21867 35547
rect 26249 35513 26283 35547
rect 26801 35513 26835 35547
rect 6101 35445 6135 35479
rect 7297 35445 7331 35479
rect 12449 35445 12483 35479
rect 15301 35445 15335 35479
rect 20913 35445 20947 35479
rect 21189 35445 21223 35479
rect 23857 35445 23891 35479
rect 25145 35445 25179 35479
rect 26341 35445 26375 35479
rect 1593 35241 1627 35275
rect 4353 35241 4387 35275
rect 7113 35241 7147 35275
rect 13277 35241 13311 35275
rect 14749 35241 14783 35275
rect 15301 35241 15335 35275
rect 19717 35241 19751 35275
rect 21189 35241 21223 35275
rect 23489 35241 23523 35275
rect 24869 35241 24903 35275
rect 25237 35241 25271 35275
rect 35541 35241 35575 35275
rect 9689 35173 9723 35207
rect 22376 35173 22410 35207
rect 1409 35105 1443 35139
rect 4169 35105 4203 35139
rect 5529 35105 5563 35139
rect 8309 35105 8343 35139
rect 9873 35105 9907 35139
rect 11796 35105 11830 35139
rect 13737 35105 13771 35139
rect 15669 35105 15703 35139
rect 17233 35105 17267 35139
rect 18429 35105 18463 35139
rect 21005 35105 21039 35139
rect 26781 35105 26815 35139
rect 35357 35105 35391 35139
rect 5273 35037 5307 35071
rect 11529 35037 11563 35071
rect 15761 35037 15795 35071
rect 15853 35037 15887 35071
rect 17325 35037 17359 35071
rect 17417 35037 17451 35071
rect 22109 35037 22143 35071
rect 24777 35037 24811 35071
rect 25329 35037 25363 35071
rect 25421 35037 25455 35071
rect 26525 35037 26559 35071
rect 16865 34969 16899 35003
rect 18153 34969 18187 35003
rect 24317 34969 24351 35003
rect 6653 34901 6687 34935
rect 7481 34901 7515 34935
rect 8493 34901 8527 34935
rect 10057 34901 10091 34935
rect 10333 34901 10367 34935
rect 12909 34901 12943 34935
rect 13921 34901 13955 34935
rect 18613 34901 18647 34935
rect 21557 34901 21591 34935
rect 24041 34901 24075 34935
rect 27905 34901 27939 34935
rect 1593 34697 1627 34731
rect 2053 34697 2087 34731
rect 3801 34697 3835 34731
rect 4261 34697 4295 34731
rect 9137 34697 9171 34731
rect 9505 34697 9539 34731
rect 10609 34697 10643 34731
rect 11713 34697 11747 34731
rect 14197 34697 14231 34731
rect 14657 34697 14691 34731
rect 16129 34697 16163 34731
rect 16405 34697 16439 34731
rect 17417 34697 17451 34731
rect 19165 34697 19199 34731
rect 21005 34697 21039 34731
rect 22569 34697 22603 34731
rect 22845 34697 22879 34731
rect 23949 34697 23983 34731
rect 25789 34697 25823 34731
rect 26157 34697 26191 34731
rect 26525 34697 26559 34731
rect 27997 34697 28031 34731
rect 35633 34697 35667 34731
rect 36737 34697 36771 34731
rect 2697 34629 2731 34663
rect 5181 34629 5215 34663
rect 8769 34629 8803 34663
rect 13921 34629 13955 34663
rect 16773 34629 16807 34663
rect 18061 34629 18095 34663
rect 19625 34629 19659 34663
rect 3157 34561 3191 34595
rect 4629 34561 4663 34595
rect 5825 34561 5859 34595
rect 10149 34561 10183 34595
rect 12265 34561 12299 34595
rect 14749 34561 14783 34595
rect 16957 34561 16991 34595
rect 18521 34561 18555 34595
rect 18705 34561 18739 34595
rect 20177 34561 20211 34595
rect 20729 34561 20763 34595
rect 24317 34561 24351 34595
rect 1409 34493 1443 34527
rect 2513 34493 2547 34527
rect 3617 34493 3651 34527
rect 6561 34493 6595 34527
rect 7389 34493 7423 34527
rect 10057 34493 10091 34527
rect 10977 34493 11011 34527
rect 12541 34493 12575 34527
rect 12808 34493 12842 34527
rect 17785 34493 17819 34527
rect 19441 34493 19475 34527
rect 19993 34493 20027 34527
rect 21189 34493 21223 34527
rect 21456 34493 21490 34527
rect 24409 34493 24443 34527
rect 24665 34493 24699 34527
rect 26617 34493 26651 34527
rect 26873 34493 26907 34527
rect 35357 34493 35391 34527
rect 35449 34493 35483 34527
rect 36001 34493 36035 34527
rect 36553 34493 36587 34527
rect 37105 34493 37139 34527
rect 5549 34425 5583 34459
rect 7634 34425 7668 34459
rect 9965 34425 9999 34459
rect 14994 34425 15028 34459
rect 18429 34425 18463 34459
rect 20085 34425 20119 34459
rect 5089 34357 5123 34391
rect 5641 34357 5675 34391
rect 6285 34357 6319 34391
rect 7205 34357 7239 34391
rect 9597 34357 9631 34391
rect 11161 34357 11195 34391
rect 28365 34357 28399 34391
rect 4537 34153 4571 34187
rect 5641 34153 5675 34187
rect 6009 34153 6043 34187
rect 9137 34153 9171 34187
rect 13277 34153 13311 34187
rect 14013 34153 14047 34187
rect 14105 34153 14139 34187
rect 20085 34153 20119 34187
rect 22293 34153 22327 34187
rect 23581 34153 23615 34187
rect 25053 34153 25087 34187
rect 25513 34153 25547 34187
rect 35633 34153 35667 34187
rect 1685 34085 1719 34119
rect 6368 34085 6402 34119
rect 9505 34085 9539 34119
rect 9956 34085 9990 34119
rect 18052 34085 18086 34119
rect 19717 34085 19751 34119
rect 23918 34085 23952 34119
rect 27138 34085 27172 34119
rect 4905 34017 4939 34051
rect 8493 34017 8527 34051
rect 11529 34017 11563 34051
rect 12153 34017 12187 34051
rect 15557 34017 15591 34051
rect 21169 34017 21203 34051
rect 22661 34017 22695 34051
rect 23673 34017 23707 34051
rect 35449 34017 35483 34051
rect 4997 33949 5031 33983
rect 5089 33949 5123 33983
rect 6101 33949 6135 33983
rect 9689 33949 9723 33983
rect 11897 33949 11931 33983
rect 15301 33949 15335 33983
rect 17785 33949 17819 33983
rect 20913 33949 20947 33983
rect 26893 33949 26927 33983
rect 4445 33881 4479 33915
rect 2973 33813 3007 33847
rect 3893 33813 3927 33847
rect 7481 33813 7515 33847
rect 8677 33813 8711 33847
rect 11069 33813 11103 33847
rect 14749 33813 14783 33847
rect 16681 33813 16715 33847
rect 17049 33813 17083 33847
rect 17417 33813 17451 33847
rect 19165 33813 19199 33847
rect 25881 33813 25915 33847
rect 26801 33813 26835 33847
rect 28273 33813 28307 33847
rect 5825 33609 5859 33643
rect 6101 33609 6135 33643
rect 6837 33609 6871 33643
rect 9965 33609 9999 33643
rect 10241 33609 10275 33643
rect 15117 33609 15151 33643
rect 17877 33609 17911 33643
rect 20177 33609 20211 33643
rect 22017 33609 22051 33643
rect 22385 33609 22419 33643
rect 22753 33609 22787 33643
rect 23489 33609 23523 33643
rect 25237 33609 25271 33643
rect 25421 33609 25455 33643
rect 26801 33609 26835 33643
rect 35633 33609 35667 33643
rect 6561 33541 6595 33575
rect 10793 33541 10827 33575
rect 23121 33541 23155 33575
rect 2421 33473 2455 33507
rect 3525 33473 3559 33507
rect 7389 33473 7423 33507
rect 8493 33473 8527 33507
rect 11345 33473 11379 33507
rect 11805 33473 11839 33507
rect 13001 33473 13035 33507
rect 13461 33473 13495 33507
rect 15672 33473 15706 33507
rect 15945 33473 15979 33507
rect 24225 33473 24259 33507
rect 25973 33473 26007 33507
rect 36001 33473 36035 33507
rect 3249 33405 3283 33439
rect 4445 33405 4479 33439
rect 8585 33405 8619 33439
rect 8852 33405 8886 33439
rect 10701 33405 10735 33439
rect 11161 33405 11195 33439
rect 11253 33405 11287 33439
rect 12817 33405 12851 33439
rect 14105 33405 14139 33439
rect 14933 33405 14967 33439
rect 15209 33405 15243 33439
rect 15532 33405 15566 33439
rect 18061 33405 18095 33439
rect 20637 33405 20671 33439
rect 25789 33405 25823 33439
rect 26525 33405 26559 33439
rect 26985 33405 27019 33439
rect 27252 33405 27286 33439
rect 35449 33405 35483 33439
rect 2789 33337 2823 33371
rect 3985 33337 4019 33371
rect 4353 33337 4387 33371
rect 4712 33337 4746 33371
rect 7297 33337 7331 33371
rect 7849 33337 7883 33371
rect 12265 33337 12299 33371
rect 12909 33337 12943 33371
rect 14749 33337 14783 33371
rect 18328 33337 18362 33371
rect 20545 33337 20579 33371
rect 20904 33337 20938 33371
rect 24133 33337 24167 33371
rect 25881 33337 25915 33371
rect 1777 33269 1811 33303
rect 2881 33269 2915 33303
rect 3341 33269 3375 33303
rect 7205 33269 7239 33303
rect 12449 33269 12483 33303
rect 14197 33269 14231 33303
rect 14933 33269 14967 33303
rect 17049 33269 17083 33303
rect 17509 33269 17543 33303
rect 19441 33269 19475 33303
rect 19809 33269 19843 33303
rect 23673 33269 23707 33303
rect 24041 33269 24075 33303
rect 24685 33269 24719 33303
rect 28365 33269 28399 33303
rect 28641 33269 28675 33303
rect 35357 33269 35391 33303
rect 3801 33065 3835 33099
rect 5457 33065 5491 33099
rect 6469 33065 6503 33099
rect 7573 33065 7607 33099
rect 9045 33065 9079 33099
rect 10885 33065 10919 33099
rect 11253 33065 11287 33099
rect 12357 33065 12391 33099
rect 12909 33065 12943 33099
rect 13645 33065 13679 33099
rect 14749 33065 14783 33099
rect 15117 33065 15151 33099
rect 19349 33065 19383 33099
rect 22293 33065 22327 33099
rect 23489 33065 23523 33099
rect 24685 33065 24719 33099
rect 24869 33065 24903 33099
rect 27077 33065 27111 33099
rect 6009 32997 6043 33031
rect 9413 32997 9447 33031
rect 10241 32997 10275 33031
rect 12265 32997 12299 33031
rect 27436 32997 27470 33031
rect 2033 32929 2067 32963
rect 4333 32929 4367 32963
rect 6929 32929 6963 32963
rect 8493 32929 8527 32963
rect 9689 32929 9723 32963
rect 14013 32929 14047 32963
rect 15301 32929 15335 32963
rect 15624 32929 15658 32963
rect 16037 32929 16071 32963
rect 18236 32929 18270 32963
rect 21169 32929 21203 32963
rect 25237 32929 25271 32963
rect 27169 32929 27203 32963
rect 29377 32929 29411 32963
rect 1777 32861 1811 32895
rect 4077 32861 4111 32895
rect 7021 32861 7055 32895
rect 7205 32861 7239 32895
rect 12541 32861 12575 32895
rect 14105 32861 14139 32895
rect 14289 32861 14323 32895
rect 15764 32861 15798 32895
rect 17785 32861 17819 32895
rect 17969 32861 18003 32895
rect 20913 32861 20947 32895
rect 23581 32861 23615 32895
rect 23673 32861 23707 32895
rect 25329 32861 25363 32895
rect 25421 32861 25455 32895
rect 3157 32793 3191 32827
rect 8677 32793 8711 32827
rect 11897 32793 11931 32827
rect 23121 32793 23155 32827
rect 1593 32725 1627 32759
rect 3525 32725 3559 32759
rect 6561 32725 6595 32759
rect 9873 32725 9907 32759
rect 11713 32725 11747 32759
rect 17141 32725 17175 32759
rect 20637 32725 20671 32759
rect 24133 32725 24167 32759
rect 28549 32725 28583 32759
rect 29561 32725 29595 32759
rect 1777 32521 1811 32555
rect 3249 32521 3283 32555
rect 5549 32521 5583 32555
rect 6285 32521 6319 32555
rect 7849 32521 7883 32555
rect 11621 32521 11655 32555
rect 12633 32521 12667 32555
rect 13277 32521 13311 32555
rect 14197 32521 14231 32555
rect 14381 32521 14415 32555
rect 15485 32521 15519 32555
rect 16221 32521 16255 32555
rect 20177 32521 20211 32555
rect 20637 32521 20671 32555
rect 22477 32521 22511 32555
rect 23213 32521 23247 32555
rect 25237 32521 25271 32555
rect 26249 32521 26283 32555
rect 26801 32521 26835 32555
rect 27813 32521 27847 32555
rect 28641 32521 28675 32555
rect 29469 32521 29503 32555
rect 3893 32453 3927 32487
rect 5825 32453 5859 32487
rect 6837 32453 6871 32487
rect 8309 32453 8343 32487
rect 11989 32453 12023 32487
rect 15761 32453 15795 32487
rect 22753 32453 22787 32487
rect 28181 32453 28215 32487
rect 4629 32385 4663 32419
rect 7389 32385 7423 32419
rect 8953 32385 8987 32419
rect 13737 32385 13771 32419
rect 14933 32385 14967 32419
rect 16957 32385 16991 32419
rect 21097 32385 21131 32419
rect 24225 32385 24259 32419
rect 25789 32385 25823 32419
rect 26709 32385 26743 32419
rect 27261 32385 27295 32419
rect 27353 32385 27387 32419
rect 1869 32317 1903 32351
rect 4445 32317 4479 32351
rect 5641 32317 5675 32351
rect 8769 32317 8803 32351
rect 9689 32317 9723 32351
rect 14749 32317 14783 32351
rect 14841 32317 14875 32351
rect 16405 32317 16439 32351
rect 16681 32317 16715 32351
rect 18061 32317 18095 32351
rect 19809 32317 19843 32351
rect 24041 32317 24075 32351
rect 27169 32317 27203 32351
rect 2136 32249 2170 32283
rect 7297 32249 7331 32283
rect 8861 32249 8895 32283
rect 17509 32249 17543 32283
rect 18306 32249 18340 32283
rect 21342 32249 21376 32283
rect 24777 32249 24811 32283
rect 25605 32249 25639 32283
rect 3617 32181 3651 32215
rect 4077 32181 4111 32215
rect 4537 32181 4571 32215
rect 5089 32181 5123 32215
rect 6561 32181 6595 32215
rect 7205 32181 7239 32215
rect 8401 32181 8435 32215
rect 17877 32181 17911 32215
rect 19441 32181 19475 32215
rect 20913 32181 20947 32215
rect 23673 32181 23707 32215
rect 24133 32181 24167 32215
rect 25145 32181 25179 32215
rect 25697 32181 25731 32215
rect 2789 31977 2823 32011
rect 3249 31977 3283 32011
rect 4077 31977 4111 32011
rect 5181 31977 5215 32011
rect 5825 31977 5859 32011
rect 6929 31977 6963 32011
rect 7297 31977 7331 32011
rect 9045 31977 9079 32011
rect 13737 31977 13771 32011
rect 14841 31977 14875 32011
rect 16129 31977 16163 32011
rect 17785 31977 17819 32011
rect 18889 31977 18923 32011
rect 22477 31977 22511 32011
rect 23121 31977 23155 32011
rect 23489 31977 23523 32011
rect 23949 31977 23983 32011
rect 24225 31977 24259 32011
rect 24777 31977 24811 32011
rect 25881 31977 25915 32011
rect 26893 31977 26927 32011
rect 35633 31977 35667 32011
rect 4445 31909 4479 31943
rect 6561 31909 6595 31943
rect 7573 31909 7607 31943
rect 11244 31909 11278 31943
rect 14473 31909 14507 31943
rect 15853 31909 15887 31943
rect 20729 31909 20763 31943
rect 25329 31909 25363 31943
rect 27344 31909 27378 31943
rect 1676 31841 1710 31875
rect 4537 31841 4571 31875
rect 5641 31841 5675 31875
rect 8493 31841 8527 31875
rect 10977 31841 11011 31875
rect 18153 31841 18187 31875
rect 21364 31841 21398 31875
rect 23305 31841 23339 31875
rect 25237 31841 25271 31875
rect 27077 31841 27111 31875
rect 35449 31841 35483 31875
rect 1409 31773 1443 31807
rect 4629 31773 4663 31807
rect 9505 31773 9539 31807
rect 15301 31773 15335 31807
rect 18245 31773 18279 31807
rect 18337 31773 18371 31807
rect 21097 31773 21131 31807
rect 25513 31773 25547 31807
rect 8677 31705 8711 31739
rect 3709 31637 3743 31671
rect 12357 31637 12391 31671
rect 24869 31637 24903 31671
rect 28457 31637 28491 31671
rect 3433 31433 3467 31467
rect 4721 31433 4755 31467
rect 6193 31433 6227 31467
rect 7021 31433 7055 31467
rect 8493 31433 8527 31467
rect 8769 31433 8803 31467
rect 10885 31433 10919 31467
rect 11897 31433 11931 31467
rect 12633 31433 12667 31467
rect 13093 31433 13127 31467
rect 16497 31433 16531 31467
rect 17049 31433 17083 31467
rect 17877 31433 17911 31467
rect 18613 31433 18647 31467
rect 20821 31433 20855 31467
rect 21465 31433 21499 31467
rect 23397 31433 23431 31467
rect 24133 31433 24167 31467
rect 25605 31433 25639 31467
rect 26249 31433 26283 31467
rect 26709 31433 26743 31467
rect 2789 31365 2823 31399
rect 12173 31365 12207 31399
rect 14749 31365 14783 31399
rect 16865 31365 16899 31399
rect 25329 31365 25363 31399
rect 1409 31297 1443 31331
rect 3157 31297 3191 31331
rect 4169 31297 4203 31331
rect 5733 31297 5767 31331
rect 9965 31297 9999 31331
rect 22017 31297 22051 31331
rect 6837 31229 6871 31263
rect 7389 31229 7423 31263
rect 8217 31229 8251 31263
rect 8953 31229 8987 31263
rect 10517 31229 10551 31263
rect 11161 31229 11195 31263
rect 11253 31229 11287 31263
rect 12449 31229 12483 31263
rect 13553 31229 13587 31263
rect 14105 31229 14139 31263
rect 14933 31229 14967 31263
rect 15209 31229 15243 31263
rect 15485 31229 15519 31263
rect 16037 31229 16071 31263
rect 17233 31229 17267 31263
rect 21833 31229 21867 31263
rect 24593 31229 24627 31263
rect 26801 31229 26835 31263
rect 27057 31229 27091 31263
rect 1676 31161 1710 31195
rect 3985 31161 4019 31195
rect 5641 31161 5675 31195
rect 9321 31161 9355 31195
rect 9873 31161 9907 31195
rect 18245 31161 18279 31195
rect 21189 31161 21223 31195
rect 21925 31161 21959 31195
rect 24501 31161 24535 31195
rect 24777 31161 24811 31195
rect 3617 31093 3651 31127
rect 4077 31093 4111 31127
rect 5089 31093 5123 31127
rect 5181 31093 5215 31127
rect 5549 31093 5583 31127
rect 9413 31093 9447 31127
rect 9781 31093 9815 31127
rect 10977 31093 11011 31127
rect 11437 31093 11471 31127
rect 13737 31093 13771 31127
rect 15669 31093 15703 31127
rect 24961 31093 24995 31127
rect 28181 31093 28215 31127
rect 35449 31093 35483 31127
rect 2053 30889 2087 30923
rect 3709 30889 3743 30923
rect 4445 30889 4479 30923
rect 10701 30889 10735 30923
rect 12725 30889 12759 30923
rect 13093 30889 13127 30923
rect 13553 30889 13587 30923
rect 14381 30889 14415 30923
rect 17785 30889 17819 30923
rect 21097 30889 21131 30923
rect 21557 30889 21591 30923
rect 21925 30889 21959 30923
rect 22753 30889 22787 30923
rect 24317 30889 24351 30923
rect 24777 30889 24811 30923
rect 25513 30889 25547 30923
rect 35633 30889 35667 30923
rect 2329 30821 2363 30855
rect 5632 30821 5666 30855
rect 12909 30821 12943 30855
rect 13369 30821 13403 30855
rect 15822 30821 15856 30855
rect 4261 30753 4295 30787
rect 4905 30753 4939 30787
rect 8677 30753 8711 30787
rect 9689 30753 9723 30787
rect 10241 30753 10275 30787
rect 10793 30753 10827 30787
rect 11049 30753 11083 30787
rect 5365 30685 5399 30719
rect 9505 30685 9539 30719
rect 13185 30753 13219 30787
rect 14565 30753 14599 30787
rect 15117 30753 15151 30787
rect 17509 30753 17543 30787
rect 18153 30753 18187 30787
rect 18245 30753 18279 30787
rect 22569 30753 22603 30787
rect 26525 30753 26559 30787
rect 35449 30753 35483 30787
rect 15577 30685 15611 30719
rect 1685 30617 1719 30651
rect 7021 30617 7055 30651
rect 9873 30617 9907 30651
rect 12173 30617 12207 30651
rect 12909 30617 12943 30651
rect 16957 30617 16991 30651
rect 18337 30685 18371 30719
rect 24869 30685 24903 30719
rect 25053 30685 25087 30719
rect 26709 30617 26743 30651
rect 3065 30549 3099 30583
rect 5273 30549 5307 30583
rect 6745 30549 6779 30583
rect 8493 30549 8527 30583
rect 14289 30549 14323 30583
rect 17233 30549 17267 30583
rect 17509 30549 17543 30583
rect 17601 30549 17635 30583
rect 18889 30549 18923 30583
rect 24409 30549 24443 30583
rect 27077 30549 27111 30583
rect 27445 30549 27479 30583
rect 32505 30549 32539 30583
rect 1593 30345 1627 30379
rect 2973 30345 3007 30379
rect 3985 30345 4019 30379
rect 6837 30345 6871 30379
rect 9873 30345 9907 30379
rect 13737 30345 13771 30379
rect 22569 30345 22603 30379
rect 24685 30345 24719 30379
rect 26525 30345 26559 30379
rect 2513 30277 2547 30311
rect 5917 30277 5951 30311
rect 10793 30277 10827 30311
rect 22109 30277 22143 30311
rect 35633 30277 35667 30311
rect 3525 30209 3559 30243
rect 7481 30209 7515 30243
rect 7849 30209 7883 30243
rect 11437 30209 11471 30243
rect 13185 30209 13219 30243
rect 16957 30209 16991 30243
rect 18061 30209 18095 30243
rect 18524 30209 18558 30243
rect 18797 30209 18831 30243
rect 33057 30209 33091 30243
rect 3341 30141 3375 30175
rect 4537 30141 4571 30175
rect 7205 30141 7239 30175
rect 8493 30141 8527 30175
rect 11161 30141 11195 30175
rect 11805 30141 11839 30175
rect 14013 30141 14047 30175
rect 14197 30141 14231 30175
rect 14453 30141 14487 30175
rect 16313 30141 16347 30175
rect 16773 30141 16807 30175
rect 20269 30141 20303 30175
rect 20729 30141 20763 30175
rect 23673 30141 23707 30175
rect 24225 30141 24259 30175
rect 24777 30141 24811 30175
rect 25033 30141 25067 30175
rect 26985 30141 27019 30175
rect 27537 30141 27571 30175
rect 35449 30141 35483 30175
rect 36001 30141 36035 30175
rect 2881 30073 2915 30107
rect 3433 30073 3467 30107
rect 4445 30073 4479 30107
rect 4782 30073 4816 30107
rect 6561 30073 6595 30107
rect 7297 30073 7331 30107
rect 8738 30073 8772 30107
rect 11253 30073 11287 30107
rect 12265 30073 12299 30107
rect 13093 30073 13127 30107
rect 17785 30073 17819 30107
rect 20974 30073 21008 30107
rect 23489 30073 23523 30107
rect 32873 30073 32907 30107
rect 6285 30005 6319 30039
rect 8401 30005 8435 30039
rect 10241 30005 10275 30039
rect 10701 30005 10735 30039
rect 12633 30005 12667 30039
rect 13001 30005 13035 30039
rect 15577 30005 15611 30039
rect 15853 30005 15887 30039
rect 16405 30005 16439 30039
rect 16865 30005 16899 30039
rect 17509 30005 17543 30039
rect 18527 30005 18561 30039
rect 19901 30005 19935 30039
rect 20545 30005 20579 30039
rect 23857 30005 23891 30039
rect 26157 30005 26191 30039
rect 27169 30005 27203 30039
rect 32229 30005 32263 30039
rect 32413 30005 32447 30039
rect 32781 30005 32815 30039
rect 35357 30005 35391 30039
rect 2329 29801 2363 29835
rect 2421 29801 2455 29835
rect 6009 29801 6043 29835
rect 7849 29801 7883 29835
rect 8861 29801 8895 29835
rect 11069 29801 11103 29835
rect 11437 29801 11471 29835
rect 14197 29801 14231 29835
rect 16135 29801 16169 29835
rect 17509 29801 17543 29835
rect 18521 29801 18555 29835
rect 22293 29801 22327 29835
rect 24961 29801 24995 29835
rect 25053 29801 25087 29835
rect 35909 29801 35943 29835
rect 4506 29733 4540 29767
rect 9934 29733 9968 29767
rect 13062 29733 13096 29767
rect 18153 29733 18187 29767
rect 24133 29733 24167 29767
rect 24409 29733 24443 29767
rect 2789 29665 2823 29699
rect 3893 29665 3927 29699
rect 4261 29665 4295 29699
rect 6725 29665 6759 29699
rect 8585 29665 8619 29699
rect 9689 29665 9723 29699
rect 14841 29665 14875 29699
rect 16405 29665 16439 29699
rect 19625 29665 19659 29699
rect 20913 29665 20947 29699
rect 21180 29665 21214 29699
rect 32505 29665 32539 29699
rect 33773 29665 33807 29699
rect 35725 29665 35759 29699
rect 2881 29597 2915 29631
rect 2973 29597 3007 29631
rect 6377 29597 6411 29631
rect 6469 29597 6503 29631
rect 8217 29597 8251 29631
rect 12173 29597 12207 29631
rect 12817 29597 12851 29631
rect 15577 29597 15611 29631
rect 15669 29597 15703 29631
rect 16175 29597 16209 29631
rect 19717 29597 19751 29631
rect 19809 29597 19843 29631
rect 25145 29597 25179 29631
rect 25605 29597 25639 29631
rect 26525 29597 26559 29631
rect 33517 29597 33551 29631
rect 5641 29529 5675 29563
rect 12541 29461 12575 29495
rect 14473 29461 14507 29495
rect 19165 29461 19199 29495
rect 19257 29461 19291 29495
rect 24593 29461 24627 29495
rect 27077 29461 27111 29495
rect 34897 29461 34931 29495
rect 35265 29461 35299 29495
rect 2513 29257 2547 29291
rect 4077 29257 4111 29291
rect 4445 29257 4479 29291
rect 5181 29257 5215 29291
rect 6561 29257 6595 29291
rect 9965 29257 9999 29291
rect 11345 29257 11379 29291
rect 11805 29257 11839 29291
rect 13461 29257 13495 29291
rect 15577 29257 15611 29291
rect 17049 29257 17083 29291
rect 17325 29257 17359 29291
rect 17785 29257 17819 29291
rect 18429 29257 18463 29291
rect 18889 29257 18923 29291
rect 21833 29257 21867 29291
rect 24593 29257 24627 29291
rect 26157 29257 26191 29291
rect 26433 29257 26467 29291
rect 26801 29257 26835 29291
rect 9781 29189 9815 29223
rect 12449 29189 12483 29223
rect 14013 29189 14047 29223
rect 19165 29189 19199 29223
rect 21189 29189 21223 29223
rect 23857 29189 23891 29223
rect 24317 29189 24351 29223
rect 26985 29189 27019 29223
rect 34897 29189 34931 29223
rect 5089 29121 5123 29155
rect 5641 29121 5675 29155
rect 5733 29121 5767 29155
rect 7113 29121 7147 29155
rect 7757 29121 7791 29155
rect 10609 29121 10643 29155
rect 13093 29121 13127 29155
rect 14565 29121 14599 29155
rect 15669 29121 15703 29155
rect 19812 29121 19846 29155
rect 20085 29121 20119 29155
rect 27537 29121 27571 29155
rect 35541 29121 35575 29155
rect 2697 29053 2731 29087
rect 5549 29053 5583 29087
rect 10333 29053 10367 29087
rect 10977 29053 11011 29087
rect 12817 29053 12851 29087
rect 15209 29053 15243 29087
rect 15936 29053 15970 29087
rect 19349 29053 19383 29087
rect 21465 29053 21499 29087
rect 23489 29053 23523 29087
rect 23673 29053 23707 29087
rect 24777 29053 24811 29087
rect 27353 29053 27387 29087
rect 31493 29053 31527 29087
rect 34345 29053 34379 29087
rect 35265 29053 35299 29087
rect 1777 28985 1811 29019
rect 2145 28985 2179 29019
rect 2942 28985 2976 29019
rect 7665 28985 7699 29019
rect 8002 28985 8036 29019
rect 12173 28985 12207 29019
rect 12909 28985 12943 29019
rect 13829 28985 13863 29019
rect 14381 28985 14415 29019
rect 22017 28985 22051 29019
rect 25022 28985 25056 29019
rect 27445 28985 27479 29019
rect 31738 28985 31772 29019
rect 35357 28985 35391 29019
rect 35909 28985 35943 29019
rect 9137 28917 9171 28951
rect 10425 28917 10459 28951
rect 14473 28917 14507 28951
rect 19815 28917 19849 28951
rect 31309 28917 31343 28951
rect 32873 28917 32907 28951
rect 33609 28917 33643 28951
rect 33977 28917 34011 28951
rect 34713 28917 34747 28951
rect 3157 28713 3191 28747
rect 3341 28713 3375 28747
rect 3525 28713 3559 28747
rect 3893 28713 3927 28747
rect 5457 28713 5491 28747
rect 5825 28713 5859 28747
rect 8493 28713 8527 28747
rect 9873 28713 9907 28747
rect 10609 28713 10643 28747
rect 13369 28713 13403 28747
rect 14105 28713 14139 28747
rect 15669 28713 15703 28747
rect 18797 28713 18831 28747
rect 19257 28713 19291 28747
rect 19625 28713 19659 28747
rect 20729 28713 20763 28747
rect 22293 28713 22327 28747
rect 23673 28713 23707 28747
rect 24133 28713 24167 28747
rect 31217 28713 31251 28747
rect 33793 28713 33827 28747
rect 36001 28713 36035 28747
rect 2044 28645 2078 28679
rect 1777 28509 1811 28543
rect 4322 28645 4356 28679
rect 11244 28645 11278 28679
rect 14381 28645 14415 28679
rect 15761 28645 15795 28679
rect 19073 28645 19107 28679
rect 24492 28645 24526 28679
rect 4077 28577 4111 28611
rect 8401 28577 8435 28611
rect 9689 28577 9723 28611
rect 13185 28577 13219 28611
rect 20913 28577 20947 28611
rect 21180 28577 21214 28611
rect 24225 28577 24259 28611
rect 26781 28577 26815 28611
rect 30093 28577 30127 28611
rect 32669 28577 32703 28611
rect 34877 28577 34911 28611
rect 7481 28509 7515 28543
rect 8677 28509 8711 28543
rect 9505 28509 9539 28543
rect 10977 28509 11011 28543
rect 15853 28509 15887 28543
rect 16865 28509 16899 28543
rect 19717 28509 19751 28543
rect 19809 28509 19843 28543
rect 23213 28509 23247 28543
rect 26525 28509 26559 28543
rect 29745 28509 29779 28543
rect 29837 28509 29871 28543
rect 32413 28509 32447 28543
rect 34621 28509 34655 28543
rect 8033 28441 8067 28475
rect 10241 28441 10275 28475
rect 15301 28441 15335 28475
rect 25881 28441 25915 28475
rect 3341 28373 3375 28407
rect 7849 28373 7883 28407
rect 12357 28373 12391 28407
rect 12633 28373 12667 28407
rect 13001 28373 13035 28407
rect 15117 28373 15151 28407
rect 16313 28373 16347 28407
rect 20361 28373 20395 28407
rect 25605 28373 25639 28407
rect 27905 28373 27939 28407
rect 31585 28373 31619 28407
rect 34437 28373 34471 28407
rect 1869 28169 1903 28203
rect 4169 28169 4203 28203
rect 4537 28169 4571 28203
rect 7297 28169 7331 28203
rect 8769 28169 8803 28203
rect 9873 28169 9907 28203
rect 11897 28169 11931 28203
rect 12265 28169 12299 28203
rect 13461 28169 13495 28203
rect 14657 28169 14691 28203
rect 15301 28169 15335 28203
rect 15485 28169 15519 28203
rect 16497 28169 16531 28203
rect 19349 28169 19383 28203
rect 20085 28169 20119 28203
rect 23857 28169 23891 28203
rect 27261 28169 27295 28203
rect 29653 28169 29687 28203
rect 31493 28169 31527 28203
rect 32229 28169 32263 28203
rect 34713 28169 34747 28203
rect 9597 28101 9631 28135
rect 10793 28101 10827 28135
rect 12449 28101 12483 28135
rect 18981 28101 19015 28135
rect 24041 28101 24075 28135
rect 8401 28033 8435 28067
rect 10701 28033 10735 28067
rect 11253 28033 11287 28067
rect 11345 28033 11379 28067
rect 12909 28033 12943 28067
rect 13001 28033 13035 28067
rect 15945 28033 15979 28067
rect 16129 28033 16163 28067
rect 16313 28033 16347 28067
rect 19625 28033 19659 28067
rect 23489 28033 23523 28067
rect 24685 28033 24719 28067
rect 25513 28033 25547 28067
rect 31953 28033 31987 28067
rect 32965 28033 32999 28067
rect 8217 27965 8251 27999
rect 9689 27965 9723 27999
rect 12817 27965 12851 27999
rect 15853 27965 15887 27999
rect 20729 27965 20763 27999
rect 24409 27965 24443 27999
rect 25605 27965 25639 27999
rect 25872 27965 25906 27999
rect 29101 27965 29135 27999
rect 30113 27965 30147 27999
rect 34989 27965 35023 27999
rect 35256 27965 35290 27999
rect 8125 27897 8159 27931
rect 15025 27897 15059 27931
rect 16313 27897 16347 27931
rect 20996 27897 21030 27931
rect 22385 27897 22419 27931
rect 25145 27897 25179 27931
rect 30021 27897 30055 27931
rect 30358 27897 30392 27931
rect 31861 27897 31895 27931
rect 31953 27897 31987 27931
rect 32781 27897 32815 27931
rect 36645 27897 36679 27931
rect 2145 27829 2179 27863
rect 7573 27829 7607 27863
rect 7757 27829 7791 27863
rect 9229 27829 9263 27863
rect 10241 27829 10275 27863
rect 11161 27829 11195 27863
rect 20637 27829 20671 27863
rect 22109 27829 22143 27863
rect 24501 27829 24535 27863
rect 26985 27829 27019 27863
rect 32321 27829 32355 27863
rect 32689 27829 32723 27863
rect 33333 27829 33367 27863
rect 33793 27829 33827 27863
rect 34161 27829 34195 27863
rect 36369 27829 36403 27863
rect 2789 27625 2823 27659
rect 8585 27625 8619 27659
rect 9505 27625 9539 27659
rect 15577 27625 15611 27659
rect 15853 27625 15887 27659
rect 21925 27625 21959 27659
rect 23765 27625 23799 27659
rect 24869 27625 24903 27659
rect 31033 27625 31067 27659
rect 32597 27625 32631 27659
rect 35081 27625 35115 27659
rect 10885 27557 10919 27591
rect 21281 27557 21315 27591
rect 24133 27557 24167 27591
rect 25237 27557 25271 27591
rect 31953 27557 31987 27591
rect 32505 27557 32539 27591
rect 1409 27489 1443 27523
rect 1676 27489 1710 27523
rect 7205 27489 7239 27523
rect 7461 27489 7495 27523
rect 9965 27489 9999 27523
rect 11069 27489 11103 27523
rect 11336 27489 11370 27523
rect 13277 27489 13311 27523
rect 16497 27489 16531 27523
rect 19625 27489 19659 27523
rect 22845 27489 22879 27523
rect 29561 27489 29595 27523
rect 29653 27489 29687 27523
rect 29920 27489 29954 27523
rect 31585 27489 31619 27523
rect 34069 27489 34103 27523
rect 35440 27489 35474 27523
rect 19717 27421 19751 27455
rect 19901 27421 19935 27455
rect 20729 27421 20763 27455
rect 21373 27421 21407 27455
rect 21557 27421 21591 27455
rect 22937 27421 22971 27455
rect 23121 27421 23155 27455
rect 25329 27421 25363 27455
rect 25421 27421 25455 27455
rect 26525 27421 26559 27455
rect 32781 27421 32815 27455
rect 35173 27421 35207 27455
rect 10149 27353 10183 27387
rect 13461 27353 13495 27387
rect 19257 27353 19291 27387
rect 20913 27353 20947 27387
rect 22477 27353 22511 27387
rect 24777 27353 24811 27387
rect 34621 27353 34655 27387
rect 12449 27285 12483 27319
rect 12817 27285 12851 27319
rect 16221 27285 16255 27319
rect 16681 27285 16715 27319
rect 20361 27285 20395 27319
rect 25881 27285 25915 27319
rect 26985 27285 27019 27319
rect 32137 27285 32171 27319
rect 33241 27285 33275 27319
rect 34253 27285 34287 27319
rect 36553 27285 36587 27319
rect 36829 27285 36863 27319
rect 2053 27081 2087 27115
rect 6653 27081 6687 27115
rect 7757 27081 7791 27115
rect 8217 27081 8251 27115
rect 9965 27081 9999 27115
rect 10701 27081 10735 27115
rect 11805 27081 11839 27115
rect 12449 27081 12483 27115
rect 13461 27081 13495 27115
rect 15301 27081 15335 27115
rect 17141 27081 17175 27115
rect 18981 27081 19015 27115
rect 19349 27081 19383 27115
rect 20361 27081 20395 27115
rect 21833 27081 21867 27115
rect 23213 27081 23247 27115
rect 25421 27081 25455 27115
rect 27813 27081 27847 27115
rect 30849 27081 30883 27115
rect 31125 27081 31159 27115
rect 31493 27081 31527 27115
rect 31677 27081 31711 27115
rect 32689 27081 32723 27115
rect 34345 27081 34379 27115
rect 34713 27081 34747 27115
rect 36001 27081 36035 27115
rect 36369 27081 36403 27115
rect 37473 27081 37507 27115
rect 22109 27013 22143 27047
rect 8861 26945 8895 26979
rect 11345 26945 11379 26979
rect 13001 26945 13035 26979
rect 19441 26945 19475 26979
rect 24593 26945 24627 26979
rect 28733 26945 28767 26979
rect 32137 26945 32171 26979
rect 32321 26945 32355 26979
rect 33793 26945 33827 26979
rect 35357 26945 35391 26979
rect 35449 26945 35483 26979
rect 37013 26945 37047 26979
rect 8585 26877 8619 26911
rect 9689 26877 9723 26911
rect 12909 26877 12943 26911
rect 14381 26877 14415 26911
rect 15393 26877 15427 26911
rect 15649 26877 15683 26911
rect 20453 26877 20487 26911
rect 24501 26877 24535 26911
rect 25605 26877 25639 26911
rect 27997 26877 28031 26911
rect 28273 26877 28307 26911
rect 29469 26877 29503 26911
rect 33609 26877 33643 26911
rect 36921 26877 36955 26911
rect 1685 26809 1719 26843
rect 8677 26809 8711 26843
rect 10609 26809 10643 26843
rect 11161 26809 11195 26843
rect 19993 26809 20027 26843
rect 20720 26809 20754 26843
rect 22845 26809 22879 26843
rect 23949 26809 23983 26843
rect 25145 26809 25179 26843
rect 25872 26809 25906 26843
rect 29101 26809 29135 26843
rect 29714 26809 29748 26843
rect 33701 26809 33735 26843
rect 35265 26809 35299 26843
rect 7297 26741 7331 26775
rect 8033 26741 8067 26775
rect 11069 26741 11103 26775
rect 12173 26741 12207 26775
rect 12817 26741 12851 26775
rect 14197 26741 14231 26775
rect 14749 26741 14783 26775
rect 16773 26741 16807 26775
rect 22569 26741 22603 26775
rect 24041 26741 24075 26775
rect 24409 26741 24443 26775
rect 26985 26741 27019 26775
rect 32045 26741 32079 26775
rect 33057 26741 33091 26775
rect 33241 26741 33275 26775
rect 34897 26741 34931 26775
rect 36461 26741 36495 26775
rect 36829 26741 36863 26775
rect 8309 26537 8343 26571
rect 8677 26537 8711 26571
rect 10425 26537 10459 26571
rect 15945 26537 15979 26571
rect 19257 26537 19291 26571
rect 19625 26537 19659 26571
rect 20545 26537 20579 26571
rect 22293 26537 22327 26571
rect 23857 26537 23891 26571
rect 24869 26537 24903 26571
rect 25237 26537 25271 26571
rect 30849 26537 30883 26571
rect 31677 26537 31711 26571
rect 32137 26537 32171 26571
rect 34989 26537 35023 26571
rect 7174 26469 7208 26503
rect 10793 26469 10827 26503
rect 19165 26469 19199 26503
rect 24777 26469 24811 26503
rect 32505 26469 32539 26503
rect 34161 26469 34195 26503
rect 11336 26401 11370 26435
rect 15853 26401 15887 26435
rect 17049 26401 17083 26435
rect 18797 26401 18831 26435
rect 21169 26401 21203 26435
rect 27261 26401 27295 26435
rect 29725 26401 29759 26435
rect 33517 26401 33551 26435
rect 34069 26401 34103 26435
rect 35521 26401 35555 26435
rect 6929 26333 6963 26367
rect 11069 26333 11103 26367
rect 15117 26333 15151 26367
rect 16129 26333 16163 26367
rect 19717 26333 19751 26367
rect 19809 26333 19843 26367
rect 20913 26333 20947 26367
rect 25329 26333 25363 26367
rect 25513 26333 25547 26367
rect 26249 26333 26283 26367
rect 26525 26333 26559 26367
rect 26848 26333 26882 26367
rect 26988 26333 27022 26367
rect 29377 26333 29411 26367
rect 29469 26333 29503 26367
rect 31309 26333 31343 26367
rect 32597 26333 32631 26367
rect 32781 26333 32815 26367
rect 34253 26333 34287 26367
rect 35265 26333 35299 26367
rect 12449 26265 12483 26299
rect 12725 26265 12759 26299
rect 15485 26265 15519 26299
rect 17233 26265 17267 26299
rect 24225 26265 24259 26299
rect 25973 26265 26007 26299
rect 28365 26265 28399 26299
rect 29009 26265 29043 26299
rect 36645 26265 36679 26299
rect 36921 26265 36955 26299
rect 33149 26197 33183 26231
rect 33701 26197 33735 26231
rect 6653 25993 6687 26027
rect 8309 25993 8343 26027
rect 11805 25993 11839 26027
rect 12449 25993 12483 26027
rect 17049 25993 17083 26027
rect 20729 25993 20763 26027
rect 22661 25993 22695 26027
rect 26801 25993 26835 26027
rect 28181 25993 28215 26027
rect 28733 25993 28767 26027
rect 30849 25993 30883 26027
rect 31217 25993 31251 26027
rect 31585 25993 31619 26027
rect 32321 25993 32355 26027
rect 32689 25993 32723 26027
rect 34713 25993 34747 26027
rect 36093 25993 36127 26027
rect 19349 25925 19383 25959
rect 25973 25925 26007 25959
rect 31861 25925 31895 25959
rect 10057 25857 10091 25891
rect 13001 25857 13035 25891
rect 14841 25857 14875 25891
rect 15209 25857 15243 25891
rect 20361 25857 20395 25891
rect 21327 25857 21361 25891
rect 23489 25857 23523 25891
rect 24596 25857 24630 25891
rect 24869 25857 24903 25891
rect 27445 25857 27479 25891
rect 29469 25857 29503 25891
rect 33425 25857 33459 25891
rect 6285 25789 6319 25823
rect 6929 25789 6963 25823
rect 8677 25789 8711 25823
rect 9689 25789 9723 25823
rect 10149 25789 10183 25823
rect 10416 25789 10450 25823
rect 14105 25789 14139 25823
rect 14473 25789 14507 25823
rect 15301 25789 15335 25823
rect 15568 25789 15602 25823
rect 18061 25789 18095 25823
rect 18613 25789 18647 25823
rect 19165 25789 19199 25823
rect 20821 25789 20855 25823
rect 21557 25789 21591 25823
rect 24133 25789 24167 25823
rect 27261 25789 27295 25823
rect 31677 25789 31711 25823
rect 33149 25789 33183 25823
rect 35357 25789 35391 25823
rect 35633 25789 35667 25823
rect 35817 25789 35851 25823
rect 36645 25789 36679 25823
rect 37197 25789 37231 25823
rect 7174 25721 7208 25755
rect 12909 25721 12943 25755
rect 19809 25721 19843 25755
rect 27169 25721 27203 25755
rect 27813 25721 27847 25755
rect 29101 25721 29135 25755
rect 29714 25721 29748 25755
rect 35449 25721 35483 25755
rect 11529 25653 11563 25687
rect 12173 25653 12207 25687
rect 12817 25653 12851 25687
rect 16681 25653 16715 25687
rect 18245 25653 18279 25687
rect 19073 25653 19107 25687
rect 21287 25653 21321 25687
rect 24041 25653 24075 25687
rect 24599 25653 24633 25687
rect 26617 25653 26651 25687
rect 32781 25653 32815 25687
rect 33241 25653 33275 25687
rect 33793 25653 33827 25687
rect 34161 25653 34195 25687
rect 36461 25653 36495 25687
rect 36829 25653 36863 25687
rect 10609 25449 10643 25483
rect 12541 25449 12575 25483
rect 19257 25449 19291 25483
rect 20729 25449 20763 25483
rect 21097 25449 21131 25483
rect 21557 25449 21591 25483
rect 23673 25449 23707 25483
rect 25881 25449 25915 25483
rect 26249 25449 26283 25483
rect 26893 25449 26927 25483
rect 27537 25449 27571 25483
rect 29285 25449 29319 25483
rect 30757 25449 30791 25483
rect 32505 25449 32539 25483
rect 34437 25449 34471 25483
rect 14013 25381 14047 25415
rect 20361 25381 20395 25415
rect 21833 25381 21867 25415
rect 24133 25381 24167 25415
rect 24492 25381 24526 25415
rect 27169 25381 27203 25415
rect 33333 25381 33367 25415
rect 35256 25381 35290 25415
rect 7113 25313 7147 25347
rect 7369 25313 7403 25347
rect 10957 25313 10991 25347
rect 15557 25313 15591 25347
rect 18153 25313 18187 25347
rect 19625 25313 19659 25347
rect 19717 25313 19751 25347
rect 20913 25313 20947 25347
rect 28181 25313 28215 25347
rect 28273 25313 28307 25347
rect 29633 25313 29667 25347
rect 31769 25313 31803 25347
rect 32321 25313 32355 25347
rect 33793 25313 33827 25347
rect 10701 25245 10735 25279
rect 14105 25245 14139 25279
rect 14289 25245 14323 25279
rect 15301 25245 15335 25279
rect 16957 25245 16991 25279
rect 19165 25245 19199 25279
rect 19809 25245 19843 25279
rect 23213 25245 23247 25279
rect 24225 25245 24259 25279
rect 28457 25245 28491 25279
rect 29377 25245 29411 25279
rect 33885 25245 33919 25279
rect 34069 25245 34103 25279
rect 34989 25245 35023 25279
rect 31585 25177 31619 25211
rect 7021 25109 7055 25143
rect 8493 25109 8527 25143
rect 10149 25109 10183 25143
rect 12081 25109 12115 25143
rect 12909 25109 12943 25143
rect 13645 25109 13679 25143
rect 14749 25109 14783 25143
rect 15025 25109 15059 25143
rect 16681 25109 16715 25143
rect 17417 25109 17451 25143
rect 18337 25109 18371 25143
rect 18705 25109 18739 25143
rect 25605 25109 25639 25143
rect 27813 25109 27847 25143
rect 32873 25109 32907 25143
rect 33425 25109 33459 25143
rect 34805 25109 34839 25143
rect 36369 25109 36403 25143
rect 6653 24905 6687 24939
rect 9689 24905 9723 24939
rect 10057 24905 10091 24939
rect 12449 24905 12483 24939
rect 14749 24905 14783 24939
rect 18337 24905 18371 24939
rect 19809 24905 19843 24939
rect 21281 24905 21315 24939
rect 23489 24905 23523 24939
rect 24225 24905 24259 24939
rect 27537 24905 27571 24939
rect 30665 24905 30699 24939
rect 32505 24905 32539 24939
rect 33149 24905 33183 24939
rect 33885 24905 33919 24939
rect 34713 24905 34747 24939
rect 36369 24905 36403 24939
rect 36645 24905 36679 24939
rect 17049 24837 17083 24871
rect 21557 24837 21591 24871
rect 31033 24837 31067 24871
rect 11897 24769 11931 24803
rect 13001 24769 13035 24803
rect 13737 24769 13771 24803
rect 16589 24769 16623 24803
rect 16957 24769 16991 24803
rect 18981 24769 19015 24803
rect 21925 24769 21959 24803
rect 23949 24769 23983 24803
rect 28733 24769 28767 24803
rect 31401 24769 31435 24803
rect 31953 24769 31987 24803
rect 32045 24769 32079 24803
rect 34253 24769 34287 24803
rect 35541 24769 35575 24803
rect 37105 24769 37139 24803
rect 7389 24701 7423 24735
rect 10149 24701 10183 24735
rect 14841 24701 14875 24735
rect 17233 24701 17267 24735
rect 19901 24701 19935 24735
rect 20157 24701 20191 24735
rect 24501 24701 24535 24735
rect 24757 24701 24791 24735
rect 29285 24701 29319 24735
rect 33609 24701 33643 24735
rect 33701 24701 33735 24735
rect 35265 24701 35299 24735
rect 36461 24701 36495 24735
rect 7297 24633 7331 24667
rect 7656 24633 7690 24667
rect 10394 24633 10428 24667
rect 12909 24633 12943 24667
rect 15108 24633 15142 24667
rect 18797 24633 18831 24667
rect 19441 24633 19475 24667
rect 22109 24633 22143 24667
rect 26249 24633 26283 24667
rect 27905 24633 27939 24667
rect 29101 24633 29135 24667
rect 29530 24633 29564 24667
rect 35357 24633 35391 24667
rect 35909 24633 35943 24667
rect 8769 24565 8803 24599
rect 11529 24565 11563 24599
rect 12173 24565 12207 24599
rect 12817 24565 12851 24599
rect 14105 24565 14139 24599
rect 16221 24565 16255 24599
rect 17785 24565 17819 24599
rect 18705 24565 18739 24599
rect 25881 24565 25915 24599
rect 28273 24565 28307 24599
rect 31493 24565 31527 24599
rect 31861 24565 31895 24599
rect 34897 24565 34931 24599
rect 7205 24361 7239 24395
rect 7849 24361 7883 24395
rect 10241 24361 10275 24395
rect 11989 24361 12023 24395
rect 15301 24361 15335 24395
rect 15669 24361 15703 24395
rect 15761 24361 15795 24395
rect 16865 24361 16899 24395
rect 18061 24361 18095 24395
rect 19993 24361 20027 24395
rect 20269 24361 20303 24395
rect 20913 24361 20947 24395
rect 24317 24361 24351 24395
rect 27261 24361 27295 24395
rect 29193 24361 29227 24395
rect 30665 24361 30699 24395
rect 31493 24361 31527 24395
rect 31953 24361 31987 24395
rect 32321 24361 32355 24395
rect 33517 24361 33551 24395
rect 33885 24361 33919 24395
rect 36645 24361 36679 24395
rect 8309 24293 8343 24327
rect 12541 24293 12575 24327
rect 14933 24293 14967 24327
rect 18337 24293 18371 24327
rect 20637 24293 20671 24327
rect 21281 24293 21315 24327
rect 24685 24293 24719 24327
rect 34520 24293 34554 24327
rect 8217 24225 8251 24259
rect 10865 24225 10899 24259
rect 14105 24225 14139 24259
rect 17233 24225 17267 24259
rect 18880 24225 18914 24259
rect 24777 24225 24811 24259
rect 27445 24225 27479 24259
rect 29552 24225 29586 24259
rect 32137 24225 32171 24259
rect 34253 24225 34287 24259
rect 36461 24225 36495 24259
rect 8493 24157 8527 24191
rect 10609 24157 10643 24191
rect 15853 24157 15887 24191
rect 17325 24157 17359 24191
rect 17509 24157 17543 24191
rect 18613 24157 18647 24191
rect 21373 24157 21407 24191
rect 21465 24157 21499 24191
rect 24869 24157 24903 24191
rect 29285 24157 29319 24191
rect 7573 24089 7607 24123
rect 14289 24089 14323 24123
rect 16497 24089 16531 24123
rect 13737 24021 13771 24055
rect 25329 24021 25363 24055
rect 35633 24021 35667 24055
rect 7941 23817 7975 23851
rect 8217 23817 8251 23851
rect 8585 23817 8619 23851
rect 10701 23817 10735 23851
rect 11345 23817 11379 23851
rect 13277 23817 13311 23851
rect 15393 23817 15427 23851
rect 15761 23817 15795 23851
rect 16405 23817 16439 23851
rect 17417 23817 17451 23851
rect 17785 23817 17819 23851
rect 18245 23817 18279 23851
rect 19625 23817 19659 23851
rect 19993 23817 20027 23851
rect 20729 23817 20763 23851
rect 22109 23817 22143 23851
rect 24133 23817 24167 23851
rect 24685 23817 24719 23851
rect 27353 23817 27387 23851
rect 28733 23817 28767 23851
rect 28917 23817 28951 23851
rect 29561 23817 29595 23851
rect 31309 23817 31343 23851
rect 32137 23817 32171 23851
rect 32781 23817 32815 23851
rect 33149 23817 33183 23851
rect 33517 23817 33551 23851
rect 33885 23817 33919 23851
rect 35909 23817 35943 23851
rect 36461 23817 36495 23851
rect 11069 23749 11103 23783
rect 15945 23749 15979 23783
rect 20269 23749 20303 23783
rect 26433 23749 26467 23783
rect 29929 23749 29963 23783
rect 30941 23749 30975 23783
rect 13645 23681 13679 23715
rect 17049 23681 17083 23715
rect 23489 23681 23523 23715
rect 30389 23681 30423 23715
rect 30573 23681 30607 23715
rect 34345 23681 34379 23715
rect 35541 23681 35575 23715
rect 11529 23613 11563 23647
rect 11805 23613 11839 23647
rect 12909 23613 12943 23647
rect 13737 23613 13771 23647
rect 14004 23613 14038 23647
rect 16129 23613 16163 23647
rect 18061 23613 18095 23647
rect 18613 23613 18647 23647
rect 19165 23613 19199 23647
rect 19441 23613 19475 23647
rect 24869 23613 24903 23647
rect 25145 23613 25179 23647
rect 25421 23613 25455 23647
rect 25973 23613 26007 23647
rect 29101 23613 29135 23647
rect 32597 23613 32631 23647
rect 33701 23613 33735 23647
rect 35357 23613 35391 23647
rect 16773 23545 16807 23579
rect 19257 23545 19291 23579
rect 20821 23545 20855 23579
rect 24593 23545 24627 23579
rect 24961 23545 24995 23579
rect 25329 23545 25363 23579
rect 30297 23545 30331 23579
rect 34713 23545 34747 23579
rect 35265 23545 35299 23579
rect 15117 23477 15151 23511
rect 16865 23477 16899 23511
rect 25605 23477 25639 23511
rect 28457 23477 28491 23511
rect 34897 23477 34931 23511
rect 10425 23273 10459 23307
rect 12541 23273 12575 23307
rect 15117 23273 15151 23307
rect 15301 23273 15335 23307
rect 18797 23273 18831 23307
rect 20545 23273 20579 23307
rect 21189 23273 21223 23307
rect 28089 23273 28123 23307
rect 30297 23273 30331 23307
rect 30573 23273 30607 23307
rect 34069 23273 34103 23307
rect 35817 23273 35851 23307
rect 36369 23273 36403 23307
rect 19432 23205 19466 23239
rect 24952 23205 24986 23239
rect 33701 23205 33735 23239
rect 34428 23205 34462 23239
rect 10609 23137 10643 23171
rect 12725 23137 12759 23171
rect 13268 23137 13302 23171
rect 15669 23137 15703 23171
rect 17233 23137 17267 23171
rect 19165 23137 19199 23171
rect 24685 23137 24719 23171
rect 28273 23137 28307 23171
rect 29184 23137 29218 23171
rect 33057 23137 33091 23171
rect 13001 23069 13035 23103
rect 15761 23069 15795 23103
rect 15945 23069 15979 23103
rect 17325 23069 17359 23103
rect 17417 23069 17451 23103
rect 17877 23069 17911 23103
rect 28917 23069 28951 23103
rect 34161 23069 34195 23103
rect 14749 23001 14783 23035
rect 12449 22933 12483 22967
rect 14381 22933 14415 22967
rect 16405 22933 16439 22967
rect 16865 22933 16899 22967
rect 18429 22933 18463 22967
rect 21557 22933 21591 22967
rect 22109 22933 22143 22967
rect 24317 22933 24351 22967
rect 26065 22933 26099 22967
rect 33241 22933 33275 22967
rect 35541 22933 35575 22967
rect 10517 22729 10551 22763
rect 12265 22729 12299 22763
rect 13001 22729 13035 22763
rect 13921 22729 13955 22763
rect 15393 22729 15427 22763
rect 16497 22729 16531 22763
rect 17325 22729 17359 22763
rect 17601 22729 17635 22763
rect 19717 22729 19751 22763
rect 19993 22729 20027 22763
rect 20821 22729 20855 22763
rect 23949 22729 23983 22763
rect 25697 22729 25731 22763
rect 30757 22729 30791 22763
rect 31217 22729 31251 22763
rect 31769 22729 31803 22763
rect 32781 22729 32815 22763
rect 34345 22729 34379 22763
rect 12725 22661 12759 22695
rect 15485 22661 15519 22695
rect 13461 22593 13495 22627
rect 13829 22593 13863 22627
rect 14381 22593 14415 22627
rect 14565 22593 14599 22627
rect 16037 22593 16071 22627
rect 21557 22593 21591 22627
rect 22661 22593 22695 22627
rect 29929 22593 29963 22627
rect 30297 22593 30331 22627
rect 32413 22593 32447 22627
rect 33793 22593 33827 22627
rect 34621 22593 34655 22627
rect 12817 22525 12851 22559
rect 18337 22525 18371 22559
rect 18593 22525 18627 22559
rect 22385 22525 22419 22559
rect 26893 22525 26927 22559
rect 27445 22525 27479 22559
rect 28733 22525 28767 22559
rect 31401 22525 31435 22559
rect 33149 22525 33183 22559
rect 33701 22525 33735 22559
rect 34897 22525 34931 22559
rect 35153 22525 35187 22559
rect 15853 22457 15887 22491
rect 16865 22457 16899 22491
rect 21925 22457 21959 22491
rect 24409 22457 24443 22491
rect 29101 22457 29135 22491
rect 29653 22457 29687 22491
rect 33609 22457 33643 22491
rect 36553 22457 36587 22491
rect 14289 22389 14323 22423
rect 14933 22389 14967 22423
rect 15945 22389 15979 22423
rect 20361 22389 20395 22423
rect 22017 22389 22051 22423
rect 22477 22389 22511 22423
rect 24225 22389 24259 22423
rect 27077 22389 27111 22423
rect 28089 22389 28123 22423
rect 29285 22389 29319 22423
rect 29745 22389 29779 22423
rect 33241 22389 33275 22423
rect 36277 22389 36311 22423
rect 12633 22185 12667 22219
rect 14657 22185 14691 22219
rect 15025 22185 15059 22219
rect 15301 22185 15335 22219
rect 16865 22185 16899 22219
rect 18429 22185 18463 22219
rect 18797 22185 18831 22219
rect 19901 22185 19935 22219
rect 24869 22185 24903 22219
rect 29101 22185 29135 22219
rect 33241 22185 33275 22219
rect 34253 22185 34287 22219
rect 34529 22185 34563 22219
rect 34621 22185 34655 22219
rect 27629 22117 27663 22151
rect 30205 22117 30239 22151
rect 12817 22049 12851 22083
rect 13176 22049 13210 22083
rect 15669 22049 15703 22083
rect 17233 22049 17267 22083
rect 21169 22049 21203 22083
rect 23745 22049 23779 22083
rect 26525 22049 26559 22083
rect 28549 22049 28583 22083
rect 29009 22049 29043 22083
rect 29745 22049 29779 22083
rect 33609 22049 33643 22083
rect 35072 22049 35106 22083
rect 12909 21981 12943 22015
rect 15761 21981 15795 22015
rect 15853 21981 15887 22015
rect 17325 21981 17359 22015
rect 17509 21981 17543 22015
rect 18153 21981 18187 22015
rect 18889 21981 18923 22015
rect 19073 21981 19107 22015
rect 19441 21981 19475 22015
rect 20913 21981 20947 22015
rect 23489 21981 23523 22015
rect 29193 21981 29227 22015
rect 33701 21981 33735 22015
rect 33885 21981 33919 22015
rect 34529 21981 34563 22015
rect 34805 21981 34839 22015
rect 14289 21913 14323 21947
rect 16773 21913 16807 21947
rect 12541 21845 12575 21879
rect 16313 21845 16347 21879
rect 22293 21845 22327 21879
rect 25237 21845 25271 21879
rect 25605 21845 25639 21879
rect 26709 21845 26743 21879
rect 28641 21845 28675 21879
rect 30113 21845 30147 21879
rect 31493 21845 31527 21879
rect 33149 21845 33183 21879
rect 36185 21845 36219 21879
rect 11805 21641 11839 21675
rect 12909 21641 12943 21675
rect 14381 21641 14415 21675
rect 14749 21641 14783 21675
rect 15117 21641 15151 21675
rect 15209 21641 15243 21675
rect 16681 21641 16715 21675
rect 16957 21641 16991 21675
rect 17693 21641 17727 21675
rect 19441 21641 19475 21675
rect 20085 21641 20119 21675
rect 22753 21641 22787 21675
rect 23121 21641 23155 21675
rect 23857 21641 23891 21675
rect 24041 21641 24075 21675
rect 27261 21641 27295 21675
rect 28457 21641 28491 21675
rect 28825 21641 28859 21675
rect 30665 21641 30699 21675
rect 32781 21641 32815 21675
rect 34345 21641 34379 21675
rect 34713 21641 34747 21675
rect 36645 21641 36679 21675
rect 31493 21573 31527 21607
rect 12265 21505 12299 21539
rect 15853 21505 15887 21539
rect 24501 21505 24535 21539
rect 24685 21505 24719 21539
rect 32045 21505 32079 21539
rect 33793 21505 33827 21539
rect 13001 21437 13035 21471
rect 13268 21437 13302 21471
rect 16773 21437 16807 21471
rect 18061 21437 18095 21471
rect 21373 21437 21407 21471
rect 21640 21437 21674 21471
rect 25605 21437 25639 21471
rect 27813 21437 27847 21471
rect 29285 21437 29319 21471
rect 29552 21437 29586 21471
rect 31401 21437 31435 21471
rect 31861 21437 31895 21471
rect 33609 21437 33643 21471
rect 34989 21437 35023 21471
rect 35245 21437 35279 21471
rect 15577 21369 15611 21403
rect 16221 21369 16255 21403
rect 18328 21369 18362 21403
rect 20637 21369 20671 21403
rect 25850 21369 25884 21403
rect 27721 21369 27755 21403
rect 31033 21369 31067 21403
rect 33149 21369 33183 21403
rect 15669 21301 15703 21335
rect 17325 21301 17359 21335
rect 19717 21301 19751 21335
rect 20913 21301 20947 21335
rect 23489 21301 23523 21335
rect 24409 21301 24443 21335
rect 25421 21301 25455 21335
rect 26985 21301 27019 21335
rect 27997 21301 28031 21335
rect 31953 21301 31987 21335
rect 33241 21301 33275 21335
rect 33701 21301 33735 21335
rect 36369 21301 36403 21335
rect 12725 21097 12759 21131
rect 14381 21097 14415 21131
rect 15577 21097 15611 21131
rect 15945 21097 15979 21131
rect 17601 21097 17635 21131
rect 18061 21097 18095 21131
rect 23673 21097 23707 21131
rect 24133 21097 24167 21131
rect 25237 21097 25271 21131
rect 25329 21097 25363 21131
rect 29285 21097 29319 21131
rect 31033 21097 31067 21131
rect 31585 21097 31619 21131
rect 32137 21097 32171 21131
rect 32965 21097 32999 21131
rect 33333 21097 33367 21131
rect 35357 21097 35391 21131
rect 35633 21097 35667 21131
rect 13268 21029 13302 21063
rect 15117 21029 15151 21063
rect 22560 21029 22594 21063
rect 28733 21029 28767 21063
rect 29920 21029 29954 21063
rect 36185 21029 36219 21063
rect 16488 20961 16522 20995
rect 18429 20961 18463 20995
rect 21189 20961 21223 20995
rect 22201 20961 22235 20995
rect 22293 20961 22327 20995
rect 24501 20961 24535 20995
rect 27068 20961 27102 20995
rect 34253 20961 34287 20995
rect 13001 20893 13035 20927
rect 16221 20893 16255 20927
rect 20177 20893 20211 20927
rect 20545 20893 20579 20927
rect 21741 20893 21775 20927
rect 25421 20893 25455 20927
rect 26801 20893 26835 20927
rect 29653 20893 29687 20927
rect 33517 20893 33551 20927
rect 33840 20893 33874 20927
rect 33980 20893 34014 20927
rect 21373 20757 21407 20791
rect 24869 20757 24903 20791
rect 26065 20757 26099 20791
rect 28181 20757 28215 20791
rect 13369 20553 13403 20587
rect 15301 20553 15335 20587
rect 16129 20553 16163 20587
rect 17693 20553 17727 20587
rect 19441 20553 19475 20587
rect 21925 20553 21959 20587
rect 22385 20553 22419 20587
rect 24961 20553 24995 20587
rect 25329 20553 25363 20587
rect 27629 20553 27663 20587
rect 31401 20553 31435 20587
rect 31585 20553 31619 20587
rect 33701 20553 33735 20587
rect 33977 20553 34011 20587
rect 34345 20553 34379 20587
rect 13093 20485 13127 20519
rect 17233 20485 17267 20519
rect 19533 20485 19567 20519
rect 13829 20417 13863 20451
rect 16681 20417 16715 20451
rect 18061 20417 18095 20451
rect 20085 20417 20119 20451
rect 23121 20417 23155 20451
rect 24317 20417 24351 20451
rect 26525 20417 26559 20451
rect 26617 20417 26651 20451
rect 27077 20417 27111 20451
rect 28273 20417 28307 20451
rect 29748 20417 29782 20451
rect 13921 20349 13955 20383
rect 14188 20349 14222 20383
rect 17877 20349 17911 20383
rect 18317 20349 18351 20383
rect 19901 20349 19935 20383
rect 20545 20349 20579 20383
rect 24041 20349 24075 20383
rect 25973 20349 26007 20383
rect 26433 20349 26467 20383
rect 28733 20349 28767 20383
rect 29285 20349 29319 20383
rect 30021 20349 30055 20383
rect 16037 20281 16071 20315
rect 16589 20281 16623 20315
rect 20790 20281 20824 20315
rect 22753 20281 22787 20315
rect 24133 20281 24167 20315
rect 27537 20281 27571 20315
rect 27997 20281 28031 20315
rect 31960 20417 31994 20451
rect 35081 20349 35115 20383
rect 35348 20349 35382 20383
rect 31769 20281 31803 20315
rect 32198 20281 32232 20315
rect 36737 20281 36771 20315
rect 15669 20213 15703 20247
rect 16497 20213 16531 20247
rect 17509 20213 17543 20247
rect 19993 20213 20027 20247
rect 23489 20213 23523 20247
rect 23673 20213 23707 20247
rect 26065 20213 26099 20247
rect 28089 20213 28123 20247
rect 29101 20213 29135 20247
rect 29751 20213 29785 20247
rect 31125 20213 31159 20247
rect 31585 20213 31619 20247
rect 33333 20213 33367 20247
rect 36461 20213 36495 20247
rect 37289 20213 37323 20247
rect 13921 20009 13955 20043
rect 16681 20009 16715 20043
rect 16957 20009 16991 20043
rect 17417 20009 17451 20043
rect 18889 20009 18923 20043
rect 19625 20009 19659 20043
rect 21189 20009 21223 20043
rect 21925 20009 21959 20043
rect 23673 20009 23707 20043
rect 24041 20009 24075 20043
rect 25145 20009 25179 20043
rect 26157 20009 26191 20043
rect 29009 20009 29043 20043
rect 29745 20009 29779 20043
rect 31217 20009 31251 20043
rect 32321 20009 32355 20043
rect 33431 20009 33465 20043
rect 34805 20009 34839 20043
rect 35173 20009 35207 20043
rect 15568 19941 15602 19975
rect 17754 19941 17788 19975
rect 19901 19941 19935 19975
rect 23397 19941 23431 19975
rect 27537 19941 27571 19975
rect 30104 19941 30138 19975
rect 17509 19873 17543 19907
rect 22293 19873 22327 19907
rect 24409 19873 24443 19907
rect 26525 19873 26559 19907
rect 27896 19873 27930 19907
rect 29837 19873 29871 19907
rect 36001 19873 36035 19907
rect 15301 19805 15335 19839
rect 21833 19805 21867 19839
rect 22385 19805 22419 19839
rect 22569 19805 22603 19839
rect 24501 19805 24535 19839
rect 24593 19805 24627 19839
rect 27169 19805 27203 19839
rect 27629 19805 27663 19839
rect 32965 19805 32999 19839
rect 33471 19805 33505 19839
rect 33701 19805 33735 19839
rect 36093 19805 36127 19839
rect 36277 19805 36311 19839
rect 35449 19737 35483 19771
rect 35633 19737 35667 19771
rect 19257 19669 19291 19703
rect 20545 19669 20579 19703
rect 26709 19669 26743 19703
rect 29377 19669 29411 19703
rect 32873 19669 32907 19703
rect 15945 19465 15979 19499
rect 17601 19465 17635 19499
rect 18245 19465 18279 19499
rect 18613 19465 18647 19499
rect 22017 19465 22051 19499
rect 26525 19465 26559 19499
rect 27905 19465 27939 19499
rect 33057 19465 33091 19499
rect 14565 19329 14599 19363
rect 19533 19329 19567 19363
rect 19993 19329 20027 19363
rect 24777 19329 24811 19363
rect 28181 19329 28215 19363
rect 29837 19329 29871 19363
rect 30252 19329 30286 19363
rect 30435 19329 30469 19363
rect 30665 19329 30699 19363
rect 34713 19329 34747 19363
rect 35449 19329 35483 19363
rect 14832 19261 14866 19295
rect 22201 19261 22235 19295
rect 22753 19261 22787 19295
rect 25789 19261 25823 19295
rect 26893 19261 26927 19295
rect 27445 19261 27479 19295
rect 29929 19261 29963 19295
rect 32689 19261 32723 19295
rect 35716 19261 35750 19295
rect 37105 19261 37139 19295
rect 14473 19193 14507 19227
rect 19901 19193 19935 19227
rect 20260 19193 20294 19227
rect 23489 19193 23523 19227
rect 25329 19193 25363 19227
rect 29101 19193 29135 19227
rect 33793 19193 33827 19227
rect 16221 19125 16255 19159
rect 16589 19125 16623 19159
rect 21373 19125 21407 19159
rect 22385 19125 22419 19159
rect 24041 19125 24075 19159
rect 24225 19125 24259 19159
rect 24593 19125 24627 19159
rect 24685 19125 24719 19159
rect 25697 19125 25731 19159
rect 25973 19125 26007 19159
rect 27077 19125 27111 19159
rect 28641 19125 28675 19159
rect 31769 19125 31803 19159
rect 33425 19125 33459 19159
rect 35357 19125 35391 19159
rect 36829 19125 36863 19159
rect 14565 18921 14599 18955
rect 15577 18921 15611 18955
rect 22569 18921 22603 18955
rect 24225 18921 24259 18955
rect 24593 18921 24627 18955
rect 24777 18921 24811 18955
rect 25973 18921 26007 18955
rect 26709 18921 26743 18955
rect 27629 18921 27663 18955
rect 28733 18921 28767 18955
rect 29193 18921 29227 18955
rect 29929 18921 29963 18955
rect 30757 18921 30791 18955
rect 30849 18921 30883 18955
rect 31493 18921 31527 18955
rect 33149 18921 33183 18955
rect 34529 18921 34563 18955
rect 36001 18921 36035 18955
rect 19717 18853 19751 18887
rect 29101 18853 29135 18887
rect 36093 18853 36127 18887
rect 19625 18785 19659 18819
rect 21180 18785 21214 18819
rect 23489 18785 23523 18819
rect 25145 18785 25179 18819
rect 26525 18785 26559 18819
rect 27813 18785 27847 18819
rect 34437 18785 34471 18819
rect 19901 18717 19935 18751
rect 20913 18717 20947 18751
rect 23581 18717 23615 18751
rect 23673 18717 23707 18751
rect 25237 18717 25271 18751
rect 25329 18717 25363 18751
rect 28089 18717 28123 18751
rect 29285 18717 29319 18751
rect 31033 18717 31067 18751
rect 34621 18717 34655 18751
rect 35449 18717 35483 18751
rect 36185 18717 36219 18751
rect 23121 18649 23155 18683
rect 30389 18649 30423 18683
rect 34069 18649 34103 18683
rect 19257 18581 19291 18615
rect 22293 18581 22327 18615
rect 32781 18581 32815 18615
rect 35633 18581 35667 18615
rect 19349 18377 19383 18411
rect 19625 18377 19659 18411
rect 21189 18377 21223 18411
rect 22017 18377 22051 18411
rect 23213 18377 23247 18411
rect 24869 18377 24903 18411
rect 28365 18377 28399 18411
rect 28825 18377 28859 18411
rect 29469 18377 29503 18411
rect 30481 18377 30515 18411
rect 31125 18377 31159 18411
rect 33793 18377 33827 18411
rect 34069 18377 34103 18411
rect 34437 18377 34471 18411
rect 35725 18377 35759 18411
rect 36001 18377 36035 18411
rect 36369 18377 36403 18411
rect 25789 18309 25823 18343
rect 27997 18309 28031 18343
rect 29929 18309 29963 18343
rect 21925 18241 21959 18275
rect 22477 18241 22511 18275
rect 22569 18241 22603 18275
rect 27721 18241 27755 18275
rect 30757 18241 30791 18275
rect 32229 18241 32263 18275
rect 33241 18241 33275 18275
rect 19809 18173 19843 18207
rect 22385 18173 22419 18207
rect 23857 18173 23891 18207
rect 25973 18173 26007 18207
rect 33057 18173 33091 18207
rect 18981 18105 19015 18139
rect 20076 18105 20110 18139
rect 24409 18105 24443 18139
rect 32597 18105 32631 18139
rect 33149 18105 33183 18139
rect 18613 18037 18647 18071
rect 21557 18037 21591 18071
rect 25237 18037 25271 18071
rect 32689 18037 32723 18071
rect 22293 17833 22327 17867
rect 22569 17833 22603 17867
rect 23305 17833 23339 17867
rect 23673 17833 23707 17867
rect 27905 17833 27939 17867
rect 34805 17833 34839 17867
rect 19625 17765 19659 17799
rect 21180 17765 21214 17799
rect 24501 17765 24535 17799
rect 24860 17765 24894 17799
rect 26770 17765 26804 17799
rect 22937 17697 22971 17731
rect 23121 17697 23155 17731
rect 24593 17697 24627 17731
rect 26525 17697 26559 17731
rect 32505 17697 32539 17731
rect 32597 17697 32631 17731
rect 34713 17697 34747 17731
rect 35909 17697 35943 17731
rect 19717 17629 19751 17663
rect 19901 17629 19935 17663
rect 20913 17629 20947 17663
rect 30297 17629 30331 17663
rect 32689 17629 32723 17663
rect 34897 17629 34931 17663
rect 29377 17561 29411 17595
rect 19257 17493 19291 17527
rect 20269 17493 20303 17527
rect 20637 17493 20671 17527
rect 25973 17493 26007 17527
rect 29745 17493 29779 17527
rect 31677 17493 31711 17527
rect 32137 17493 32171 17527
rect 34345 17493 34379 17527
rect 35541 17493 35575 17527
rect 36093 17493 36127 17527
rect 18981 17289 19015 17323
rect 21097 17289 21131 17323
rect 25237 17289 25271 17323
rect 26709 17289 26743 17323
rect 26985 17289 27019 17323
rect 28733 17289 28767 17323
rect 34345 17289 34379 17323
rect 36553 17289 36587 17323
rect 21925 17221 21959 17255
rect 29285 17221 29319 17255
rect 22569 17153 22603 17187
rect 29837 17153 29871 17187
rect 35909 17153 35943 17187
rect 36001 17153 36035 17187
rect 19717 17085 19751 17119
rect 19984 17085 20018 17119
rect 22293 17085 22327 17119
rect 22937 17085 22971 17119
rect 23857 17085 23891 17119
rect 25329 17085 25363 17119
rect 27905 17085 27939 17119
rect 28181 17085 28215 17119
rect 28365 17085 28399 17119
rect 31585 17085 31619 17119
rect 36829 17085 36863 17119
rect 21741 17017 21775 17051
rect 22385 17017 22419 17051
rect 23489 17017 23523 17051
rect 24124 17017 24158 17051
rect 25574 17017 25608 17051
rect 27997 17017 28031 17051
rect 29653 17017 29687 17051
rect 31401 17017 31435 17051
rect 31852 17017 31886 17051
rect 33241 17017 33275 17051
rect 33793 17017 33827 17051
rect 35357 17017 35391 17051
rect 18613 16949 18647 16983
rect 19349 16949 19383 16983
rect 21373 16949 21407 16983
rect 27353 16949 27387 16983
rect 29009 16949 29043 16983
rect 29745 16949 29779 16983
rect 31125 16949 31159 16983
rect 32965 16949 32999 16983
rect 33609 16949 33643 16983
rect 35449 16949 35483 16983
rect 35817 16949 35851 16983
rect 19257 16745 19291 16779
rect 20361 16745 20395 16779
rect 22293 16745 22327 16779
rect 22569 16745 22603 16779
rect 23121 16745 23155 16779
rect 23949 16745 23983 16779
rect 24317 16745 24351 16779
rect 24409 16745 24443 16779
rect 24869 16745 24903 16779
rect 25513 16745 25547 16779
rect 25881 16745 25915 16779
rect 27077 16745 27111 16779
rect 27445 16745 27479 16779
rect 29745 16745 29779 16779
rect 31953 16745 31987 16779
rect 32413 16745 32447 16779
rect 33247 16745 33281 16779
rect 34621 16745 34655 16779
rect 34897 16745 34931 16779
rect 36829 16745 36863 16779
rect 19165 16677 19199 16711
rect 24777 16677 24811 16711
rect 28610 16677 28644 16711
rect 35694 16677 35728 16711
rect 19625 16609 19659 16643
rect 21180 16609 21214 16643
rect 27261 16609 27295 16643
rect 28365 16609 28399 16643
rect 30573 16609 30607 16643
rect 31125 16609 31159 16643
rect 32781 16609 32815 16643
rect 33517 16609 33551 16643
rect 19717 16541 19751 16575
rect 19901 16541 19935 16575
rect 20913 16541 20947 16575
rect 24961 16541 24995 16575
rect 33244 16541 33278 16575
rect 35449 16541 35483 16575
rect 20729 16405 20763 16439
rect 30757 16405 30791 16439
rect 35357 16405 35391 16439
rect 19349 16201 19383 16235
rect 19625 16201 19659 16235
rect 21373 16201 21407 16235
rect 24133 16201 24167 16235
rect 24225 16201 24259 16235
rect 24501 16201 24535 16235
rect 25237 16201 25271 16235
rect 28365 16201 28399 16235
rect 28641 16201 28675 16235
rect 31953 16201 31987 16235
rect 33885 16201 33919 16235
rect 34529 16201 34563 16235
rect 35357 16201 35391 16235
rect 19993 15997 20027 16031
rect 20260 15997 20294 16031
rect 32045 16065 32079 16099
rect 32508 16065 32542 16099
rect 34161 16065 34195 16099
rect 25513 15997 25547 16031
rect 26065 15997 26099 16031
rect 26985 15997 27019 16031
rect 29101 15997 29135 16031
rect 29561 15997 29595 16031
rect 32781 15997 32815 16031
rect 35449 15997 35483 16031
rect 35705 15997 35739 16031
rect 24225 15929 24259 15963
rect 27230 15929 27264 15963
rect 29806 15929 29840 15963
rect 37105 15929 37139 15963
rect 18981 15861 19015 15895
rect 21741 15861 21775 15895
rect 22109 15861 22143 15895
rect 24961 15861 24995 15895
rect 25697 15861 25731 15895
rect 26801 15861 26835 15895
rect 30941 15861 30975 15895
rect 31585 15861 31619 15895
rect 32511 15861 32545 15895
rect 36829 15861 36863 15895
rect 20085 15657 20119 15691
rect 22293 15657 22327 15691
rect 23949 15657 23983 15691
rect 24869 15657 24903 15691
rect 26893 15657 26927 15691
rect 27629 15657 27663 15691
rect 28733 15657 28767 15691
rect 29653 15657 29687 15691
rect 30665 15657 30699 15691
rect 31585 15657 31619 15691
rect 35817 15657 35851 15691
rect 36645 15657 36679 15691
rect 21158 15589 21192 15623
rect 25973 15589 26007 15623
rect 26985 15589 27019 15623
rect 28641 15589 28675 15623
rect 30757 15589 30791 15623
rect 32474 15589 32508 15623
rect 36093 15589 36127 15623
rect 23857 15521 23891 15555
rect 24133 15521 24167 15555
rect 24777 15521 24811 15555
rect 25237 15521 25271 15555
rect 32229 15521 32263 15555
rect 34693 15521 34727 15555
rect 20453 15453 20487 15487
rect 20913 15453 20947 15487
rect 25329 15453 25363 15487
rect 25513 15453 25547 15487
rect 27169 15453 27203 15487
rect 28917 15453 28951 15487
rect 30941 15453 30975 15487
rect 34437 15453 34471 15487
rect 26525 15385 26559 15419
rect 30021 15385 30055 15419
rect 28273 15317 28307 15351
rect 30297 15317 30331 15351
rect 31953 15317 31987 15351
rect 33609 15317 33643 15351
rect 20913 15113 20947 15147
rect 23857 15113 23891 15147
rect 24961 15113 24995 15147
rect 27537 15113 27571 15147
rect 28457 15113 28491 15147
rect 28733 15113 28767 15147
rect 29469 15113 29503 15147
rect 29837 15113 29871 15147
rect 30389 15113 30423 15147
rect 30757 15113 30791 15147
rect 31033 15113 31067 15147
rect 32597 15113 32631 15147
rect 32873 15113 32907 15147
rect 33241 15113 33275 15147
rect 34253 15113 34287 15147
rect 34529 15113 34563 15147
rect 34621 15113 34655 15147
rect 21281 15045 21315 15079
rect 24409 14977 24443 15011
rect 33425 14977 33459 15011
rect 35449 14977 35483 15011
rect 25421 14909 25455 14943
rect 27813 14909 27847 14943
rect 29285 14909 29319 14943
rect 31217 14909 31251 14943
rect 31473 14909 31507 14943
rect 34529 14909 34563 14943
rect 35265 14909 35299 14943
rect 24317 14841 24351 14875
rect 25329 14841 25363 14875
rect 25666 14841 25700 14875
rect 35357 14841 35391 14875
rect 23029 14773 23063 14807
rect 23489 14773 23523 14807
rect 24225 14773 24259 14807
rect 26801 14773 26835 14807
rect 27077 14773 27111 14807
rect 27997 14773 28031 14807
rect 33885 14773 33919 14807
rect 34897 14773 34931 14807
rect 23305 14569 23339 14603
rect 23949 14569 23983 14603
rect 25605 14569 25639 14603
rect 26709 14569 26743 14603
rect 27077 14569 27111 14603
rect 28365 14569 28399 14603
rect 29285 14569 29319 14603
rect 29929 14569 29963 14603
rect 30665 14569 30699 14603
rect 32229 14569 32263 14603
rect 34897 14569 34931 14603
rect 35265 14569 35299 14603
rect 24470 14501 24504 14535
rect 25881 14501 25915 14535
rect 32689 14501 32723 14535
rect 23121 14433 23155 14467
rect 24225 14433 24259 14467
rect 27445 14433 27479 14467
rect 28641 14433 28675 14467
rect 29745 14433 29779 14467
rect 32597 14433 32631 14467
rect 27537 14365 27571 14399
rect 27721 14365 27755 14399
rect 32873 14365 32907 14399
rect 21373 14229 21407 14263
rect 28825 14229 28859 14263
rect 30389 14229 30423 14263
rect 31309 14229 31343 14263
rect 34437 14229 34471 14263
rect 23489 14025 23523 14059
rect 25053 14025 25087 14059
rect 25421 14025 25455 14059
rect 25697 14025 25731 14059
rect 25881 14025 25915 14059
rect 27169 14025 27203 14059
rect 27629 14025 27663 14059
rect 28365 14025 28399 14059
rect 29101 14025 29135 14059
rect 29745 14025 29779 14059
rect 31309 14025 31343 14059
rect 31493 14025 31527 14059
rect 32689 14025 32723 14059
rect 32965 14025 32999 14059
rect 28549 13957 28583 13991
rect 21373 13889 21407 13923
rect 26341 13889 26375 13923
rect 26433 13889 26467 13923
rect 30389 13889 30423 13923
rect 30573 13889 30607 13923
rect 23121 13821 23155 13855
rect 23673 13821 23707 13855
rect 23929 13821 23963 13855
rect 27445 13821 27479 13855
rect 27997 13821 28031 13855
rect 28733 13821 28767 13855
rect 30297 13821 30331 13855
rect 31033 13821 31067 13855
rect 31677 13821 31711 13855
rect 21281 13753 21315 13787
rect 21618 13753 21652 13787
rect 22753 13685 22787 13719
rect 26249 13685 26283 13719
rect 29929 13685 29963 13719
rect 32321 13685 32355 13719
rect 34897 13685 34931 13719
rect 21649 13481 21683 13515
rect 24133 13481 24167 13515
rect 24409 13481 24443 13515
rect 25053 13481 25087 13515
rect 25513 13481 25547 13515
rect 27169 13481 27203 13515
rect 28641 13481 28675 13515
rect 29009 13481 29043 13515
rect 30481 13481 30515 13515
rect 30941 13481 30975 13515
rect 32597 13481 32631 13515
rect 35817 13481 35851 13515
rect 25973 13413 26007 13447
rect 21557 13345 21591 13379
rect 23020 13345 23054 13379
rect 25237 13345 25271 13379
rect 25329 13345 25363 13379
rect 27721 13345 27755 13379
rect 29285 13345 29319 13379
rect 29837 13345 29871 13379
rect 33865 13345 33899 13379
rect 36185 13345 36219 13379
rect 21741 13277 21775 13311
rect 22753 13277 22787 13311
rect 24869 13277 24903 13311
rect 27813 13277 27847 13311
rect 27905 13277 27939 13311
rect 29929 13277 29963 13311
rect 30021 13277 30055 13311
rect 33609 13277 33643 13311
rect 36277 13277 36311 13311
rect 36461 13277 36495 13311
rect 29101 13209 29135 13243
rect 31493 13209 31527 13243
rect 21189 13141 21223 13175
rect 22569 13141 22603 13175
rect 27353 13141 27387 13175
rect 29469 13141 29503 13175
rect 34989 13141 35023 13175
rect 35357 13141 35391 13175
rect 20545 12937 20579 12971
rect 22753 12937 22787 12971
rect 23029 12937 23063 12971
rect 23673 12937 23707 12971
rect 24777 12937 24811 12971
rect 25145 12937 25179 12971
rect 26801 12937 26835 12971
rect 27813 12937 27847 12971
rect 28181 12937 28215 12971
rect 29101 12937 29135 12971
rect 32137 12937 32171 12971
rect 34713 12937 34747 12971
rect 36921 12937 36955 12971
rect 37565 12937 37599 12971
rect 20913 12869 20947 12903
rect 21281 12869 21315 12903
rect 26341 12869 26375 12903
rect 28733 12869 28767 12903
rect 31769 12869 31803 12903
rect 32413 12869 32447 12903
rect 32597 12869 32631 12903
rect 36553 12869 36587 12903
rect 21373 12801 21407 12835
rect 24317 12801 24351 12835
rect 26709 12801 26743 12835
rect 27261 12801 27295 12835
rect 27445 12801 27479 12835
rect 30392 12801 30426 12835
rect 33149 12801 33183 12835
rect 33609 12801 33643 12835
rect 37105 12801 37139 12835
rect 25421 12733 25455 12767
rect 29929 12733 29963 12767
rect 30665 12733 30699 12767
rect 33057 12733 33091 12767
rect 34069 12733 34103 12767
rect 34897 12733 34931 12767
rect 35153 12733 35187 12767
rect 21618 12665 21652 12699
rect 23489 12665 23523 12699
rect 24133 12665 24167 12699
rect 25697 12665 25731 12699
rect 32965 12665 32999 12699
rect 24041 12597 24075 12631
rect 25237 12597 25271 12631
rect 27169 12597 27203 12631
rect 29837 12597 29871 12631
rect 30395 12597 30429 12631
rect 36277 12597 36311 12631
rect 21465 12393 21499 12427
rect 23397 12393 23431 12427
rect 23673 12393 23707 12427
rect 24041 12393 24075 12427
rect 24225 12393 24259 12427
rect 25237 12393 25271 12427
rect 28733 12393 28767 12427
rect 29193 12393 29227 12427
rect 29561 12393 29595 12427
rect 31125 12393 31159 12427
rect 36829 12393 36863 12427
rect 27261 12325 27295 12359
rect 35357 12325 35391 12359
rect 35716 12325 35750 12359
rect 22273 12257 22307 12291
rect 24593 12257 24627 12291
rect 27620 12257 27654 12291
rect 30012 12257 30046 12291
rect 33104 12257 33138 12291
rect 34897 12257 34931 12291
rect 35449 12257 35483 12291
rect 22017 12189 22051 12223
rect 24685 12189 24719 12223
rect 24777 12189 24811 12223
rect 27353 12189 27387 12223
rect 29745 12189 29779 12223
rect 32781 12189 32815 12223
rect 33244 12189 33278 12223
rect 33517 12189 33551 12223
rect 21833 12053 21867 12087
rect 26893 12053 26927 12087
rect 31953 12053 31987 12087
rect 32505 12053 32539 12087
rect 34621 12053 34655 12087
rect 22109 11849 22143 11883
rect 23397 11849 23431 11883
rect 23673 11849 23707 11883
rect 25053 11849 25087 11883
rect 26617 11849 26651 11883
rect 30665 11849 30699 11883
rect 32413 11849 32447 11883
rect 33885 11849 33919 11883
rect 34161 11849 34195 11883
rect 36001 11849 36035 11883
rect 36277 11849 36311 11883
rect 31401 11781 31435 11815
rect 34621 11781 34655 11815
rect 23121 11713 23155 11747
rect 24225 11713 24259 11747
rect 28733 11713 28767 11747
rect 32505 11713 32539 11747
rect 35357 11713 35391 11747
rect 35541 11713 35575 11747
rect 24041 11645 24075 11679
rect 25881 11645 25915 11679
rect 26249 11645 26283 11679
rect 26709 11645 26743 11679
rect 29285 11645 29319 11679
rect 29552 11645 29586 11679
rect 32045 11645 32079 11679
rect 35265 11645 35299 11679
rect 36461 11645 36495 11679
rect 37013 11645 37047 11679
rect 24133 11577 24167 11611
rect 26954 11577 26988 11611
rect 30941 11577 30975 11611
rect 32750 11577 32784 11611
rect 22385 11509 22419 11543
rect 24685 11509 24719 11543
rect 28089 11509 28123 11543
rect 29101 11509 29135 11543
rect 31493 11509 31527 11543
rect 34897 11509 34931 11543
rect 36645 11509 36679 11543
rect 23581 11305 23615 11339
rect 24317 11305 24351 11339
rect 24409 11305 24443 11339
rect 30665 11305 30699 11339
rect 31953 11305 31987 11339
rect 33517 11305 33551 11339
rect 34897 11305 34931 11339
rect 36461 11305 36495 11339
rect 27344 11237 27378 11271
rect 29552 11237 29586 11271
rect 34345 11237 34379 11271
rect 34989 11237 35023 11271
rect 36093 11237 36127 11271
rect 22457 11169 22491 11203
rect 24777 11169 24811 11203
rect 27077 11169 27111 11203
rect 32404 11169 32438 11203
rect 36277 11169 36311 11203
rect 22201 11101 22235 11135
rect 24869 11101 24903 11135
rect 25053 11101 25087 11135
rect 29285 11101 29319 11135
rect 32137 11101 32171 11135
rect 35081 11101 35115 11135
rect 28457 11033 28491 11067
rect 34529 11033 34563 11067
rect 26801 10965 26835 10999
rect 35633 10965 35667 10999
rect 22293 10761 22327 10795
rect 25421 10761 25455 10795
rect 27629 10761 27663 10795
rect 29929 10761 29963 10795
rect 31769 10761 31803 10795
rect 31953 10761 31987 10795
rect 34529 10761 34563 10795
rect 29469 10625 29503 10659
rect 31493 10625 31527 10659
rect 32505 10625 32539 10659
rect 33057 10625 33091 10659
rect 22661 10557 22695 10591
rect 23121 10557 23155 10591
rect 23673 10557 23707 10591
rect 25881 10557 25915 10591
rect 30665 10557 30699 10591
rect 30849 10557 30883 10591
rect 32321 10557 32355 10591
rect 33517 10557 33551 10591
rect 34069 10557 34103 10591
rect 35449 10557 35483 10591
rect 23489 10489 23523 10523
rect 23918 10489 23952 10523
rect 25789 10489 25823 10523
rect 26148 10489 26182 10523
rect 30389 10489 30423 10523
rect 33425 10489 33459 10523
rect 35357 10489 35391 10523
rect 35716 10489 35750 10523
rect 25053 10421 25087 10455
rect 27261 10421 27295 10455
rect 27997 10421 28031 10455
rect 29009 10421 29043 10455
rect 30481 10421 30515 10455
rect 31033 10421 31067 10455
rect 32413 10421 32447 10455
rect 33701 10421 33735 10455
rect 36829 10421 36863 10455
rect 37105 10421 37139 10455
rect 24133 10217 24167 10251
rect 24777 10217 24811 10251
rect 26985 10217 27019 10251
rect 27353 10217 27387 10251
rect 30573 10217 30607 10251
rect 31493 10217 31527 10251
rect 31953 10217 31987 10251
rect 32413 10217 32447 10251
rect 32873 10217 32907 10251
rect 34161 10217 34195 10251
rect 34621 10217 34655 10251
rect 36093 10217 36127 10251
rect 32781 10149 32815 10183
rect 22753 10081 22787 10115
rect 23009 10081 23043 10115
rect 24409 10081 24443 10115
rect 33517 10081 33551 10115
rect 33977 10081 34011 10115
rect 35449 10081 35483 10115
rect 36553 10081 36587 10115
rect 27445 10013 27479 10047
rect 27537 10013 27571 10047
rect 33057 10013 33091 10047
rect 35265 9945 35299 9979
rect 25881 9877 25915 9911
rect 31125 9877 31159 9911
rect 35633 9877 35667 9911
rect 36737 9877 36771 9911
rect 22845 9673 22879 9707
rect 26157 9673 26191 9707
rect 26525 9673 26559 9707
rect 32505 9673 32539 9707
rect 33977 9673 34011 9707
rect 36553 9673 36587 9707
rect 22477 9605 22511 9639
rect 28365 9605 28399 9639
rect 29653 9605 29687 9639
rect 30849 9605 30883 9639
rect 32137 9605 32171 9639
rect 32873 9605 32907 9639
rect 35173 9605 35207 9639
rect 36277 9605 36311 9639
rect 37289 9605 37323 9639
rect 26893 9537 26927 9571
rect 27905 9537 27939 9571
rect 31493 9537 31527 9571
rect 31585 9537 31619 9571
rect 33425 9537 33459 9571
rect 35725 9537 35759 9571
rect 23765 9469 23799 9503
rect 29469 9469 29503 9503
rect 30021 9469 30055 9503
rect 31401 9469 31435 9503
rect 33241 9469 33275 9503
rect 36737 9469 36771 9503
rect 23489 9401 23523 9435
rect 24032 9401 24066 9435
rect 27261 9401 27295 9435
rect 27813 9401 27847 9435
rect 30573 9401 30607 9435
rect 35633 9401 35667 9435
rect 25145 9333 25179 9367
rect 27353 9333 27387 9367
rect 27721 9333 27755 9367
rect 31033 9333 31067 9367
rect 33333 9333 33367 9367
rect 34621 9333 34655 9367
rect 35541 9333 35575 9367
rect 36921 9333 36955 9367
rect 24133 9129 24167 9163
rect 27445 9129 27479 9163
rect 31033 9129 31067 9163
rect 33241 9129 33275 9163
rect 34345 9129 34379 9163
rect 36829 9129 36863 9163
rect 24501 9061 24535 9095
rect 24593 9061 24627 9095
rect 31953 9061 31987 9095
rect 32965 9061 32999 9095
rect 34897 9061 34931 9095
rect 23857 8993 23891 9027
rect 28089 8993 28123 9027
rect 29193 8993 29227 9027
rect 29653 8993 29687 9027
rect 30849 8993 30883 9027
rect 32137 8993 32171 9027
rect 33609 8993 33643 9027
rect 35449 8993 35483 9027
rect 35716 8993 35750 9027
rect 24685 8925 24719 8959
rect 28181 8925 28215 8959
rect 28273 8925 28307 8959
rect 29745 8925 29779 8959
rect 29929 8925 29963 8959
rect 33701 8925 33735 8959
rect 33885 8925 33919 8959
rect 27077 8857 27111 8891
rect 29285 8857 29319 8891
rect 27721 8789 27755 8823
rect 28825 8789 28859 8823
rect 30297 8789 30331 8823
rect 32321 8789 32355 8823
rect 35265 8789 35299 8823
rect 24501 8585 24535 8619
rect 26709 8585 26743 8619
rect 27169 8585 27203 8619
rect 27537 8585 27571 8619
rect 29653 8585 29687 8619
rect 30665 8585 30699 8619
rect 33241 8585 33275 8619
rect 34713 8585 34747 8619
rect 36829 8585 36863 8619
rect 25145 8517 25179 8551
rect 27629 8517 27663 8551
rect 28641 8517 28675 8551
rect 24225 8449 24259 8483
rect 28089 8449 28123 8483
rect 28273 8449 28307 8483
rect 30205 8449 30239 8483
rect 32045 8449 32079 8483
rect 32597 8449 32631 8483
rect 32689 8449 32723 8483
rect 25329 8381 25363 8415
rect 25585 8381 25619 8415
rect 27997 8381 28031 8415
rect 29101 8381 29135 8415
rect 30021 8381 30055 8415
rect 31677 8381 31711 8415
rect 32505 8381 32539 8415
rect 33701 8381 33735 8415
rect 34253 8381 34287 8415
rect 35449 8381 35483 8415
rect 29561 8313 29595 8347
rect 30113 8313 30147 8347
rect 31309 8313 31343 8347
rect 35357 8313 35391 8347
rect 35716 8313 35750 8347
rect 32137 8245 32171 8279
rect 33885 8245 33919 8279
rect 37105 8245 37139 8279
rect 24225 8041 24259 8075
rect 28181 8041 28215 8075
rect 28549 8041 28583 8075
rect 30849 8041 30883 8075
rect 31861 8041 31895 8075
rect 32597 8041 32631 8075
rect 33333 8041 33367 8075
rect 33701 8041 33735 8075
rect 34069 8041 34103 8075
rect 36645 8041 36679 8075
rect 26770 7973 26804 8007
rect 29000 7905 29034 7939
rect 32505 7905 32539 7939
rect 34989 7905 35023 7939
rect 35265 7905 35299 7939
rect 35532 7905 35566 7939
rect 25421 7837 25455 7871
rect 26525 7837 26559 7871
rect 28733 7837 28767 7871
rect 32781 7837 32815 7871
rect 34161 7837 34195 7871
rect 34345 7837 34379 7871
rect 32137 7769 32171 7803
rect 27905 7701 27939 7735
rect 30113 7701 30147 7735
rect 26249 7497 26283 7531
rect 26617 7497 26651 7531
rect 28273 7497 28307 7531
rect 28733 7497 28767 7531
rect 30665 7497 30699 7531
rect 33149 7497 33183 7531
rect 34161 7497 34195 7531
rect 37013 7497 37047 7531
rect 31309 7429 31343 7463
rect 32873 7429 32907 7463
rect 29009 7361 29043 7395
rect 26893 7293 26927 7327
rect 27160 7293 27194 7327
rect 29285 7293 29319 7327
rect 29541 7293 29575 7327
rect 31493 7293 31527 7327
rect 34897 7293 34931 7327
rect 31738 7225 31772 7259
rect 35142 7225 35176 7259
rect 33793 7157 33827 7191
rect 34621 7157 34655 7191
rect 36277 7157 36311 7191
rect 36553 7157 36587 7191
rect 26985 6953 27019 6987
rect 31953 6953 31987 6987
rect 32321 6953 32355 6987
rect 34253 6953 34287 6987
rect 36093 6953 36127 6987
rect 29736 6885 29770 6919
rect 27528 6817 27562 6851
rect 29009 6817 29043 6851
rect 29377 6817 29411 6851
rect 29469 6817 29503 6851
rect 32772 6817 32806 6851
rect 34713 6817 34747 6851
rect 34969 6817 35003 6851
rect 27261 6749 27295 6783
rect 31585 6749 31619 6783
rect 32505 6749 32539 6783
rect 28641 6681 28675 6715
rect 30849 6613 30883 6647
rect 33885 6613 33919 6647
rect 27353 6409 27387 6443
rect 29101 6409 29135 6443
rect 30941 6409 30975 6443
rect 33149 6409 33183 6443
rect 36277 6409 36311 6443
rect 36645 6409 36679 6443
rect 31677 6273 31711 6307
rect 34345 6273 34379 6307
rect 26985 6205 27019 6239
rect 27721 6205 27755 6239
rect 28733 6205 28767 6239
rect 29561 6205 29595 6239
rect 29828 6205 29862 6239
rect 31769 6205 31803 6239
rect 32036 6205 32070 6239
rect 34897 6205 34931 6239
rect 35164 6205 35198 6239
rect 34621 6069 34655 6103
rect 28825 5865 28859 5899
rect 29193 5865 29227 5899
rect 29837 5865 29871 5899
rect 32597 5865 32631 5899
rect 33241 5865 33275 5899
rect 34897 5865 34931 5899
rect 35265 5865 35299 5899
rect 29285 5797 29319 5831
rect 30297 5797 30331 5831
rect 31861 5797 31895 5831
rect 32965 5797 32999 5831
rect 34805 5797 34839 5831
rect 35357 5797 35391 5831
rect 33609 5729 33643 5763
rect 29377 5661 29411 5695
rect 33701 5661 33735 5695
rect 33793 5661 33827 5695
rect 35449 5661 35483 5695
rect 28549 5321 28583 5355
rect 28917 5321 28951 5355
rect 29469 5321 29503 5355
rect 33333 5321 33367 5355
rect 33977 5321 34011 5355
rect 34621 5321 34655 5355
rect 35541 5321 35575 5355
rect 33609 5253 33643 5287
rect 35173 5253 35207 5287
rect 33885 2601 33919 2635
rect 33333 2465 33367 2499
rect 33517 2329 33551 2363
rect 8401 2261 8435 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 7009 36907 7067 36913
rect 7009 36873 7021 36907
rect 7055 36904 7067 36907
rect 7190 36904 7196 36916
rect 7055 36876 7196 36904
rect 7055 36873 7067 36876
rect 7009 36867 7067 36873
rect 7190 36864 7196 36876
rect 7248 36864 7254 36916
rect 6825 36703 6883 36709
rect 6825 36669 6837 36703
rect 6871 36700 6883 36703
rect 6871 36672 7512 36700
rect 6871 36669 6883 36672
rect 6825 36663 6883 36669
rect 7484 36576 7512 36672
rect 7466 36564 7472 36576
rect 7427 36536 7472 36564
rect 7466 36524 7472 36536
rect 7524 36524 7530 36576
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 22649 36295 22707 36301
rect 22649 36261 22661 36295
rect 22695 36292 22707 36295
rect 22830 36292 22836 36304
rect 22695 36264 22836 36292
rect 22695 36261 22707 36264
rect 22649 36255 22707 36261
rect 22830 36252 22836 36264
rect 22888 36252 22894 36304
rect 6822 36224 6828 36236
rect 6783 36196 6828 36224
rect 6822 36184 6828 36196
rect 6880 36184 6886 36236
rect 15654 36224 15660 36236
rect 15615 36196 15660 36224
rect 15654 36184 15660 36196
rect 15712 36184 15718 36236
rect 23845 36227 23903 36233
rect 23845 36193 23857 36227
rect 23891 36224 23903 36227
rect 24762 36224 24768 36236
rect 23891 36196 24768 36224
rect 23891 36193 23903 36196
rect 23845 36187 23903 36193
rect 24762 36184 24768 36196
rect 24820 36184 24826 36236
rect 15746 36156 15752 36168
rect 15707 36128 15752 36156
rect 15746 36116 15752 36128
rect 15804 36116 15810 36168
rect 15930 36156 15936 36168
rect 15891 36128 15936 36156
rect 15930 36116 15936 36128
rect 15988 36116 15994 36168
rect 22462 36116 22468 36168
rect 22520 36156 22526 36168
rect 22741 36159 22799 36165
rect 22741 36156 22753 36159
rect 22520 36128 22753 36156
rect 22520 36116 22526 36128
rect 22741 36125 22753 36128
rect 22787 36125 22799 36159
rect 22922 36156 22928 36168
rect 22883 36128 22928 36156
rect 22741 36119 22799 36125
rect 22922 36116 22928 36128
rect 22980 36116 22986 36168
rect 7009 36023 7067 36029
rect 7009 35989 7021 36023
rect 7055 36020 7067 36023
rect 7374 36020 7380 36032
rect 7055 35992 7380 36020
rect 7055 35989 7067 35992
rect 7009 35983 7067 35989
rect 7374 35980 7380 35992
rect 7432 35980 7438 36032
rect 13998 36020 14004 36032
rect 13959 35992 14004 36020
rect 13998 35980 14004 35992
rect 14056 35980 14062 36032
rect 15194 35980 15200 36032
rect 15252 36020 15258 36032
rect 15289 36023 15347 36029
rect 15289 36020 15301 36023
rect 15252 35992 15301 36020
rect 15252 35980 15258 35992
rect 15289 35989 15301 35992
rect 15335 35989 15347 36023
rect 15289 35983 15347 35989
rect 21453 36023 21511 36029
rect 21453 35989 21465 36023
rect 21499 36020 21511 36023
rect 21726 36020 21732 36032
rect 21499 35992 21732 36020
rect 21499 35989 21511 35992
rect 21453 35983 21511 35989
rect 21726 35980 21732 35992
rect 21784 35980 21790 36032
rect 22278 36020 22284 36032
rect 22239 35992 22284 36020
rect 22278 35980 22284 35992
rect 22336 35980 22342 36032
rect 24029 36023 24087 36029
rect 24029 35989 24041 36023
rect 24075 36020 24087 36023
rect 24210 36020 24216 36032
rect 24075 35992 24216 36020
rect 24075 35989 24087 35992
rect 24029 35983 24087 35989
rect 24210 35980 24216 35992
rect 24268 35980 24274 36032
rect 24946 36020 24952 36032
rect 24907 35992 24952 36020
rect 24946 35980 24952 35992
rect 25004 35980 25010 36032
rect 26234 35980 26240 36032
rect 26292 36020 26298 36032
rect 26697 36023 26755 36029
rect 26697 36020 26709 36023
rect 26292 35992 26709 36020
rect 26292 35980 26298 35992
rect 26697 35989 26709 35992
rect 26743 35989 26755 36023
rect 26697 35983 26755 35989
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 5629 35819 5687 35825
rect 5629 35785 5641 35819
rect 5675 35816 5687 35819
rect 6086 35816 6092 35828
rect 5675 35788 6092 35816
rect 5675 35785 5687 35788
rect 5629 35779 5687 35785
rect 6086 35776 6092 35788
rect 6144 35776 6150 35828
rect 6822 35776 6828 35828
rect 6880 35816 6886 35828
rect 7742 35816 7748 35828
rect 6880 35788 7748 35816
rect 6880 35776 6886 35788
rect 7742 35776 7748 35788
rect 7800 35776 7806 35828
rect 8294 35776 8300 35828
rect 8352 35816 8358 35828
rect 8389 35819 8447 35825
rect 8389 35816 8401 35819
rect 8352 35788 8401 35816
rect 8352 35776 8358 35788
rect 8389 35785 8401 35788
rect 8435 35785 8447 35819
rect 8389 35779 8447 35785
rect 15746 35776 15752 35828
rect 15804 35816 15810 35828
rect 15933 35819 15991 35825
rect 15933 35816 15945 35819
rect 15804 35788 15945 35816
rect 15804 35776 15810 35788
rect 15933 35785 15945 35788
rect 15979 35785 15991 35819
rect 22462 35816 22468 35828
rect 22423 35788 22468 35816
rect 15933 35779 15991 35785
rect 22462 35776 22468 35788
rect 22520 35776 22526 35828
rect 22830 35816 22836 35828
rect 22791 35788 22836 35816
rect 22830 35776 22836 35788
rect 22888 35776 22894 35828
rect 24673 35819 24731 35825
rect 24673 35785 24685 35819
rect 24719 35816 24731 35819
rect 24762 35816 24768 35828
rect 24719 35788 24768 35816
rect 24719 35785 24731 35788
rect 24673 35779 24731 35785
rect 24762 35776 24768 35788
rect 24820 35776 24826 35828
rect 35618 35816 35624 35828
rect 35579 35788 35624 35816
rect 35618 35776 35624 35788
rect 35676 35776 35682 35828
rect 15654 35748 15660 35760
rect 15615 35720 15660 35748
rect 15654 35708 15660 35720
rect 15712 35708 15718 35760
rect 20162 35708 20168 35760
rect 20220 35748 20226 35760
rect 21361 35751 21419 35757
rect 21361 35748 21373 35751
rect 20220 35720 21373 35748
rect 20220 35708 20226 35720
rect 21361 35717 21373 35720
rect 21407 35717 21419 35751
rect 22922 35748 22928 35760
rect 21361 35711 21419 35717
rect 22020 35720 22928 35748
rect 22020 35692 22048 35720
rect 22922 35708 22928 35720
rect 22980 35748 22986 35760
rect 23109 35751 23167 35757
rect 23109 35748 23121 35751
rect 22980 35720 23121 35748
rect 22980 35708 22986 35720
rect 23109 35717 23121 35720
rect 23155 35717 23167 35751
rect 23109 35711 23167 35717
rect 22002 35680 22008 35692
rect 21963 35652 22008 35680
rect 22002 35640 22008 35652
rect 22060 35640 22066 35692
rect 26234 35640 26240 35692
rect 26292 35680 26298 35692
rect 26881 35683 26939 35689
rect 26881 35680 26893 35683
rect 26292 35652 26893 35680
rect 26292 35640 26298 35652
rect 26881 35649 26893 35652
rect 26927 35649 26939 35683
rect 26881 35643 26939 35649
rect 5445 35615 5503 35621
rect 5445 35581 5457 35615
rect 5491 35612 5503 35615
rect 7098 35612 7104 35624
rect 5491 35584 6132 35612
rect 7059 35584 7104 35612
rect 5491 35581 5503 35584
rect 5445 35575 5503 35581
rect 6104 35488 6132 35584
rect 7098 35572 7104 35584
rect 7156 35572 7162 35624
rect 8205 35615 8263 35621
rect 8205 35581 8217 35615
rect 8251 35612 8263 35615
rect 13909 35615 13967 35621
rect 8251 35584 8892 35612
rect 8251 35581 8263 35584
rect 8205 35575 8263 35581
rect 8864 35556 8892 35584
rect 13909 35581 13921 35615
rect 13955 35612 13967 35615
rect 13998 35612 14004 35624
rect 13955 35584 14004 35612
rect 13955 35581 13967 35584
rect 13909 35575 13967 35581
rect 13998 35572 14004 35584
rect 14056 35572 14062 35624
rect 15378 35572 15384 35624
rect 15436 35612 15442 35624
rect 15930 35612 15936 35624
rect 15436 35584 15936 35612
rect 15436 35572 15442 35584
rect 15930 35572 15936 35584
rect 15988 35612 15994 35624
rect 16301 35615 16359 35621
rect 16301 35612 16313 35615
rect 15988 35584 16313 35612
rect 15988 35572 15994 35584
rect 16301 35581 16313 35584
rect 16347 35581 16359 35615
rect 21726 35612 21732 35624
rect 21687 35584 21732 35612
rect 16301 35575 16359 35581
rect 21726 35572 21732 35584
rect 21784 35572 21790 35624
rect 23661 35615 23719 35621
rect 23661 35581 23673 35615
rect 23707 35612 23719 35615
rect 23842 35612 23848 35624
rect 23707 35584 23848 35612
rect 23707 35581 23719 35584
rect 23661 35575 23719 35581
rect 23842 35572 23848 35584
rect 23900 35612 23906 35624
rect 24213 35615 24271 35621
rect 24213 35612 24225 35615
rect 23900 35584 24225 35612
rect 23900 35572 23906 35584
rect 24213 35581 24225 35584
rect 24259 35581 24271 35615
rect 24946 35612 24952 35624
rect 24907 35584 24952 35612
rect 24213 35575 24271 35581
rect 24946 35572 24952 35584
rect 25004 35572 25010 35624
rect 25869 35615 25927 35621
rect 25869 35581 25881 35615
rect 25915 35612 25927 35615
rect 26694 35612 26700 35624
rect 25915 35584 26700 35612
rect 25915 35581 25927 35584
rect 25869 35575 25927 35581
rect 26694 35572 26700 35584
rect 26752 35572 26758 35624
rect 34514 35572 34520 35624
rect 34572 35612 34578 35624
rect 35437 35615 35495 35621
rect 35437 35612 35449 35615
rect 34572 35584 35449 35612
rect 34572 35572 34578 35584
rect 35437 35581 35449 35584
rect 35483 35612 35495 35615
rect 35989 35615 36047 35621
rect 35989 35612 36001 35615
rect 35483 35584 36001 35612
rect 35483 35581 35495 35584
rect 35437 35575 35495 35581
rect 35989 35581 36001 35584
rect 36035 35581 36047 35615
rect 35989 35575 36047 35581
rect 8846 35544 8852 35556
rect 8807 35516 8852 35544
rect 8846 35504 8852 35516
rect 8904 35504 8910 35556
rect 13817 35547 13875 35553
rect 13817 35513 13829 35547
rect 13863 35544 13875 35547
rect 14154 35547 14212 35553
rect 14154 35544 14166 35547
rect 13863 35516 14166 35544
rect 13863 35513 13875 35516
rect 13817 35507 13875 35513
rect 14154 35513 14166 35516
rect 14200 35544 14212 35547
rect 15838 35544 15844 35556
rect 14200 35516 15844 35544
rect 14200 35513 14212 35516
rect 14154 35507 14212 35513
rect 15838 35504 15844 35516
rect 15896 35504 15902 35556
rect 21821 35547 21879 35553
rect 21821 35544 21833 35547
rect 21192 35516 21833 35544
rect 6086 35476 6092 35488
rect 6047 35448 6092 35476
rect 6086 35436 6092 35448
rect 6144 35436 6150 35488
rect 7282 35476 7288 35488
rect 7243 35448 7288 35476
rect 7282 35436 7288 35448
rect 7340 35436 7346 35488
rect 12250 35436 12256 35488
rect 12308 35476 12314 35488
rect 12437 35479 12495 35485
rect 12437 35476 12449 35479
rect 12308 35448 12449 35476
rect 12308 35436 12314 35448
rect 12437 35445 12449 35448
rect 12483 35445 12495 35479
rect 12437 35439 12495 35445
rect 15289 35479 15347 35485
rect 15289 35445 15301 35479
rect 15335 35476 15347 35479
rect 15378 35476 15384 35488
rect 15335 35448 15384 35476
rect 15335 35445 15347 35448
rect 15289 35439 15347 35445
rect 15378 35436 15384 35448
rect 15436 35436 15442 35488
rect 20898 35476 20904 35488
rect 20859 35448 20904 35476
rect 20898 35436 20904 35448
rect 20956 35436 20962 35488
rect 21082 35436 21088 35488
rect 21140 35476 21146 35488
rect 21192 35485 21220 35516
rect 21821 35513 21833 35516
rect 21867 35513 21879 35547
rect 21821 35507 21879 35513
rect 26237 35547 26295 35553
rect 26237 35513 26249 35547
rect 26283 35544 26295 35547
rect 26510 35544 26516 35556
rect 26283 35516 26516 35544
rect 26283 35513 26295 35516
rect 26237 35507 26295 35513
rect 26510 35504 26516 35516
rect 26568 35544 26574 35556
rect 26789 35547 26847 35553
rect 26789 35544 26801 35547
rect 26568 35516 26801 35544
rect 26568 35504 26574 35516
rect 26789 35513 26801 35516
rect 26835 35513 26847 35547
rect 26789 35507 26847 35513
rect 21177 35479 21235 35485
rect 21177 35476 21189 35479
rect 21140 35448 21189 35476
rect 21140 35436 21146 35448
rect 21177 35445 21189 35448
rect 21223 35445 21235 35479
rect 21177 35439 21235 35445
rect 23566 35436 23572 35488
rect 23624 35476 23630 35488
rect 23845 35479 23903 35485
rect 23845 35476 23857 35479
rect 23624 35448 23857 35476
rect 23624 35436 23630 35448
rect 23845 35445 23857 35448
rect 23891 35445 23903 35479
rect 25130 35476 25136 35488
rect 25091 35448 25136 35476
rect 23845 35439 23903 35445
rect 25130 35436 25136 35448
rect 25188 35436 25194 35488
rect 26326 35476 26332 35488
rect 26287 35448 26332 35476
rect 26326 35436 26332 35448
rect 26384 35436 26390 35488
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 1581 35275 1639 35281
rect 1581 35241 1593 35275
rect 1627 35272 1639 35275
rect 1670 35272 1676 35284
rect 1627 35244 1676 35272
rect 1627 35241 1639 35244
rect 1581 35235 1639 35241
rect 1670 35232 1676 35244
rect 1728 35232 1734 35284
rect 4341 35275 4399 35281
rect 4341 35241 4353 35275
rect 4387 35272 4399 35275
rect 4982 35272 4988 35284
rect 4387 35244 4988 35272
rect 4387 35241 4399 35244
rect 4341 35235 4399 35241
rect 4982 35232 4988 35244
rect 5040 35232 5046 35284
rect 7098 35272 7104 35284
rect 7059 35244 7104 35272
rect 7098 35232 7104 35244
rect 7156 35232 7162 35284
rect 12526 35232 12532 35284
rect 12584 35272 12590 35284
rect 13265 35275 13323 35281
rect 13265 35272 13277 35275
rect 12584 35244 13277 35272
rect 12584 35232 12590 35244
rect 13265 35241 13277 35244
rect 13311 35272 13323 35275
rect 13998 35272 14004 35284
rect 13311 35244 14004 35272
rect 13311 35241 13323 35244
rect 13265 35235 13323 35241
rect 13998 35232 14004 35244
rect 14056 35272 14062 35284
rect 14734 35272 14740 35284
rect 14056 35244 14740 35272
rect 14056 35232 14062 35244
rect 14734 35232 14740 35244
rect 14792 35232 14798 35284
rect 15286 35272 15292 35284
rect 15247 35244 15292 35272
rect 15286 35232 15292 35244
rect 15344 35232 15350 35284
rect 19705 35275 19763 35281
rect 19705 35241 19717 35275
rect 19751 35272 19763 35275
rect 20254 35272 20260 35284
rect 19751 35244 20260 35272
rect 19751 35241 19763 35244
rect 19705 35235 19763 35241
rect 20254 35232 20260 35244
rect 20312 35232 20318 35284
rect 20898 35232 20904 35284
rect 20956 35272 20962 35284
rect 21177 35275 21235 35281
rect 21177 35272 21189 35275
rect 20956 35244 21189 35272
rect 20956 35232 20962 35244
rect 21177 35241 21189 35244
rect 21223 35272 21235 35275
rect 22002 35272 22008 35284
rect 21223 35244 22008 35272
rect 21223 35241 21235 35244
rect 21177 35235 21235 35241
rect 22002 35232 22008 35244
rect 22060 35232 22066 35284
rect 22830 35232 22836 35284
rect 22888 35272 22894 35284
rect 23474 35272 23480 35284
rect 22888 35244 23480 35272
rect 22888 35232 22894 35244
rect 23474 35232 23480 35244
rect 23532 35232 23538 35284
rect 24857 35275 24915 35281
rect 24857 35241 24869 35275
rect 24903 35272 24915 35275
rect 24946 35272 24952 35284
rect 24903 35244 24952 35272
rect 24903 35241 24915 35244
rect 24857 35235 24915 35241
rect 24946 35232 24952 35244
rect 25004 35232 25010 35284
rect 25038 35232 25044 35284
rect 25096 35272 25102 35284
rect 25225 35275 25283 35281
rect 25225 35272 25237 35275
rect 25096 35244 25237 35272
rect 25096 35232 25102 35244
rect 25225 35241 25237 35244
rect 25271 35272 25283 35275
rect 26326 35272 26332 35284
rect 25271 35244 26332 35272
rect 25271 35241 25283 35244
rect 25225 35235 25283 35241
rect 26326 35232 26332 35244
rect 26384 35232 26390 35284
rect 35526 35272 35532 35284
rect 35487 35244 35532 35272
rect 35526 35232 35532 35244
rect 35584 35232 35590 35284
rect 9490 35164 9496 35216
rect 9548 35204 9554 35216
rect 9677 35207 9735 35213
rect 9677 35204 9689 35207
rect 9548 35176 9689 35204
rect 9548 35164 9554 35176
rect 9677 35173 9689 35176
rect 9723 35204 9735 35207
rect 10686 35204 10692 35216
rect 9723 35176 10692 35204
rect 9723 35173 9735 35176
rect 9677 35167 9735 35173
rect 10686 35164 10692 35176
rect 10744 35164 10750 35216
rect 22364 35207 22422 35213
rect 22364 35173 22376 35207
rect 22410 35204 22422 35207
rect 22462 35204 22468 35216
rect 22410 35176 22468 35204
rect 22410 35173 22422 35176
rect 22364 35167 22422 35173
rect 22462 35164 22468 35176
rect 22520 35164 22526 35216
rect 1394 35136 1400 35148
rect 1355 35108 1400 35136
rect 1394 35096 1400 35108
rect 1452 35096 1458 35148
rect 4157 35139 4215 35145
rect 4157 35105 4169 35139
rect 4203 35136 4215 35139
rect 4706 35136 4712 35148
rect 4203 35108 4712 35136
rect 4203 35105 4215 35108
rect 4157 35099 4215 35105
rect 4706 35096 4712 35108
rect 4764 35096 4770 35148
rect 5166 35096 5172 35148
rect 5224 35136 5230 35148
rect 5517 35139 5575 35145
rect 5517 35136 5529 35139
rect 5224 35108 5529 35136
rect 5224 35096 5230 35108
rect 5517 35105 5529 35108
rect 5563 35105 5575 35139
rect 5517 35099 5575 35105
rect 8297 35139 8355 35145
rect 8297 35105 8309 35139
rect 8343 35136 8355 35139
rect 9122 35136 9128 35148
rect 8343 35108 9128 35136
rect 8343 35105 8355 35108
rect 8297 35099 8355 35105
rect 9122 35096 9128 35108
rect 9180 35096 9186 35148
rect 9858 35136 9864 35148
rect 9819 35108 9864 35136
rect 9858 35096 9864 35108
rect 9916 35096 9922 35148
rect 11790 35145 11796 35148
rect 11784 35136 11796 35145
rect 11751 35108 11796 35136
rect 11784 35099 11796 35108
rect 11790 35096 11796 35099
rect 11848 35096 11854 35148
rect 13725 35139 13783 35145
rect 13725 35105 13737 35139
rect 13771 35136 13783 35139
rect 14182 35136 14188 35148
rect 13771 35108 14188 35136
rect 13771 35105 13783 35108
rect 13725 35099 13783 35105
rect 14182 35096 14188 35108
rect 14240 35096 14246 35148
rect 14642 35096 14648 35148
rect 14700 35136 14706 35148
rect 15657 35139 15715 35145
rect 15657 35136 15669 35139
rect 14700 35108 15669 35136
rect 14700 35096 14706 35108
rect 15657 35105 15669 35108
rect 15703 35105 15715 35139
rect 17218 35136 17224 35148
rect 17179 35108 17224 35136
rect 15657 35099 15715 35105
rect 17218 35096 17224 35108
rect 17276 35096 17282 35148
rect 18417 35139 18475 35145
rect 18417 35105 18429 35139
rect 18463 35136 18475 35139
rect 19150 35136 19156 35148
rect 18463 35108 19156 35136
rect 18463 35105 18475 35108
rect 18417 35099 18475 35105
rect 19150 35096 19156 35108
rect 19208 35096 19214 35148
rect 20990 35136 20996 35148
rect 20951 35108 20996 35136
rect 20990 35096 20996 35108
rect 21048 35096 21054 35148
rect 26142 35096 26148 35148
rect 26200 35136 26206 35148
rect 26769 35139 26827 35145
rect 26769 35136 26781 35139
rect 26200 35108 26781 35136
rect 26200 35096 26206 35108
rect 26769 35105 26781 35108
rect 26815 35105 26827 35139
rect 26769 35099 26827 35105
rect 35345 35139 35403 35145
rect 35345 35105 35357 35139
rect 35391 35136 35403 35139
rect 35710 35136 35716 35148
rect 35391 35108 35716 35136
rect 35391 35105 35403 35108
rect 35345 35099 35403 35105
rect 35710 35096 35716 35108
rect 35768 35096 35774 35148
rect 5261 35071 5319 35077
rect 5261 35037 5273 35071
rect 5307 35037 5319 35071
rect 11514 35068 11520 35080
rect 11475 35040 11520 35068
rect 5261 35031 5319 35037
rect 5276 34932 5304 35031
rect 11514 35028 11520 35040
rect 11572 35028 11578 35080
rect 15746 35068 15752 35080
rect 15707 35040 15752 35068
rect 15746 35028 15752 35040
rect 15804 35028 15810 35080
rect 15838 35028 15844 35080
rect 15896 35068 15902 35080
rect 17310 35068 17316 35080
rect 15896 35040 15941 35068
rect 17271 35040 17316 35068
rect 15896 35028 15902 35040
rect 17310 35028 17316 35040
rect 17368 35028 17374 35080
rect 17405 35071 17463 35077
rect 17405 35037 17417 35071
rect 17451 35037 17463 35071
rect 22097 35071 22155 35077
rect 22097 35068 22109 35071
rect 17405 35031 17463 35037
rect 21560 35040 22109 35068
rect 16850 35000 16856 35012
rect 16811 34972 16856 35000
rect 16850 34960 16856 34972
rect 16908 34960 16914 35012
rect 17034 34960 17040 35012
rect 17092 35000 17098 35012
rect 17420 35000 17448 35031
rect 17092 34972 17448 35000
rect 18141 35003 18199 35009
rect 17092 34960 17098 34972
rect 18141 34969 18153 35003
rect 18187 35000 18199 35003
rect 18690 35000 18696 35012
rect 18187 34972 18696 35000
rect 18187 34969 18199 34972
rect 18141 34963 18199 34969
rect 18690 34960 18696 34972
rect 18748 34960 18754 35012
rect 5902 34932 5908 34944
rect 5276 34904 5908 34932
rect 5902 34892 5908 34904
rect 5960 34892 5966 34944
rect 6638 34932 6644 34944
rect 6599 34904 6644 34932
rect 6638 34892 6644 34904
rect 6696 34892 6702 34944
rect 7466 34932 7472 34944
rect 7427 34904 7472 34932
rect 7466 34892 7472 34904
rect 7524 34892 7530 34944
rect 8294 34892 8300 34944
rect 8352 34932 8358 34944
rect 8481 34935 8539 34941
rect 8481 34932 8493 34935
rect 8352 34904 8493 34932
rect 8352 34892 8358 34904
rect 8481 34901 8493 34904
rect 8527 34901 8539 34935
rect 8481 34895 8539 34901
rect 9674 34892 9680 34944
rect 9732 34932 9738 34944
rect 10045 34935 10103 34941
rect 10045 34932 10057 34935
rect 9732 34904 10057 34932
rect 9732 34892 9738 34904
rect 10045 34901 10057 34904
rect 10091 34901 10103 34935
rect 10318 34932 10324 34944
rect 10279 34904 10324 34932
rect 10045 34895 10103 34901
rect 10318 34892 10324 34904
rect 10376 34892 10382 34944
rect 12802 34892 12808 34944
rect 12860 34932 12866 34944
rect 12897 34935 12955 34941
rect 12897 34932 12909 34935
rect 12860 34904 12909 34932
rect 12860 34892 12866 34904
rect 12897 34901 12909 34904
rect 12943 34901 12955 34935
rect 12897 34895 12955 34901
rect 13814 34892 13820 34944
rect 13872 34932 13878 34944
rect 13909 34935 13967 34941
rect 13909 34932 13921 34935
rect 13872 34904 13921 34932
rect 13872 34892 13878 34904
rect 13909 34901 13921 34904
rect 13955 34901 13967 34935
rect 13909 34895 13967 34901
rect 18046 34892 18052 34944
rect 18104 34932 18110 34944
rect 18601 34935 18659 34941
rect 18601 34932 18613 34935
rect 18104 34904 18613 34932
rect 18104 34892 18110 34904
rect 18601 34901 18613 34904
rect 18647 34901 18659 34935
rect 18601 34895 18659 34901
rect 20898 34892 20904 34944
rect 20956 34932 20962 34944
rect 21560 34941 21588 35040
rect 22097 35037 22109 35040
rect 22143 35037 22155 35071
rect 22097 35031 22155 35037
rect 24765 35071 24823 35077
rect 24765 35037 24777 35071
rect 24811 35068 24823 35071
rect 25314 35068 25320 35080
rect 24811 35040 25320 35068
rect 24811 35037 24823 35040
rect 24765 35031 24823 35037
rect 25314 35028 25320 35040
rect 25372 35028 25378 35080
rect 25409 35071 25467 35077
rect 25409 35037 25421 35071
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 23566 34960 23572 35012
rect 23624 35000 23630 35012
rect 24305 35003 24363 35009
rect 24305 35000 24317 35003
rect 23624 34972 24317 35000
rect 23624 34960 23630 34972
rect 24305 34969 24317 34972
rect 24351 35000 24363 35003
rect 25424 35000 25452 35031
rect 26418 35028 26424 35080
rect 26476 35068 26482 35080
rect 26513 35071 26571 35077
rect 26513 35068 26525 35071
rect 26476 35040 26525 35068
rect 26476 35028 26482 35040
rect 26513 35037 26525 35040
rect 26559 35037 26571 35071
rect 26513 35031 26571 35037
rect 24351 34972 25452 35000
rect 24351 34969 24363 34972
rect 24305 34963 24363 34969
rect 21545 34935 21603 34941
rect 21545 34932 21557 34935
rect 20956 34904 21557 34932
rect 20956 34892 20962 34904
rect 21545 34901 21557 34904
rect 21591 34901 21603 34935
rect 24026 34932 24032 34944
rect 23987 34904 24032 34932
rect 21545 34895 21603 34901
rect 24026 34892 24032 34904
rect 24084 34892 24090 34944
rect 26510 34892 26516 34944
rect 26568 34932 26574 34944
rect 27893 34935 27951 34941
rect 27893 34932 27905 34935
rect 26568 34904 27905 34932
rect 26568 34892 26574 34904
rect 27893 34901 27905 34904
rect 27939 34901 27951 34935
rect 27893 34895 27951 34901
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 566 34688 572 34740
rect 624 34728 630 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 624 34700 1593 34728
rect 624 34688 630 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 2038 34728 2044 34740
rect 1999 34700 2044 34728
rect 1581 34691 1639 34697
rect 2038 34688 2044 34700
rect 2096 34688 2102 34740
rect 3789 34731 3847 34737
rect 3789 34697 3801 34731
rect 3835 34728 3847 34731
rect 3878 34728 3884 34740
rect 3835 34700 3884 34728
rect 3835 34697 3847 34700
rect 3789 34691 3847 34697
rect 3878 34688 3884 34700
rect 3936 34688 3942 34740
rect 4249 34731 4307 34737
rect 4249 34697 4261 34731
rect 4295 34728 4307 34731
rect 4614 34728 4620 34740
rect 4295 34700 4620 34728
rect 4295 34697 4307 34700
rect 4249 34691 4307 34697
rect 2682 34660 2688 34672
rect 2643 34632 2688 34660
rect 2682 34620 2688 34632
rect 2740 34620 2746 34672
rect 3142 34592 3148 34604
rect 2516 34564 3148 34592
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 2038 34524 2044 34536
rect 1443 34496 2044 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2516 34533 2544 34564
rect 3142 34552 3148 34564
rect 3200 34552 3206 34604
rect 2501 34527 2559 34533
rect 2501 34493 2513 34527
rect 2547 34493 2559 34527
rect 2501 34487 2559 34493
rect 3605 34527 3663 34533
rect 3605 34493 3617 34527
rect 3651 34524 3663 34527
rect 4264 34524 4292 34691
rect 4614 34688 4620 34700
rect 4672 34688 4678 34740
rect 9122 34728 9128 34740
rect 9083 34700 9128 34728
rect 9122 34688 9128 34700
rect 9180 34688 9186 34740
rect 9490 34728 9496 34740
rect 9451 34700 9496 34728
rect 9490 34688 9496 34700
rect 9548 34688 9554 34740
rect 9858 34688 9864 34740
rect 9916 34728 9922 34740
rect 10597 34731 10655 34737
rect 10597 34728 10609 34731
rect 9916 34700 10609 34728
rect 9916 34688 9922 34700
rect 10597 34697 10609 34700
rect 10643 34697 10655 34731
rect 10597 34691 10655 34697
rect 11701 34731 11759 34737
rect 11701 34697 11713 34731
rect 11747 34728 11759 34731
rect 11790 34728 11796 34740
rect 11747 34700 11796 34728
rect 11747 34697 11759 34700
rect 11701 34691 11759 34697
rect 11790 34688 11796 34700
rect 11848 34728 11854 34740
rect 12434 34728 12440 34740
rect 11848 34700 12440 34728
rect 11848 34688 11854 34700
rect 12434 34688 12440 34700
rect 12492 34688 12498 34740
rect 14182 34728 14188 34740
rect 14143 34700 14188 34728
rect 14182 34688 14188 34700
rect 14240 34688 14246 34740
rect 14642 34728 14648 34740
rect 14603 34700 14648 34728
rect 14642 34688 14648 34700
rect 14700 34688 14706 34740
rect 15838 34688 15844 34740
rect 15896 34728 15902 34740
rect 16117 34731 16175 34737
rect 16117 34728 16129 34731
rect 15896 34700 16129 34728
rect 15896 34688 15902 34700
rect 16117 34697 16129 34700
rect 16163 34728 16175 34731
rect 16393 34731 16451 34737
rect 16393 34728 16405 34731
rect 16163 34700 16405 34728
rect 16163 34697 16175 34700
rect 16117 34691 16175 34697
rect 16393 34697 16405 34700
rect 16439 34697 16451 34731
rect 17218 34728 17224 34740
rect 16393 34691 16451 34697
rect 16960 34700 17224 34728
rect 5169 34663 5227 34669
rect 5169 34629 5181 34663
rect 5215 34660 5227 34663
rect 5442 34660 5448 34672
rect 5215 34632 5448 34660
rect 5215 34629 5227 34632
rect 5169 34623 5227 34629
rect 5442 34620 5448 34632
rect 5500 34620 5506 34672
rect 8757 34663 8815 34669
rect 8757 34629 8769 34663
rect 8803 34660 8815 34663
rect 8846 34660 8852 34672
rect 8803 34632 8852 34660
rect 8803 34629 8815 34632
rect 8757 34623 8815 34629
rect 8846 34620 8852 34632
rect 8904 34660 8910 34672
rect 9876 34660 9904 34688
rect 8904 34632 9904 34660
rect 13909 34663 13967 34669
rect 8904 34620 8910 34632
rect 13909 34629 13921 34663
rect 13955 34660 13967 34663
rect 14274 34660 14280 34672
rect 13955 34632 14280 34660
rect 13955 34629 13967 34632
rect 13909 34623 13967 34629
rect 14274 34620 14280 34632
rect 14332 34620 14338 34672
rect 15746 34620 15752 34672
rect 15804 34660 15810 34672
rect 16761 34663 16819 34669
rect 16761 34660 16773 34663
rect 15804 34632 16773 34660
rect 15804 34620 15810 34632
rect 16761 34629 16773 34632
rect 16807 34629 16819 34663
rect 16761 34623 16819 34629
rect 4617 34595 4675 34601
rect 4617 34561 4629 34595
rect 4663 34592 4675 34595
rect 4706 34592 4712 34604
rect 4663 34564 4712 34592
rect 4663 34561 4675 34564
rect 4617 34555 4675 34561
rect 4706 34552 4712 34564
rect 4764 34552 4770 34604
rect 5813 34595 5871 34601
rect 5813 34561 5825 34595
rect 5859 34592 5871 34595
rect 6086 34592 6092 34604
rect 5859 34564 6092 34592
rect 5859 34561 5871 34564
rect 5813 34555 5871 34561
rect 6086 34552 6092 34564
rect 6144 34592 6150 34604
rect 7282 34592 7288 34604
rect 6144 34564 7288 34592
rect 6144 34552 6150 34564
rect 7282 34552 7288 34564
rect 7340 34552 7346 34604
rect 10134 34592 10140 34604
rect 10095 34564 10140 34592
rect 10134 34552 10140 34564
rect 10192 34552 10198 34604
rect 12253 34595 12311 34601
rect 12253 34561 12265 34595
rect 12299 34592 12311 34595
rect 12342 34592 12348 34604
rect 12299 34564 12348 34592
rect 12299 34561 12311 34564
rect 12253 34555 12311 34561
rect 12342 34552 12348 34564
rect 12400 34592 12406 34604
rect 14734 34592 14740 34604
rect 12400 34564 12664 34592
rect 14695 34564 14740 34592
rect 12400 34552 12406 34564
rect 3651 34496 4292 34524
rect 3651 34493 3663 34496
rect 3605 34487 3663 34493
rect 5902 34484 5908 34536
rect 5960 34524 5966 34536
rect 6549 34527 6607 34533
rect 6549 34524 6561 34527
rect 5960 34496 6561 34524
rect 5960 34484 5966 34496
rect 6549 34493 6561 34496
rect 6595 34524 6607 34527
rect 7377 34527 7435 34533
rect 7377 34524 7389 34527
rect 6595 34496 7389 34524
rect 6595 34493 6607 34496
rect 6549 34487 6607 34493
rect 7377 34493 7389 34496
rect 7423 34524 7435 34527
rect 7466 34524 7472 34536
rect 7423 34496 7472 34524
rect 7423 34493 7435 34496
rect 7377 34487 7435 34493
rect 7466 34484 7472 34496
rect 7524 34524 7530 34536
rect 8386 34524 8392 34536
rect 7524 34496 8392 34524
rect 7524 34484 7530 34496
rect 8386 34484 8392 34496
rect 8444 34484 8450 34536
rect 9766 34484 9772 34536
rect 9824 34524 9830 34536
rect 10045 34527 10103 34533
rect 10045 34524 10057 34527
rect 9824 34496 10057 34524
rect 9824 34484 9830 34496
rect 10045 34493 10057 34496
rect 10091 34524 10103 34527
rect 10965 34527 11023 34533
rect 10965 34524 10977 34527
rect 10091 34496 10977 34524
rect 10091 34493 10103 34496
rect 10045 34487 10103 34493
rect 10965 34493 10977 34496
rect 11011 34493 11023 34527
rect 12526 34524 12532 34536
rect 12487 34496 12532 34524
rect 10965 34487 11023 34493
rect 12526 34484 12532 34496
rect 12584 34484 12590 34536
rect 12636 34524 12664 34564
rect 14734 34552 14740 34564
rect 14792 34552 14798 34604
rect 16960 34601 16988 34700
rect 17218 34688 17224 34700
rect 17276 34728 17282 34740
rect 17405 34731 17463 34737
rect 17405 34728 17417 34731
rect 17276 34700 17417 34728
rect 17276 34688 17282 34700
rect 17405 34697 17417 34700
rect 17451 34697 17463 34731
rect 19150 34728 19156 34740
rect 19111 34700 19156 34728
rect 17405 34691 17463 34697
rect 19150 34688 19156 34700
rect 19208 34688 19214 34740
rect 20990 34728 20996 34740
rect 20951 34700 20996 34728
rect 20990 34688 20996 34700
rect 21048 34688 21054 34740
rect 22462 34688 22468 34740
rect 22520 34728 22526 34740
rect 22557 34731 22615 34737
rect 22557 34728 22569 34731
rect 22520 34700 22569 34728
rect 22520 34688 22526 34700
rect 22557 34697 22569 34700
rect 22603 34728 22615 34731
rect 22833 34731 22891 34737
rect 22833 34728 22845 34731
rect 22603 34700 22845 34728
rect 22603 34697 22615 34700
rect 22557 34691 22615 34697
rect 22833 34697 22845 34700
rect 22879 34697 22891 34731
rect 22833 34691 22891 34697
rect 23937 34731 23995 34737
rect 23937 34697 23949 34731
rect 23983 34728 23995 34731
rect 25038 34728 25044 34740
rect 23983 34700 25044 34728
rect 23983 34697 23995 34700
rect 23937 34691 23995 34697
rect 25038 34688 25044 34700
rect 25096 34688 25102 34740
rect 25777 34731 25835 34737
rect 25777 34697 25789 34731
rect 25823 34728 25835 34731
rect 26142 34728 26148 34740
rect 25823 34700 26148 34728
rect 25823 34697 25835 34700
rect 25777 34691 25835 34697
rect 26142 34688 26148 34700
rect 26200 34688 26206 34740
rect 26510 34728 26516 34740
rect 26471 34700 26516 34728
rect 26510 34688 26516 34700
rect 26568 34688 26574 34740
rect 26786 34688 26792 34740
rect 26844 34728 26850 34740
rect 27985 34731 28043 34737
rect 27985 34728 27997 34731
rect 26844 34700 27997 34728
rect 26844 34688 26850 34700
rect 27985 34697 27997 34700
rect 28031 34697 28043 34731
rect 27985 34691 28043 34697
rect 35621 34731 35679 34737
rect 35621 34697 35633 34731
rect 35667 34728 35679 34731
rect 35802 34728 35808 34740
rect 35667 34700 35808 34728
rect 35667 34697 35679 34700
rect 35621 34691 35679 34697
rect 35802 34688 35808 34700
rect 35860 34688 35866 34740
rect 36722 34728 36728 34740
rect 36683 34700 36728 34728
rect 36722 34688 36728 34700
rect 36780 34688 36786 34740
rect 18049 34663 18107 34669
rect 18049 34629 18061 34663
rect 18095 34660 18107 34663
rect 18138 34660 18144 34672
rect 18095 34632 18144 34660
rect 18095 34629 18107 34632
rect 18049 34623 18107 34629
rect 18138 34620 18144 34632
rect 18196 34620 18202 34672
rect 19613 34663 19671 34669
rect 19613 34629 19625 34663
rect 19659 34660 19671 34663
rect 20530 34660 20536 34672
rect 19659 34632 20536 34660
rect 19659 34629 19671 34632
rect 19613 34623 19671 34629
rect 20530 34620 20536 34632
rect 20588 34620 20594 34672
rect 16945 34595 17003 34601
rect 16945 34561 16957 34595
rect 16991 34561 17003 34595
rect 16945 34555 17003 34561
rect 17954 34552 17960 34604
rect 18012 34592 18018 34604
rect 18509 34595 18567 34601
rect 18509 34592 18521 34595
rect 18012 34564 18521 34592
rect 18012 34552 18018 34564
rect 18509 34561 18521 34564
rect 18555 34561 18567 34595
rect 18690 34592 18696 34604
rect 18603 34564 18696 34592
rect 18509 34555 18567 34561
rect 12802 34533 12808 34536
rect 12796 34524 12808 34533
rect 12636 34496 12808 34524
rect 12796 34487 12808 34496
rect 12802 34484 12808 34487
rect 12860 34484 12866 34536
rect 17678 34484 17684 34536
rect 17736 34524 17742 34536
rect 17773 34527 17831 34533
rect 17773 34524 17785 34527
rect 17736 34496 17785 34524
rect 17736 34484 17742 34496
rect 17773 34493 17785 34496
rect 17819 34524 17831 34527
rect 18524 34524 18552 34555
rect 18690 34552 18696 34564
rect 18748 34592 18754 34604
rect 19150 34592 19156 34604
rect 18748 34564 19156 34592
rect 18748 34552 18754 34564
rect 19150 34552 19156 34564
rect 19208 34552 19214 34604
rect 20070 34552 20076 34604
rect 20128 34592 20134 34604
rect 20165 34595 20223 34601
rect 20165 34592 20177 34595
rect 20128 34564 20177 34592
rect 20128 34552 20134 34564
rect 20165 34561 20177 34564
rect 20211 34561 20223 34595
rect 20165 34555 20223 34561
rect 20717 34595 20775 34601
rect 20717 34561 20729 34595
rect 20763 34592 20775 34595
rect 24305 34595 24363 34601
rect 20763 34564 21312 34592
rect 20763 34561 20775 34564
rect 20717 34555 20775 34561
rect 19429 34527 19487 34533
rect 19429 34524 19441 34527
rect 17819 34496 17908 34524
rect 18524 34496 19441 34524
rect 17819 34493 17831 34496
rect 17773 34487 17831 34493
rect 5537 34459 5595 34465
rect 5537 34425 5549 34459
rect 5583 34456 5595 34459
rect 7622 34459 7680 34465
rect 7622 34456 7634 34459
rect 5583 34428 6316 34456
rect 5583 34425 5595 34428
rect 5537 34419 5595 34425
rect 6288 34400 6316 34428
rect 7208 34428 7634 34456
rect 7208 34400 7236 34428
rect 7622 34425 7634 34428
rect 7668 34425 7680 34459
rect 7622 34419 7680 34425
rect 9306 34416 9312 34468
rect 9364 34456 9370 34468
rect 9953 34459 10011 34465
rect 9953 34456 9965 34459
rect 9364 34428 9965 34456
rect 9364 34416 9370 34428
rect 9953 34425 9965 34428
rect 9999 34456 10011 34459
rect 10318 34456 10324 34468
rect 9999 34428 10324 34456
rect 9999 34425 10011 34428
rect 9953 34419 10011 34425
rect 10318 34416 10324 34428
rect 10376 34416 10382 34468
rect 14274 34416 14280 34468
rect 14332 34456 14338 34468
rect 14982 34459 15040 34465
rect 14982 34456 14994 34459
rect 14332 34428 14994 34456
rect 14332 34416 14338 34428
rect 14982 34425 14994 34428
rect 15028 34425 15040 34459
rect 17880 34456 17908 34496
rect 19429 34493 19441 34496
rect 19475 34493 19487 34527
rect 19429 34487 19487 34493
rect 19981 34527 20039 34533
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20254 34524 20260 34536
rect 20027 34496 20260 34524
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 20254 34484 20260 34496
rect 20312 34484 20318 34536
rect 20898 34484 20904 34536
rect 20956 34524 20962 34536
rect 21177 34527 21235 34533
rect 21177 34524 21189 34527
rect 20956 34496 21189 34524
rect 20956 34484 20962 34496
rect 21177 34493 21189 34496
rect 21223 34493 21235 34527
rect 21284 34524 21312 34564
rect 24305 34561 24317 34595
rect 24351 34592 24363 34595
rect 26528 34592 26556 34688
rect 24351 34564 24532 34592
rect 26528 34564 26740 34592
rect 24351 34561 24363 34564
rect 24305 34555 24363 34561
rect 21444 34527 21502 34533
rect 21444 34524 21456 34527
rect 21284 34496 21456 34524
rect 21177 34487 21235 34493
rect 21444 34493 21456 34496
rect 21490 34524 21502 34527
rect 21726 34524 21732 34536
rect 21490 34496 21732 34524
rect 21490 34493 21502 34496
rect 21444 34487 21502 34493
rect 21726 34484 21732 34496
rect 21784 34524 21790 34536
rect 21784 34496 22048 34524
rect 21784 34484 21790 34496
rect 18417 34459 18475 34465
rect 18417 34456 18429 34459
rect 17880 34428 18429 34456
rect 14982 34419 15040 34425
rect 18417 34425 18429 34428
rect 18463 34425 18475 34459
rect 18417 34419 18475 34425
rect 20073 34459 20131 34465
rect 20073 34425 20085 34459
rect 20119 34456 20131 34459
rect 20162 34456 20168 34468
rect 20119 34428 20168 34456
rect 20119 34425 20131 34428
rect 20073 34419 20131 34425
rect 20162 34416 20168 34428
rect 20220 34416 20226 34468
rect 22020 34456 22048 34496
rect 24026 34484 24032 34536
rect 24084 34524 24090 34536
rect 24397 34527 24455 34533
rect 24397 34524 24409 34527
rect 24084 34496 24409 34524
rect 24084 34484 24090 34496
rect 24397 34493 24409 34496
rect 24443 34493 24455 34527
rect 24504 34524 24532 34564
rect 24653 34527 24711 34533
rect 24653 34524 24665 34527
rect 24504 34496 24665 34524
rect 24397 34487 24455 34493
rect 24653 34493 24665 34496
rect 24699 34524 24711 34527
rect 26602 34524 26608 34536
rect 24699 34496 24808 34524
rect 26563 34496 26608 34524
rect 24699 34493 24711 34496
rect 24653 34487 24711 34493
rect 22278 34456 22284 34468
rect 22020 34428 22284 34456
rect 22278 34416 22284 34428
rect 22336 34416 22342 34468
rect 24780 34456 24808 34496
rect 26602 34484 26608 34496
rect 26660 34484 26666 34536
rect 26712 34524 26740 34564
rect 26861 34527 26919 34533
rect 26861 34524 26873 34527
rect 26712 34496 26873 34524
rect 26861 34493 26873 34496
rect 26907 34493 26919 34527
rect 26861 34487 26919 34493
rect 35345 34527 35403 34533
rect 35345 34493 35357 34527
rect 35391 34524 35403 34527
rect 35437 34527 35495 34533
rect 35437 34524 35449 34527
rect 35391 34496 35449 34524
rect 35391 34493 35403 34496
rect 35345 34487 35403 34493
rect 35437 34493 35449 34496
rect 35483 34524 35495 34527
rect 35526 34524 35532 34536
rect 35483 34496 35532 34524
rect 35483 34493 35495 34496
rect 35437 34487 35495 34493
rect 35526 34484 35532 34496
rect 35584 34484 35590 34536
rect 35710 34484 35716 34536
rect 35768 34524 35774 34536
rect 35989 34527 36047 34533
rect 35989 34524 36001 34527
rect 35768 34496 36001 34524
rect 35768 34484 35774 34496
rect 35989 34493 36001 34496
rect 36035 34493 36047 34527
rect 35989 34487 36047 34493
rect 36541 34527 36599 34533
rect 36541 34493 36553 34527
rect 36587 34524 36599 34527
rect 37090 34524 37096 34536
rect 36587 34496 37096 34524
rect 36587 34493 36599 34496
rect 36541 34487 36599 34493
rect 37090 34484 37096 34496
rect 37148 34484 37154 34536
rect 25038 34456 25044 34468
rect 24780 34428 25044 34456
rect 25038 34416 25044 34428
rect 25096 34416 25102 34468
rect 5077 34391 5135 34397
rect 5077 34357 5089 34391
rect 5123 34388 5135 34391
rect 5166 34388 5172 34400
rect 5123 34360 5172 34388
rect 5123 34357 5135 34360
rect 5077 34351 5135 34357
rect 5166 34348 5172 34360
rect 5224 34348 5230 34400
rect 5626 34348 5632 34400
rect 5684 34388 5690 34400
rect 6270 34388 6276 34400
rect 5684 34360 5729 34388
rect 6231 34360 6276 34388
rect 5684 34348 5690 34360
rect 6270 34348 6276 34360
rect 6328 34348 6334 34400
rect 7190 34388 7196 34400
rect 7151 34360 7196 34388
rect 7190 34348 7196 34360
rect 7248 34348 7254 34400
rect 9582 34388 9588 34400
rect 9543 34360 9588 34388
rect 9582 34348 9588 34360
rect 9640 34348 9646 34400
rect 11146 34388 11152 34400
rect 11107 34360 11152 34388
rect 11146 34348 11152 34360
rect 11204 34348 11210 34400
rect 28353 34391 28411 34397
rect 28353 34357 28365 34391
rect 28399 34388 28411 34391
rect 28626 34388 28632 34400
rect 28399 34360 28632 34388
rect 28399 34357 28411 34360
rect 28353 34351 28411 34357
rect 28626 34348 28632 34360
rect 28684 34348 28690 34400
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 4525 34187 4583 34193
rect 4525 34153 4537 34187
rect 4571 34184 4583 34187
rect 5626 34184 5632 34196
rect 4571 34156 5632 34184
rect 4571 34153 4583 34156
rect 4525 34147 4583 34153
rect 5626 34144 5632 34156
rect 5684 34144 5690 34196
rect 5718 34144 5724 34196
rect 5776 34184 5782 34196
rect 5997 34187 6055 34193
rect 5997 34184 6009 34187
rect 5776 34156 6009 34184
rect 5776 34144 5782 34156
rect 5997 34153 6009 34156
rect 6043 34184 6055 34187
rect 6086 34184 6092 34196
rect 6043 34156 6092 34184
rect 6043 34153 6055 34156
rect 5997 34147 6055 34153
rect 6086 34144 6092 34156
rect 6144 34144 6150 34196
rect 9125 34187 9183 34193
rect 9125 34153 9137 34187
rect 9171 34184 9183 34187
rect 9582 34184 9588 34196
rect 9171 34156 9588 34184
rect 9171 34153 9183 34156
rect 9125 34147 9183 34153
rect 1394 34076 1400 34128
rect 1452 34116 1458 34128
rect 1673 34119 1731 34125
rect 1673 34116 1685 34119
rect 1452 34088 1685 34116
rect 1452 34076 1458 34088
rect 1673 34085 1685 34088
rect 1719 34116 1731 34119
rect 2866 34116 2872 34128
rect 1719 34088 2872 34116
rect 1719 34085 1731 34088
rect 1673 34079 1731 34085
rect 2866 34076 2872 34088
rect 2924 34076 2930 34128
rect 6356 34119 6414 34125
rect 6356 34085 6368 34119
rect 6402 34116 6414 34119
rect 6638 34116 6644 34128
rect 6402 34088 6644 34116
rect 6402 34085 6414 34088
rect 6356 34079 6414 34085
rect 6638 34076 6644 34088
rect 6696 34076 6702 34128
rect 4893 34051 4951 34057
rect 4893 34017 4905 34051
rect 4939 34048 4951 34051
rect 5166 34048 5172 34060
rect 4939 34020 5172 34048
rect 4939 34017 4951 34020
rect 4893 34011 4951 34017
rect 5166 34008 5172 34020
rect 5224 34048 5230 34060
rect 5810 34048 5816 34060
rect 5224 34020 5816 34048
rect 5224 34008 5230 34020
rect 5810 34008 5816 34020
rect 5868 34008 5874 34060
rect 8481 34051 8539 34057
rect 8481 34017 8493 34051
rect 8527 34048 8539 34051
rect 9140 34048 9168 34147
rect 9582 34144 9588 34156
rect 9640 34144 9646 34196
rect 12434 34144 12440 34196
rect 12492 34184 12498 34196
rect 12986 34184 12992 34196
rect 12492 34156 12992 34184
rect 12492 34144 12498 34156
rect 12986 34144 12992 34156
rect 13044 34184 13050 34196
rect 13265 34187 13323 34193
rect 13265 34184 13277 34187
rect 13044 34156 13277 34184
rect 13044 34144 13050 34156
rect 13265 34153 13277 34156
rect 13311 34153 13323 34187
rect 13998 34184 14004 34196
rect 13959 34156 14004 34184
rect 13265 34147 13323 34153
rect 13998 34144 14004 34156
rect 14056 34144 14062 34196
rect 14093 34187 14151 34193
rect 14093 34153 14105 34187
rect 14139 34184 14151 34187
rect 14642 34184 14648 34196
rect 14139 34156 14648 34184
rect 14139 34153 14151 34156
rect 14093 34147 14151 34153
rect 14642 34144 14648 34156
rect 14700 34144 14706 34196
rect 20070 34184 20076 34196
rect 20031 34156 20076 34184
rect 20070 34144 20076 34156
rect 20128 34144 20134 34196
rect 22278 34184 22284 34196
rect 22239 34156 22284 34184
rect 22278 34144 22284 34156
rect 22336 34144 22342 34196
rect 23566 34184 23572 34196
rect 23527 34156 23572 34184
rect 23566 34144 23572 34156
rect 23624 34144 23630 34196
rect 25038 34184 25044 34196
rect 24999 34156 25044 34184
rect 25038 34144 25044 34156
rect 25096 34144 25102 34196
rect 25501 34187 25559 34193
rect 25501 34153 25513 34187
rect 25547 34184 25559 34187
rect 25774 34184 25780 34196
rect 25547 34156 25780 34184
rect 25547 34153 25559 34156
rect 25501 34147 25559 34153
rect 25774 34144 25780 34156
rect 25832 34184 25838 34196
rect 26142 34184 26148 34196
rect 25832 34156 26148 34184
rect 25832 34144 25838 34156
rect 26142 34144 26148 34156
rect 26200 34144 26206 34196
rect 35434 34144 35440 34196
rect 35492 34184 35498 34196
rect 35621 34187 35679 34193
rect 35621 34184 35633 34187
rect 35492 34156 35633 34184
rect 35492 34144 35498 34156
rect 35621 34153 35633 34156
rect 35667 34153 35679 34187
rect 35621 34147 35679 34153
rect 9493 34119 9551 34125
rect 9493 34085 9505 34119
rect 9539 34116 9551 34119
rect 9944 34119 10002 34125
rect 9944 34116 9956 34119
rect 9539 34088 9956 34116
rect 9539 34085 9551 34088
rect 9493 34079 9551 34085
rect 9944 34085 9956 34088
rect 9990 34116 10002 34119
rect 10134 34116 10140 34128
rect 9990 34088 10140 34116
rect 9990 34085 10002 34088
rect 9944 34079 10002 34085
rect 10134 34076 10140 34088
rect 10192 34076 10198 34128
rect 18040 34119 18098 34125
rect 18040 34085 18052 34119
rect 18086 34116 18098 34119
rect 18138 34116 18144 34128
rect 18086 34088 18144 34116
rect 18086 34085 18098 34088
rect 18040 34079 18098 34085
rect 18138 34076 18144 34088
rect 18196 34076 18202 34128
rect 19705 34119 19763 34125
rect 19705 34085 19717 34119
rect 19751 34116 19763 34119
rect 20162 34116 20168 34128
rect 19751 34088 20168 34116
rect 19751 34085 19763 34088
rect 19705 34079 19763 34085
rect 20162 34076 20168 34088
rect 20220 34076 20226 34128
rect 23474 34076 23480 34128
rect 23532 34116 23538 34128
rect 23906 34119 23964 34125
rect 23906 34116 23918 34119
rect 23532 34088 23918 34116
rect 23532 34076 23538 34088
rect 23906 34085 23918 34088
rect 23952 34085 23964 34119
rect 23906 34079 23964 34085
rect 24026 34076 24032 34128
rect 24084 34076 24090 34128
rect 26694 34076 26700 34128
rect 26752 34116 26758 34128
rect 27126 34119 27184 34125
rect 27126 34116 27138 34119
rect 26752 34088 27138 34116
rect 26752 34076 26758 34088
rect 27126 34085 27138 34088
rect 27172 34085 27184 34119
rect 27126 34079 27184 34085
rect 11514 34048 11520 34060
rect 8527 34020 9168 34048
rect 9692 34020 11520 34048
rect 8527 34017 8539 34020
rect 8481 34011 8539 34017
rect 4706 33940 4712 33992
rect 4764 33980 4770 33992
rect 4985 33983 5043 33989
rect 4985 33980 4997 33983
rect 4764 33952 4997 33980
rect 4764 33940 4770 33952
rect 4985 33949 4997 33952
rect 5031 33949 5043 33983
rect 4985 33943 5043 33949
rect 5077 33983 5135 33989
rect 5077 33949 5089 33983
rect 5123 33980 5135 33983
rect 5534 33980 5540 33992
rect 5123 33952 5540 33980
rect 5123 33949 5135 33952
rect 5077 33943 5135 33949
rect 3510 33872 3516 33924
rect 3568 33912 3574 33924
rect 4433 33915 4491 33921
rect 4433 33912 4445 33915
rect 3568 33884 4445 33912
rect 3568 33872 3574 33884
rect 4433 33881 4445 33884
rect 4479 33912 4491 33915
rect 5092 33912 5120 33943
rect 5534 33940 5540 33952
rect 5592 33940 5598 33992
rect 5902 33940 5908 33992
rect 5960 33980 5966 33992
rect 6089 33983 6147 33989
rect 6089 33980 6101 33983
rect 5960 33952 6101 33980
rect 5960 33940 5966 33952
rect 6089 33949 6101 33952
rect 6135 33949 6147 33983
rect 6089 33943 6147 33949
rect 9398 33940 9404 33992
rect 9456 33980 9462 33992
rect 9692 33989 9720 34020
rect 11514 34008 11520 34020
rect 11572 34008 11578 34060
rect 11790 34008 11796 34060
rect 11848 34048 11854 34060
rect 12141 34051 12199 34057
rect 12141 34048 12153 34051
rect 11848 34020 12153 34048
rect 11848 34008 11854 34020
rect 12141 34017 12153 34020
rect 12187 34017 12199 34051
rect 12141 34011 12199 34017
rect 14918 34008 14924 34060
rect 14976 34048 14982 34060
rect 15378 34048 15384 34060
rect 14976 34020 15384 34048
rect 14976 34008 14982 34020
rect 15378 34008 15384 34020
rect 15436 34048 15442 34060
rect 15545 34051 15603 34057
rect 15545 34048 15557 34051
rect 15436 34020 15557 34048
rect 15436 34008 15442 34020
rect 15545 34017 15557 34020
rect 15591 34017 15603 34051
rect 15545 34011 15603 34017
rect 20990 34008 20996 34060
rect 21048 34048 21054 34060
rect 21157 34051 21215 34057
rect 21157 34048 21169 34051
rect 21048 34020 21169 34048
rect 21048 34008 21054 34020
rect 21157 34017 21169 34020
rect 21203 34017 21215 34051
rect 21157 34011 21215 34017
rect 22649 34051 22707 34057
rect 22649 34017 22661 34051
rect 22695 34048 22707 34051
rect 22738 34048 22744 34060
rect 22695 34020 22744 34048
rect 22695 34017 22707 34020
rect 22649 34011 22707 34017
rect 22738 34008 22744 34020
rect 22796 34048 22802 34060
rect 23661 34051 23719 34057
rect 23661 34048 23673 34051
rect 22796 34020 23673 34048
rect 22796 34008 22802 34020
rect 23661 34017 23673 34020
rect 23707 34048 23719 34051
rect 24044 34048 24072 34076
rect 23707 34020 24072 34048
rect 23707 34017 23719 34020
rect 23661 34011 23719 34017
rect 35250 34008 35256 34060
rect 35308 34048 35314 34060
rect 35437 34051 35495 34057
rect 35437 34048 35449 34051
rect 35308 34020 35449 34048
rect 35308 34008 35314 34020
rect 35437 34017 35449 34020
rect 35483 34017 35495 34051
rect 35437 34011 35495 34017
rect 9677 33983 9735 33989
rect 9677 33980 9689 33983
rect 9456 33952 9689 33980
rect 9456 33940 9462 33952
rect 9677 33949 9689 33952
rect 9723 33949 9735 33983
rect 11532 33980 11560 34008
rect 11885 33983 11943 33989
rect 11885 33980 11897 33983
rect 11532 33952 11897 33980
rect 9677 33943 9735 33949
rect 11885 33949 11897 33952
rect 11931 33949 11943 33983
rect 11885 33943 11943 33949
rect 14734 33940 14740 33992
rect 14792 33980 14798 33992
rect 15289 33983 15347 33989
rect 15289 33980 15301 33983
rect 14792 33952 15301 33980
rect 14792 33940 14798 33952
rect 15289 33949 15301 33952
rect 15335 33949 15347 33983
rect 15289 33943 15347 33949
rect 17773 33983 17831 33989
rect 17773 33949 17785 33983
rect 17819 33949 17831 33983
rect 17773 33943 17831 33949
rect 4479 33884 5120 33912
rect 4479 33881 4491 33884
rect 4433 33875 4491 33881
rect 2958 33844 2964 33856
rect 2919 33816 2964 33844
rect 2958 33804 2964 33816
rect 3016 33804 3022 33856
rect 3881 33847 3939 33853
rect 3881 33813 3893 33847
rect 3927 33844 3939 33847
rect 4062 33844 4068 33856
rect 3927 33816 4068 33844
rect 3927 33813 3939 33816
rect 3881 33807 3939 33813
rect 4062 33804 4068 33816
rect 4120 33804 4126 33856
rect 7190 33804 7196 33856
rect 7248 33844 7254 33856
rect 7469 33847 7527 33853
rect 7469 33844 7481 33847
rect 7248 33816 7481 33844
rect 7248 33804 7254 33816
rect 7469 33813 7481 33816
rect 7515 33813 7527 33847
rect 8662 33844 8668 33856
rect 8623 33816 8668 33844
rect 7469 33807 7527 33813
rect 8662 33804 8668 33816
rect 8720 33804 8726 33856
rect 11054 33844 11060 33856
rect 11015 33816 11060 33844
rect 11054 33804 11060 33816
rect 11112 33804 11118 33856
rect 14274 33804 14280 33856
rect 14332 33844 14338 33856
rect 14737 33847 14795 33853
rect 14737 33844 14749 33847
rect 14332 33816 14749 33844
rect 14332 33804 14338 33816
rect 14737 33813 14749 33816
rect 14783 33813 14795 33847
rect 15304 33844 15332 33943
rect 17788 33912 17816 33943
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 20898 33980 20904 33992
rect 20680 33952 20904 33980
rect 20680 33940 20686 33952
rect 20898 33940 20904 33952
rect 20956 33940 20962 33992
rect 26602 33940 26608 33992
rect 26660 33980 26666 33992
rect 26881 33983 26939 33989
rect 26881 33980 26893 33983
rect 26660 33952 26893 33980
rect 26660 33940 26666 33952
rect 16224 33884 17816 33912
rect 16224 33856 16252 33884
rect 26804 33856 26832 33952
rect 26881 33949 26893 33952
rect 26927 33949 26939 33983
rect 26881 33943 26939 33949
rect 16206 33844 16212 33856
rect 15304 33816 16212 33844
rect 14737 33807 14795 33813
rect 16206 33804 16212 33816
rect 16264 33804 16270 33856
rect 16666 33844 16672 33856
rect 16627 33816 16672 33844
rect 16666 33804 16672 33816
rect 16724 33804 16730 33856
rect 17034 33844 17040 33856
rect 16995 33816 17040 33844
rect 17034 33804 17040 33816
rect 17092 33804 17098 33856
rect 17310 33804 17316 33856
rect 17368 33844 17374 33856
rect 17405 33847 17463 33853
rect 17405 33844 17417 33847
rect 17368 33816 17417 33844
rect 17368 33804 17374 33816
rect 17405 33813 17417 33816
rect 17451 33844 17463 33847
rect 17770 33844 17776 33856
rect 17451 33816 17776 33844
rect 17451 33813 17463 33816
rect 17405 33807 17463 33813
rect 17770 33804 17776 33816
rect 17828 33804 17834 33856
rect 19150 33844 19156 33856
rect 19111 33816 19156 33844
rect 19150 33804 19156 33816
rect 19208 33804 19214 33856
rect 25866 33844 25872 33856
rect 25827 33816 25872 33844
rect 25866 33804 25872 33816
rect 25924 33844 25930 33856
rect 26234 33844 26240 33856
rect 25924 33816 26240 33844
rect 25924 33804 25930 33816
rect 26234 33804 26240 33816
rect 26292 33804 26298 33856
rect 26786 33844 26792 33856
rect 26747 33816 26792 33844
rect 26786 33804 26792 33816
rect 26844 33804 26850 33856
rect 28258 33844 28264 33856
rect 28219 33816 28264 33844
rect 28258 33804 28264 33816
rect 28316 33804 28322 33856
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 5810 33640 5816 33652
rect 5723 33612 5816 33640
rect 5810 33600 5816 33612
rect 5868 33640 5874 33652
rect 6089 33643 6147 33649
rect 6089 33640 6101 33643
rect 5868 33612 6101 33640
rect 5868 33600 5874 33612
rect 6089 33609 6101 33612
rect 6135 33609 6147 33643
rect 6089 33603 6147 33609
rect 6270 33600 6276 33652
rect 6328 33640 6334 33652
rect 6825 33643 6883 33649
rect 6825 33640 6837 33643
rect 6328 33612 6837 33640
rect 6328 33600 6334 33612
rect 6825 33609 6837 33612
rect 6871 33609 6883 33643
rect 6825 33603 6883 33609
rect 9953 33643 10011 33649
rect 9953 33609 9965 33643
rect 9999 33640 10011 33643
rect 10134 33640 10140 33652
rect 9999 33612 10140 33640
rect 9999 33609 10011 33612
rect 9953 33603 10011 33609
rect 10134 33600 10140 33612
rect 10192 33640 10198 33652
rect 10229 33643 10287 33649
rect 10229 33640 10241 33643
rect 10192 33612 10241 33640
rect 10192 33600 10198 33612
rect 10229 33609 10241 33612
rect 10275 33609 10287 33643
rect 10229 33603 10287 33609
rect 15105 33643 15163 33649
rect 15105 33609 15117 33643
rect 15151 33640 15163 33643
rect 15930 33640 15936 33652
rect 15151 33612 15936 33640
rect 15151 33609 15163 33612
rect 15105 33603 15163 33609
rect 15930 33600 15936 33612
rect 15988 33600 15994 33652
rect 17034 33600 17040 33652
rect 17092 33640 17098 33652
rect 17865 33643 17923 33649
rect 17865 33640 17877 33643
rect 17092 33612 17877 33640
rect 17092 33600 17098 33612
rect 17865 33609 17877 33612
rect 17911 33640 17923 33643
rect 18322 33640 18328 33652
rect 17911 33612 18328 33640
rect 17911 33609 17923 33612
rect 17865 33603 17923 33609
rect 18322 33600 18328 33612
rect 18380 33640 18386 33652
rect 19242 33640 19248 33652
rect 18380 33612 19248 33640
rect 18380 33600 18386 33612
rect 19242 33600 19248 33612
rect 19300 33600 19306 33652
rect 20165 33643 20223 33649
rect 20165 33609 20177 33643
rect 20211 33640 20223 33643
rect 20990 33640 20996 33652
rect 20211 33612 20996 33640
rect 20211 33609 20223 33612
rect 20165 33603 20223 33609
rect 20990 33600 20996 33612
rect 21048 33640 21054 33652
rect 22005 33643 22063 33649
rect 22005 33640 22017 33643
rect 21048 33612 22017 33640
rect 21048 33600 21054 33612
rect 22005 33609 22017 33612
rect 22051 33609 22063 33643
rect 22005 33603 22063 33609
rect 22373 33643 22431 33649
rect 22373 33609 22385 33643
rect 22419 33640 22431 33643
rect 22738 33640 22744 33652
rect 22419 33612 22744 33640
rect 22419 33609 22431 33612
rect 22373 33603 22431 33609
rect 6549 33575 6607 33581
rect 6549 33541 6561 33575
rect 6595 33572 6607 33575
rect 6638 33572 6644 33584
rect 6595 33544 6644 33572
rect 6595 33541 6607 33544
rect 6549 33535 6607 33541
rect 6638 33532 6644 33544
rect 6696 33532 6702 33584
rect 10778 33572 10784 33584
rect 10739 33544 10784 33572
rect 10778 33532 10784 33544
rect 10836 33532 10842 33584
rect 2409 33507 2467 33513
rect 2409 33473 2421 33507
rect 2455 33504 2467 33507
rect 3510 33504 3516 33516
rect 2455 33476 3516 33504
rect 2455 33473 2467 33476
rect 2409 33467 2467 33473
rect 3510 33464 3516 33476
rect 3568 33464 3574 33516
rect 7374 33504 7380 33516
rect 7335 33476 7380 33504
rect 7374 33464 7380 33476
rect 7432 33464 7438 33516
rect 8481 33507 8539 33513
rect 8481 33473 8493 33507
rect 8527 33504 8539 33507
rect 8527 33476 8708 33504
rect 8527 33473 8539 33476
rect 8481 33467 8539 33473
rect 2958 33396 2964 33448
rect 3016 33436 3022 33448
rect 3237 33439 3295 33445
rect 3237 33436 3249 33439
rect 3016 33408 3249 33436
rect 3016 33396 3022 33408
rect 3237 33405 3249 33408
rect 3283 33405 3295 33439
rect 3237 33399 3295 33405
rect 4062 33396 4068 33448
rect 4120 33436 4126 33448
rect 4433 33439 4491 33445
rect 4433 33436 4445 33439
rect 4120 33408 4445 33436
rect 4120 33396 4126 33408
rect 4433 33405 4445 33408
rect 4479 33436 4491 33439
rect 5902 33436 5908 33448
rect 4479 33408 5908 33436
rect 4479 33405 4491 33408
rect 4433 33399 4491 33405
rect 5902 33396 5908 33408
rect 5960 33396 5966 33448
rect 6822 33396 6828 33448
rect 6880 33436 6886 33448
rect 7392 33436 7420 33464
rect 6880 33408 7420 33436
rect 6880 33396 6886 33408
rect 8386 33396 8392 33448
rect 8444 33436 8450 33448
rect 8573 33439 8631 33445
rect 8573 33436 8585 33439
rect 8444 33408 8585 33436
rect 8444 33396 8450 33408
rect 8573 33405 8585 33408
rect 8619 33405 8631 33439
rect 8680 33436 8708 33476
rect 11054 33464 11060 33516
rect 11112 33504 11118 33516
rect 11333 33507 11391 33513
rect 11333 33504 11345 33507
rect 11112 33476 11345 33504
rect 11112 33464 11118 33476
rect 11333 33473 11345 33476
rect 11379 33504 11391 33507
rect 11790 33504 11796 33516
rect 11379 33476 11796 33504
rect 11379 33473 11391 33476
rect 11333 33467 11391 33473
rect 11790 33464 11796 33476
rect 11848 33464 11854 33516
rect 12986 33504 12992 33516
rect 12947 33476 12992 33504
rect 12986 33464 12992 33476
rect 13044 33504 13050 33516
rect 13449 33507 13507 33513
rect 13449 33504 13461 33507
rect 13044 33476 13461 33504
rect 13044 33464 13050 33476
rect 13449 33473 13461 33476
rect 13495 33473 13507 33507
rect 13449 33467 13507 33473
rect 15102 33464 15108 33516
rect 15160 33504 15166 33516
rect 15660 33507 15718 33513
rect 15660 33504 15672 33507
rect 15160 33476 15672 33504
rect 15160 33464 15166 33476
rect 15660 33473 15672 33476
rect 15706 33473 15718 33507
rect 15930 33504 15936 33516
rect 15891 33476 15936 33504
rect 15660 33467 15718 33473
rect 15930 33464 15936 33476
rect 15988 33464 15994 33516
rect 22388 33504 22416 33603
rect 22738 33600 22744 33612
rect 22796 33600 22802 33652
rect 23474 33640 23480 33652
rect 23435 33612 23480 33640
rect 23474 33600 23480 33612
rect 23532 33600 23538 33652
rect 25038 33600 25044 33652
rect 25096 33640 25102 33652
rect 25225 33643 25283 33649
rect 25225 33640 25237 33643
rect 25096 33612 25237 33640
rect 25096 33600 25102 33612
rect 25225 33609 25237 33612
rect 25271 33609 25283 33643
rect 25225 33603 25283 33609
rect 23109 33575 23167 33581
rect 23109 33541 23121 33575
rect 23155 33572 23167 33575
rect 24118 33572 24124 33584
rect 23155 33544 24124 33572
rect 23155 33541 23167 33544
rect 23109 33535 23167 33541
rect 21652 33476 22416 33504
rect 8846 33445 8852 33448
rect 8840 33436 8852 33445
rect 8680 33408 8852 33436
rect 8573 33399 8631 33405
rect 8840 33399 8852 33408
rect 8846 33396 8852 33399
rect 8904 33396 8910 33448
rect 10689 33439 10747 33445
rect 10689 33405 10701 33439
rect 10735 33436 10747 33439
rect 11146 33436 11152 33448
rect 10735 33408 11152 33436
rect 10735 33405 10747 33408
rect 10689 33399 10747 33405
rect 11146 33396 11152 33408
rect 11204 33396 11210 33448
rect 11238 33396 11244 33448
rect 11296 33436 11302 33448
rect 12802 33436 12808 33448
rect 11296 33408 11341 33436
rect 12763 33408 12808 33436
rect 11296 33396 11302 33408
rect 12802 33396 12808 33408
rect 12860 33396 12866 33448
rect 15562 33445 15568 33448
rect 14093 33439 14151 33445
rect 14093 33405 14105 33439
rect 14139 33436 14151 33439
rect 14921 33439 14979 33445
rect 14921 33436 14933 33439
rect 14139 33408 14933 33436
rect 14139 33405 14151 33408
rect 14093 33399 14151 33405
rect 14921 33405 14933 33408
rect 14967 33436 14979 33439
rect 15197 33439 15255 33445
rect 15197 33436 15209 33439
rect 14967 33408 15209 33436
rect 14967 33405 14979 33408
rect 14921 33399 14979 33405
rect 15197 33405 15209 33408
rect 15243 33405 15255 33439
rect 15520 33439 15568 33445
rect 15520 33436 15532 33439
rect 15197 33399 15255 33405
rect 15304 33408 15532 33436
rect 4706 33377 4712 33380
rect 2777 33371 2835 33377
rect 2777 33337 2789 33371
rect 2823 33368 2835 33371
rect 3973 33371 4031 33377
rect 2823 33340 3372 33368
rect 2823 33337 2835 33340
rect 2777 33331 2835 33337
rect 3344 33312 3372 33340
rect 3973 33337 3985 33371
rect 4019 33368 4031 33371
rect 4341 33371 4399 33377
rect 4341 33368 4353 33371
rect 4019 33340 4353 33368
rect 4019 33337 4031 33340
rect 3973 33331 4031 33337
rect 4341 33337 4353 33340
rect 4387 33368 4399 33371
rect 4700 33368 4712 33377
rect 4387 33340 4712 33368
rect 4387 33337 4399 33340
rect 4341 33331 4399 33337
rect 4700 33331 4712 33340
rect 4706 33328 4712 33331
rect 4764 33328 4770 33380
rect 6638 33328 6644 33380
rect 6696 33368 6702 33380
rect 7285 33371 7343 33377
rect 7285 33368 7297 33371
rect 6696 33340 7297 33368
rect 6696 33328 6702 33340
rect 7285 33337 7297 33340
rect 7331 33368 7343 33371
rect 7837 33371 7895 33377
rect 7837 33368 7849 33371
rect 7331 33340 7849 33368
rect 7331 33337 7343 33340
rect 7285 33331 7343 33337
rect 7837 33337 7849 33340
rect 7883 33337 7895 33371
rect 7837 33331 7895 33337
rect 12253 33371 12311 33377
rect 12253 33337 12265 33371
rect 12299 33368 12311 33371
rect 12894 33368 12900 33380
rect 12299 33340 12900 33368
rect 12299 33337 12311 33340
rect 12253 33331 12311 33337
rect 12894 33328 12900 33340
rect 12952 33328 12958 33380
rect 14737 33371 14795 33377
rect 14737 33337 14749 33371
rect 14783 33368 14795 33371
rect 15304 33368 15332 33408
rect 15520 33405 15532 33408
rect 15566 33405 15568 33439
rect 15520 33399 15568 33405
rect 15562 33396 15568 33399
rect 15620 33436 15626 33448
rect 18049 33439 18107 33445
rect 15620 33408 15668 33436
rect 15620 33396 15626 33408
rect 18049 33405 18061 33439
rect 18095 33436 18107 33439
rect 18095 33408 19840 33436
rect 18095 33405 18107 33408
rect 18049 33399 18107 33405
rect 18322 33377 18328 33380
rect 14783 33340 15332 33368
rect 14783 33337 14795 33340
rect 14737 33331 14795 33337
rect 18316 33331 18328 33377
rect 18380 33368 18386 33380
rect 18380 33340 18416 33368
rect 18322 33328 18328 33331
rect 18380 33328 18386 33340
rect 1762 33300 1768 33312
rect 1723 33272 1768 33300
rect 1762 33260 1768 33272
rect 1820 33260 1826 33312
rect 2866 33300 2872 33312
rect 2827 33272 2872 33300
rect 2866 33260 2872 33272
rect 2924 33260 2930 33312
rect 3326 33300 3332 33312
rect 3287 33272 3332 33300
rect 3326 33260 3332 33272
rect 3384 33260 3390 33312
rect 7190 33300 7196 33312
rect 7151 33272 7196 33300
rect 7190 33260 7196 33272
rect 7248 33260 7254 33312
rect 12158 33260 12164 33312
rect 12216 33300 12222 33312
rect 12437 33303 12495 33309
rect 12437 33300 12449 33303
rect 12216 33272 12449 33300
rect 12216 33260 12222 33272
rect 12437 33269 12449 33272
rect 12483 33269 12495 33303
rect 14182 33300 14188 33312
rect 14143 33272 14188 33300
rect 12437 33263 12495 33269
rect 14182 33260 14188 33272
rect 14240 33260 14246 33312
rect 14921 33303 14979 33309
rect 14921 33269 14933 33303
rect 14967 33300 14979 33303
rect 15286 33300 15292 33312
rect 14967 33272 15292 33300
rect 14967 33269 14979 33272
rect 14921 33263 14979 33269
rect 15286 33260 15292 33272
rect 15344 33260 15350 33312
rect 17034 33300 17040 33312
rect 16995 33272 17040 33300
rect 17034 33260 17040 33272
rect 17092 33260 17098 33312
rect 17497 33303 17555 33309
rect 17497 33269 17509 33303
rect 17543 33300 17555 33303
rect 18138 33300 18144 33312
rect 17543 33272 18144 33300
rect 17543 33269 17555 33272
rect 17497 33263 17555 33269
rect 18138 33260 18144 33272
rect 18196 33300 18202 33312
rect 19812 33309 19840 33408
rect 20162 33396 20168 33448
rect 20220 33436 20226 33448
rect 20622 33436 20628 33448
rect 20220 33408 20628 33436
rect 20220 33396 20226 33408
rect 20622 33396 20628 33408
rect 20680 33436 20686 33448
rect 21652 33436 21680 33476
rect 20680 33408 21680 33436
rect 20680 33396 20686 33408
rect 21818 33396 21824 33448
rect 21876 33436 21882 33448
rect 23124 33436 23152 33535
rect 24118 33532 24124 33544
rect 24176 33532 24182 33584
rect 23566 33464 23572 33516
rect 23624 33504 23630 33516
rect 24213 33507 24271 33513
rect 24213 33504 24225 33507
rect 23624 33476 24225 33504
rect 23624 33464 23630 33476
rect 24213 33473 24225 33476
rect 24259 33504 24271 33507
rect 24670 33504 24676 33516
rect 24259 33476 24676 33504
rect 24259 33473 24271 33476
rect 24213 33467 24271 33473
rect 24670 33464 24676 33476
rect 24728 33464 24734 33516
rect 21876 33408 23152 33436
rect 21876 33396 21882 33408
rect 23382 33396 23388 33448
rect 23440 33436 23446 33448
rect 23440 33408 24256 33436
rect 23440 33396 23446 33408
rect 20533 33371 20591 33377
rect 20533 33337 20545 33371
rect 20579 33368 20591 33371
rect 20892 33371 20950 33377
rect 20892 33368 20904 33371
rect 20579 33340 20904 33368
rect 20579 33337 20591 33340
rect 20533 33331 20591 33337
rect 20892 33337 20904 33340
rect 20938 33368 20950 33371
rect 21910 33368 21916 33380
rect 20938 33340 21916 33368
rect 20938 33337 20950 33340
rect 20892 33331 20950 33337
rect 21910 33328 21916 33340
rect 21968 33328 21974 33380
rect 24118 33368 24124 33380
rect 24079 33340 24124 33368
rect 24118 33328 24124 33340
rect 24176 33328 24182 33380
rect 19429 33303 19487 33309
rect 19429 33300 19441 33303
rect 18196 33272 19441 33300
rect 18196 33260 18202 33272
rect 19429 33269 19441 33272
rect 19475 33269 19487 33303
rect 19429 33263 19487 33269
rect 19797 33303 19855 33309
rect 19797 33269 19809 33303
rect 19843 33300 19855 33303
rect 19978 33300 19984 33312
rect 19843 33272 19984 33300
rect 19843 33269 19855 33272
rect 19797 33263 19855 33269
rect 19978 33260 19984 33272
rect 20036 33260 20042 33312
rect 23474 33260 23480 33312
rect 23532 33300 23538 33312
rect 23661 33303 23719 33309
rect 23661 33300 23673 33303
rect 23532 33272 23673 33300
rect 23532 33260 23538 33272
rect 23661 33269 23673 33272
rect 23707 33269 23719 33303
rect 23661 33263 23719 33269
rect 24029 33303 24087 33309
rect 24029 33269 24041 33303
rect 24075 33300 24087 33303
rect 24228 33300 24256 33408
rect 25240 33368 25268 33603
rect 25314 33600 25320 33652
rect 25372 33640 25378 33652
rect 25409 33643 25467 33649
rect 25409 33640 25421 33643
rect 25372 33612 25421 33640
rect 25372 33600 25378 33612
rect 25409 33609 25421 33612
rect 25455 33609 25467 33643
rect 25409 33603 25467 33609
rect 26694 33600 26700 33652
rect 26752 33640 26758 33652
rect 26789 33643 26847 33649
rect 26789 33640 26801 33643
rect 26752 33612 26801 33640
rect 26752 33600 26758 33612
rect 26789 33609 26801 33612
rect 26835 33609 26847 33643
rect 35618 33640 35624 33652
rect 35579 33612 35624 33640
rect 26789 33603 26847 33609
rect 35618 33600 35624 33612
rect 35676 33600 35682 33652
rect 25958 33504 25964 33516
rect 25919 33476 25964 33504
rect 25958 33464 25964 33476
rect 26016 33464 26022 33516
rect 35250 33464 35256 33516
rect 35308 33504 35314 33516
rect 35989 33507 36047 33513
rect 35989 33504 36001 33507
rect 35308 33476 36001 33504
rect 35308 33464 35314 33476
rect 35989 33473 36001 33476
rect 36035 33473 36047 33507
rect 35989 33467 36047 33473
rect 25774 33436 25780 33448
rect 25735 33408 25780 33436
rect 25774 33396 25780 33408
rect 25832 33396 25838 33448
rect 26513 33439 26571 33445
rect 26513 33405 26525 33439
rect 26559 33436 26571 33439
rect 26786 33436 26792 33448
rect 26559 33408 26792 33436
rect 26559 33405 26571 33408
rect 26513 33399 26571 33405
rect 26786 33396 26792 33408
rect 26844 33436 26850 33448
rect 26973 33439 27031 33445
rect 26973 33436 26985 33439
rect 26844 33408 26985 33436
rect 26844 33396 26850 33408
rect 26973 33405 26985 33408
rect 27019 33405 27031 33439
rect 26973 33399 27031 33405
rect 25869 33371 25927 33377
rect 25869 33368 25881 33371
rect 25240 33340 25881 33368
rect 25869 33337 25881 33340
rect 25915 33337 25927 33371
rect 26988 33368 27016 33399
rect 27062 33396 27068 33448
rect 27120 33436 27126 33448
rect 27240 33439 27298 33445
rect 27240 33436 27252 33439
rect 27120 33408 27252 33436
rect 27120 33396 27126 33408
rect 27240 33405 27252 33408
rect 27286 33436 27298 33439
rect 28258 33436 28264 33448
rect 27286 33408 28264 33436
rect 27286 33405 27298 33408
rect 27240 33399 27298 33405
rect 28258 33396 28264 33408
rect 28316 33396 28322 33448
rect 35437 33439 35495 33445
rect 35437 33436 35449 33439
rect 35360 33408 35449 33436
rect 27154 33368 27160 33380
rect 26988 33340 27160 33368
rect 25869 33331 25927 33337
rect 27154 33328 27160 33340
rect 27212 33328 27218 33380
rect 35360 33312 35388 33408
rect 35437 33405 35449 33408
rect 35483 33405 35495 33439
rect 35437 33399 35495 33405
rect 24673 33303 24731 33309
rect 24673 33300 24685 33303
rect 24075 33272 24685 33300
rect 24075 33269 24087 33272
rect 24029 33263 24087 33269
rect 24673 33269 24685 33272
rect 24719 33269 24731 33303
rect 28350 33300 28356 33312
rect 28311 33272 28356 33300
rect 24673 33263 24731 33269
rect 28350 33260 28356 33272
rect 28408 33260 28414 33312
rect 28626 33300 28632 33312
rect 28587 33272 28632 33300
rect 28626 33260 28632 33272
rect 28684 33260 28690 33312
rect 35342 33300 35348 33312
rect 35303 33272 35348 33300
rect 35342 33260 35348 33272
rect 35400 33260 35406 33312
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 3786 33096 3792 33108
rect 2924 33068 3792 33096
rect 2924 33056 2930 33068
rect 3786 33056 3792 33068
rect 3844 33056 3850 33108
rect 4706 33056 4712 33108
rect 4764 33096 4770 33108
rect 5445 33099 5503 33105
rect 5445 33096 5457 33099
rect 4764 33068 5457 33096
rect 4764 33056 4770 33068
rect 5445 33065 5457 33068
rect 5491 33065 5503 33099
rect 5445 33059 5503 33065
rect 5534 33056 5540 33108
rect 5592 33096 5598 33108
rect 6457 33099 6515 33105
rect 6457 33096 6469 33099
rect 5592 33068 6469 33096
rect 5592 33056 5598 33068
rect 6457 33065 6469 33068
rect 6503 33096 6515 33099
rect 6822 33096 6828 33108
rect 6503 33068 6828 33096
rect 6503 33065 6515 33068
rect 6457 33059 6515 33065
rect 6822 33056 6828 33068
rect 6880 33056 6886 33108
rect 7190 33056 7196 33108
rect 7248 33096 7254 33108
rect 7561 33099 7619 33105
rect 7561 33096 7573 33099
rect 7248 33068 7573 33096
rect 7248 33056 7254 33068
rect 7561 33065 7573 33068
rect 7607 33065 7619 33099
rect 7561 33059 7619 33065
rect 8386 33056 8392 33108
rect 8444 33056 8450 33108
rect 8662 33056 8668 33108
rect 8720 33096 8726 33108
rect 9033 33099 9091 33105
rect 9033 33096 9045 33099
rect 8720 33068 9045 33096
rect 8720 33056 8726 33068
rect 9033 33065 9045 33068
rect 9079 33065 9091 33099
rect 9033 33059 9091 33065
rect 10873 33099 10931 33105
rect 10873 33065 10885 33099
rect 10919 33096 10931 33099
rect 10962 33096 10968 33108
rect 10919 33068 10968 33096
rect 10919 33065 10931 33068
rect 10873 33059 10931 33065
rect 10962 33056 10968 33068
rect 11020 33056 11026 33108
rect 11238 33096 11244 33108
rect 11199 33068 11244 33096
rect 11238 33056 11244 33068
rect 11296 33056 11302 33108
rect 12158 33056 12164 33108
rect 12216 33096 12222 33108
rect 12345 33099 12403 33105
rect 12345 33096 12357 33099
rect 12216 33068 12357 33096
rect 12216 33056 12222 33068
rect 12345 33065 12357 33068
rect 12391 33065 12403 33099
rect 12345 33059 12403 33065
rect 12802 33056 12808 33108
rect 12860 33096 12866 33108
rect 12897 33099 12955 33105
rect 12897 33096 12909 33099
rect 12860 33068 12909 33096
rect 12860 33056 12866 33068
rect 12897 33065 12909 33068
rect 12943 33065 12955 33099
rect 13630 33096 13636 33108
rect 13591 33068 13636 33096
rect 12897 33059 12955 33065
rect 13630 33056 13636 33068
rect 13688 33056 13694 33108
rect 14737 33099 14795 33105
rect 14737 33065 14749 33099
rect 14783 33096 14795 33099
rect 14918 33096 14924 33108
rect 14783 33068 14924 33096
rect 14783 33065 14795 33068
rect 14737 33059 14795 33065
rect 14918 33056 14924 33068
rect 14976 33056 14982 33108
rect 15102 33096 15108 33108
rect 15063 33068 15108 33096
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 19334 33056 19340 33108
rect 19392 33096 19398 33108
rect 19392 33068 19437 33096
rect 19392 33056 19398 33068
rect 22094 33056 22100 33108
rect 22152 33096 22158 33108
rect 22281 33099 22339 33105
rect 22281 33096 22293 33099
rect 22152 33068 22293 33096
rect 22152 33056 22158 33068
rect 22281 33065 22293 33068
rect 22327 33096 22339 33099
rect 23477 33099 23535 33105
rect 23477 33096 23489 33099
rect 22327 33068 23489 33096
rect 22327 33065 22339 33068
rect 22281 33059 22339 33065
rect 23477 33065 23489 33068
rect 23523 33065 23535 33099
rect 24670 33096 24676 33108
rect 24631 33068 24676 33096
rect 23477 33059 23535 33065
rect 24670 33056 24676 33068
rect 24728 33056 24734 33108
rect 24854 33096 24860 33108
rect 24815 33068 24860 33096
rect 24854 33056 24860 33068
rect 24912 33056 24918 33108
rect 27062 33096 27068 33108
rect 27023 33068 27068 33096
rect 27062 33056 27068 33068
rect 27120 33056 27126 33108
rect 5902 32988 5908 33040
rect 5960 33028 5966 33040
rect 5997 33031 6055 33037
rect 5997 33028 6009 33031
rect 5960 33000 6009 33028
rect 5960 32988 5966 33000
rect 5997 32997 6009 33000
rect 6043 32997 6055 33031
rect 8404 33028 8432 33056
rect 9398 33028 9404 33040
rect 8404 33000 9404 33028
rect 5997 32991 6055 32997
rect 9398 32988 9404 33000
rect 9456 33028 9462 33040
rect 10229 33031 10287 33037
rect 10229 33028 10241 33031
rect 9456 33000 10241 33028
rect 9456 32988 9462 33000
rect 10229 32997 10241 33000
rect 10275 32997 10287 33031
rect 12250 33028 12256 33040
rect 12211 33000 12256 33028
rect 10229 32991 10287 32997
rect 12250 32988 12256 33000
rect 12308 32988 12314 33040
rect 24688 33028 24716 33056
rect 27424 33031 27482 33037
rect 24688 33000 25452 33028
rect 1854 32920 1860 32972
rect 1912 32960 1918 32972
rect 2021 32963 2079 32969
rect 2021 32960 2033 32963
rect 1912 32932 2033 32960
rect 1912 32920 1918 32932
rect 2021 32929 2033 32932
rect 2067 32960 2079 32963
rect 3326 32960 3332 32972
rect 2067 32932 3332 32960
rect 2067 32929 2079 32932
rect 2021 32923 2079 32929
rect 3326 32920 3332 32932
rect 3384 32920 3390 32972
rect 4321 32963 4379 32969
rect 4321 32960 4333 32963
rect 3988 32932 4333 32960
rect 1762 32892 1768 32904
rect 1596 32864 1768 32892
rect 1394 32716 1400 32768
rect 1452 32756 1458 32768
rect 1596 32765 1624 32864
rect 1762 32852 1768 32864
rect 1820 32852 1826 32904
rect 2958 32784 2964 32836
rect 3016 32824 3022 32836
rect 3145 32827 3203 32833
rect 3145 32824 3157 32827
rect 3016 32796 3157 32824
rect 3016 32784 3022 32796
rect 3145 32793 3157 32796
rect 3191 32824 3203 32827
rect 3988 32824 4016 32932
rect 4321 32929 4333 32932
rect 4367 32929 4379 32963
rect 4321 32923 4379 32929
rect 6917 32963 6975 32969
rect 6917 32929 6929 32963
rect 6963 32960 6975 32963
rect 7282 32960 7288 32972
rect 6963 32932 7288 32960
rect 6963 32929 6975 32932
rect 6917 32923 6975 32929
rect 7282 32920 7288 32932
rect 7340 32920 7346 32972
rect 8386 32920 8392 32972
rect 8444 32960 8450 32972
rect 8481 32963 8539 32969
rect 8481 32960 8493 32963
rect 8444 32932 8493 32960
rect 8444 32920 8450 32932
rect 8481 32929 8493 32932
rect 8527 32929 8539 32963
rect 9674 32960 9680 32972
rect 9635 32932 9680 32960
rect 8481 32923 8539 32929
rect 9674 32920 9680 32932
rect 9732 32920 9738 32972
rect 13262 32920 13268 32972
rect 13320 32960 13326 32972
rect 14001 32963 14059 32969
rect 14001 32960 14013 32963
rect 13320 32932 14013 32960
rect 13320 32920 13326 32932
rect 14001 32929 14013 32932
rect 14047 32929 14059 32963
rect 15286 32960 15292 32972
rect 15247 32932 15292 32960
rect 14001 32923 14059 32929
rect 15286 32920 15292 32932
rect 15344 32920 15350 32972
rect 15562 32920 15568 32972
rect 15620 32969 15626 32972
rect 15620 32963 15670 32969
rect 15620 32929 15624 32963
rect 15658 32929 15670 32963
rect 16022 32960 16028 32972
rect 15983 32932 16028 32960
rect 15620 32923 15670 32929
rect 15620 32920 15626 32923
rect 16022 32920 16028 32932
rect 16080 32920 16086 32972
rect 18230 32969 18236 32972
rect 18224 32960 18236 32969
rect 18191 32932 18236 32960
rect 18224 32923 18236 32932
rect 18230 32920 18236 32923
rect 18288 32920 18294 32972
rect 20622 32920 20628 32972
rect 20680 32960 20686 32972
rect 21157 32963 21215 32969
rect 21157 32960 21169 32963
rect 20680 32932 21169 32960
rect 20680 32920 20686 32932
rect 21157 32929 21169 32932
rect 21203 32929 21215 32963
rect 21157 32923 21215 32929
rect 22922 32920 22928 32972
rect 22980 32960 22986 32972
rect 25222 32960 25228 32972
rect 22980 32932 23704 32960
rect 25183 32932 25228 32960
rect 22980 32920 22986 32932
rect 4062 32852 4068 32904
rect 4120 32892 4126 32904
rect 4120 32864 4213 32892
rect 4120 32852 4126 32864
rect 6270 32852 6276 32904
rect 6328 32892 6334 32904
rect 7009 32895 7067 32901
rect 7009 32892 7021 32895
rect 6328 32864 7021 32892
rect 6328 32852 6334 32864
rect 7009 32861 7021 32864
rect 7055 32861 7067 32895
rect 7009 32855 7067 32861
rect 7193 32895 7251 32901
rect 7193 32861 7205 32895
rect 7239 32892 7251 32895
rect 7374 32892 7380 32904
rect 7239 32864 7380 32892
rect 7239 32861 7251 32864
rect 7193 32855 7251 32861
rect 7374 32852 7380 32864
rect 7432 32892 7438 32904
rect 8202 32892 8208 32904
rect 7432 32864 8208 32892
rect 7432 32852 7438 32864
rect 8202 32852 8208 32864
rect 8260 32852 8266 32904
rect 12342 32852 12348 32904
rect 12400 32892 12406 32904
rect 12526 32892 12532 32904
rect 12400 32864 12532 32892
rect 12400 32852 12406 32864
rect 12526 32852 12532 32864
rect 12584 32852 12590 32904
rect 14090 32892 14096 32904
rect 14051 32864 14096 32892
rect 14090 32852 14096 32864
rect 14148 32852 14154 32904
rect 14274 32892 14280 32904
rect 14235 32864 14280 32892
rect 14274 32852 14280 32864
rect 14332 32852 14338 32904
rect 15746 32852 15752 32904
rect 15804 32892 15810 32904
rect 15804 32864 15849 32892
rect 15804 32852 15810 32864
rect 16206 32852 16212 32904
rect 16264 32892 16270 32904
rect 17586 32892 17592 32904
rect 16264 32864 17592 32892
rect 16264 32852 16270 32864
rect 17586 32852 17592 32864
rect 17644 32892 17650 32904
rect 17773 32895 17831 32901
rect 17773 32892 17785 32895
rect 17644 32864 17785 32892
rect 17644 32852 17650 32864
rect 17773 32861 17785 32864
rect 17819 32861 17831 32895
rect 17773 32855 17831 32861
rect 17957 32895 18015 32901
rect 17957 32861 17969 32895
rect 18003 32861 18015 32895
rect 17957 32855 18015 32861
rect 20901 32895 20959 32901
rect 20901 32861 20913 32895
rect 20947 32861 20959 32895
rect 23566 32892 23572 32904
rect 23527 32864 23572 32892
rect 20901 32855 20959 32861
rect 3191 32796 4016 32824
rect 3191 32793 3203 32796
rect 3145 32787 3203 32793
rect 1581 32759 1639 32765
rect 1581 32756 1593 32759
rect 1452 32728 1593 32756
rect 1452 32716 1458 32728
rect 1581 32725 1593 32728
rect 1627 32725 1639 32759
rect 3510 32756 3516 32768
rect 3471 32728 3516 32756
rect 1581 32719 1639 32725
rect 3510 32716 3516 32728
rect 3568 32716 3574 32768
rect 3694 32716 3700 32768
rect 3752 32756 3758 32768
rect 4080 32756 4108 32852
rect 8665 32827 8723 32833
rect 8665 32793 8677 32827
rect 8711 32824 8723 32827
rect 9582 32824 9588 32836
rect 8711 32796 9588 32824
rect 8711 32793 8723 32796
rect 8665 32787 8723 32793
rect 9582 32784 9588 32796
rect 9640 32784 9646 32836
rect 11606 32784 11612 32836
rect 11664 32824 11670 32836
rect 11885 32827 11943 32833
rect 11885 32824 11897 32827
rect 11664 32796 11897 32824
rect 11664 32784 11670 32796
rect 11885 32793 11897 32796
rect 11931 32824 11943 32827
rect 12618 32824 12624 32836
rect 11931 32796 12624 32824
rect 11931 32793 11943 32796
rect 11885 32787 11943 32793
rect 12618 32784 12624 32796
rect 12676 32784 12682 32836
rect 3752 32728 4108 32756
rect 6549 32759 6607 32765
rect 3752 32716 3758 32728
rect 6549 32725 6561 32759
rect 6595 32756 6607 32759
rect 7834 32756 7840 32768
rect 6595 32728 7840 32756
rect 6595 32725 6607 32728
rect 6549 32719 6607 32725
rect 7834 32716 7840 32728
rect 7892 32716 7898 32768
rect 9858 32756 9864 32768
rect 9819 32728 9864 32756
rect 9858 32716 9864 32728
rect 9916 32716 9922 32768
rect 11514 32716 11520 32768
rect 11572 32756 11578 32768
rect 11701 32759 11759 32765
rect 11701 32756 11713 32759
rect 11572 32728 11713 32756
rect 11572 32716 11578 32728
rect 11701 32725 11713 32728
rect 11747 32725 11759 32759
rect 11701 32719 11759 32725
rect 16758 32716 16764 32768
rect 16816 32756 16822 32768
rect 17129 32759 17187 32765
rect 17129 32756 17141 32759
rect 16816 32728 17141 32756
rect 16816 32716 16822 32728
rect 17129 32725 17141 32728
rect 17175 32725 17187 32759
rect 17972 32756 18000 32855
rect 18138 32756 18144 32768
rect 17972 32728 18144 32756
rect 17129 32719 17187 32725
rect 18138 32716 18144 32728
rect 18196 32716 18202 32768
rect 20162 32716 20168 32768
rect 20220 32756 20226 32768
rect 20625 32759 20683 32765
rect 20625 32756 20637 32759
rect 20220 32728 20637 32756
rect 20220 32716 20226 32728
rect 20625 32725 20637 32728
rect 20671 32756 20683 32759
rect 20916 32756 20944 32855
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 23676 32901 23704 32932
rect 25222 32920 25228 32932
rect 25280 32920 25286 32972
rect 23661 32895 23719 32901
rect 23661 32861 23673 32895
rect 23707 32892 23719 32895
rect 25038 32892 25044 32904
rect 23707 32864 25044 32892
rect 23707 32861 23719 32864
rect 23661 32855 23719 32861
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 25314 32892 25320 32904
rect 25275 32864 25320 32892
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 25424 32901 25452 33000
rect 27424 32997 27436 33031
rect 27470 33028 27482 33031
rect 27798 33028 27804 33040
rect 27470 33000 27804 33028
rect 27470 32997 27482 33000
rect 27424 32991 27482 32997
rect 27798 32988 27804 33000
rect 27856 33028 27862 33040
rect 28350 33028 28356 33040
rect 27856 33000 28356 33028
rect 27856 32988 27862 33000
rect 28350 32988 28356 33000
rect 28408 32988 28414 33040
rect 27154 32960 27160 32972
rect 27067 32932 27160 32960
rect 27154 32920 27160 32932
rect 27212 32960 27218 32972
rect 28626 32960 28632 32972
rect 27212 32932 28632 32960
rect 27212 32920 27218 32932
rect 28626 32920 28632 32932
rect 28684 32920 28690 32972
rect 29362 32960 29368 32972
rect 29323 32932 29368 32960
rect 29362 32920 29368 32932
rect 29420 32920 29426 32972
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32861 25467 32895
rect 25409 32855 25467 32861
rect 23109 32827 23167 32833
rect 23109 32793 23121 32827
rect 23155 32824 23167 32827
rect 23382 32824 23388 32836
rect 23155 32796 23388 32824
rect 23155 32793 23167 32796
rect 23109 32787 23167 32793
rect 23382 32784 23388 32796
rect 23440 32784 23446 32836
rect 21082 32756 21088 32768
rect 20671 32728 21088 32756
rect 20671 32725 20683 32728
rect 20625 32719 20683 32725
rect 21082 32716 21088 32728
rect 21140 32716 21146 32768
rect 24118 32756 24124 32768
rect 24079 32728 24124 32756
rect 24118 32716 24124 32728
rect 24176 32716 24182 32768
rect 28534 32756 28540 32768
rect 28495 32728 28540 32756
rect 28534 32716 28540 32728
rect 28592 32716 28598 32768
rect 29546 32756 29552 32768
rect 29507 32728 29552 32756
rect 29546 32716 29552 32728
rect 29604 32716 29610 32768
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 1765 32555 1823 32561
rect 1765 32521 1777 32555
rect 1811 32552 1823 32555
rect 1854 32552 1860 32564
rect 1811 32524 1860 32552
rect 1811 32521 1823 32524
rect 1765 32515 1823 32521
rect 1854 32512 1860 32524
rect 1912 32512 1918 32564
rect 3237 32555 3295 32561
rect 3237 32521 3249 32555
rect 3283 32552 3295 32555
rect 3326 32552 3332 32564
rect 3283 32524 3332 32552
rect 3283 32521 3295 32524
rect 3237 32515 3295 32521
rect 3326 32512 3332 32524
rect 3384 32512 3390 32564
rect 5534 32552 5540 32564
rect 5495 32524 5540 32552
rect 5534 32512 5540 32524
rect 5592 32512 5598 32564
rect 6270 32552 6276 32564
rect 6231 32524 6276 32552
rect 6270 32512 6276 32524
rect 6328 32512 6334 32564
rect 7282 32552 7288 32564
rect 6656 32524 7288 32552
rect 2958 32444 2964 32496
rect 3016 32484 3022 32496
rect 3881 32487 3939 32493
rect 3881 32484 3893 32487
rect 3016 32456 3893 32484
rect 3016 32444 3022 32456
rect 3881 32453 3893 32456
rect 3927 32453 3939 32487
rect 3881 32447 3939 32453
rect 5813 32487 5871 32493
rect 5813 32453 5825 32487
rect 5859 32484 5871 32487
rect 6656 32484 6684 32524
rect 7282 32512 7288 32524
rect 7340 32512 7346 32564
rect 7834 32552 7840 32564
rect 7795 32524 7840 32552
rect 7834 32512 7840 32524
rect 7892 32512 7898 32564
rect 11609 32555 11667 32561
rect 11609 32521 11621 32555
rect 11655 32552 11667 32555
rect 12158 32552 12164 32564
rect 11655 32524 12164 32552
rect 11655 32521 11667 32524
rect 11609 32515 11667 32521
rect 12158 32512 12164 32524
rect 12216 32512 12222 32564
rect 12526 32512 12532 32564
rect 12584 32552 12590 32564
rect 12621 32555 12679 32561
rect 12621 32552 12633 32555
rect 12584 32524 12633 32552
rect 12584 32512 12590 32524
rect 12621 32521 12633 32524
rect 12667 32521 12679 32555
rect 13262 32552 13268 32564
rect 13223 32524 13268 32552
rect 12621 32515 12679 32521
rect 13262 32512 13268 32524
rect 13320 32512 13326 32564
rect 14182 32552 14188 32564
rect 14143 32524 14188 32552
rect 14182 32512 14188 32524
rect 14240 32512 14246 32564
rect 14369 32555 14427 32561
rect 14369 32521 14381 32555
rect 14415 32552 14427 32555
rect 15102 32552 15108 32564
rect 14415 32524 15108 32552
rect 14415 32521 14427 32524
rect 14369 32515 14427 32521
rect 15102 32512 15108 32524
rect 15160 32512 15166 32564
rect 15473 32555 15531 32561
rect 15473 32521 15485 32555
rect 15519 32552 15531 32555
rect 15562 32552 15568 32564
rect 15519 32524 15568 32552
rect 15519 32521 15531 32524
rect 15473 32515 15531 32521
rect 15562 32512 15568 32524
rect 15620 32512 15626 32564
rect 16206 32552 16212 32564
rect 16167 32524 16212 32552
rect 16206 32512 16212 32524
rect 16264 32512 16270 32564
rect 20162 32552 20168 32564
rect 20123 32524 20168 32552
rect 20162 32512 20168 32524
rect 20220 32512 20226 32564
rect 20622 32552 20628 32564
rect 20583 32524 20628 32552
rect 20622 32512 20628 32524
rect 20680 32552 20686 32564
rect 22465 32555 22523 32561
rect 22465 32552 22477 32555
rect 20680 32524 22477 32552
rect 20680 32512 20686 32524
rect 22465 32521 22477 32524
rect 22511 32552 22523 32555
rect 23201 32555 23259 32561
rect 23201 32552 23213 32555
rect 22511 32524 23213 32552
rect 22511 32521 22523 32524
rect 22465 32515 22523 32521
rect 23201 32521 23213 32524
rect 23247 32552 23259 32555
rect 23566 32552 23572 32564
rect 23247 32524 23572 32552
rect 23247 32521 23259 32524
rect 23201 32515 23259 32521
rect 23566 32512 23572 32524
rect 23624 32512 23630 32564
rect 25222 32552 25228 32564
rect 25183 32524 25228 32552
rect 25222 32512 25228 32524
rect 25280 32512 25286 32564
rect 25314 32512 25320 32564
rect 25372 32552 25378 32564
rect 26237 32555 26295 32561
rect 26237 32552 26249 32555
rect 25372 32524 26249 32552
rect 25372 32512 25378 32524
rect 26237 32521 26249 32524
rect 26283 32552 26295 32555
rect 26789 32555 26847 32561
rect 26789 32552 26801 32555
rect 26283 32524 26801 32552
rect 26283 32521 26295 32524
rect 26237 32515 26295 32521
rect 26789 32521 26801 32524
rect 26835 32521 26847 32555
rect 27798 32552 27804 32564
rect 27759 32524 27804 32552
rect 26789 32515 26847 32521
rect 27798 32512 27804 32524
rect 27856 32512 27862 32564
rect 28626 32552 28632 32564
rect 28587 32524 28632 32552
rect 28626 32512 28632 32524
rect 28684 32512 28690 32564
rect 29362 32512 29368 32564
rect 29420 32552 29426 32564
rect 29457 32555 29515 32561
rect 29457 32552 29469 32555
rect 29420 32524 29469 32552
rect 29420 32512 29426 32524
rect 29457 32521 29469 32524
rect 29503 32521 29515 32555
rect 29457 32515 29515 32521
rect 5859 32456 6684 32484
rect 6825 32487 6883 32493
rect 5859 32453 5871 32456
rect 5813 32447 5871 32453
rect 6825 32453 6837 32487
rect 6871 32484 6883 32487
rect 8297 32487 8355 32493
rect 8297 32484 8309 32487
rect 6871 32456 8309 32484
rect 6871 32453 6883 32456
rect 6825 32447 6883 32453
rect 8297 32453 8309 32456
rect 8343 32484 8355 32487
rect 8478 32484 8484 32496
rect 8343 32456 8484 32484
rect 8343 32453 8355 32456
rect 8297 32447 8355 32453
rect 8478 32444 8484 32456
rect 8536 32444 8542 32496
rect 11977 32487 12035 32493
rect 11977 32453 11989 32487
rect 12023 32484 12035 32487
rect 12250 32484 12256 32496
rect 12023 32456 12256 32484
rect 12023 32453 12035 32456
rect 11977 32447 12035 32453
rect 12250 32444 12256 32456
rect 12308 32444 12314 32496
rect 13280 32484 13308 32512
rect 15746 32484 15752 32496
rect 13280 32456 15752 32484
rect 15746 32444 15752 32456
rect 15804 32444 15810 32496
rect 22094 32444 22100 32496
rect 22152 32484 22158 32496
rect 22741 32487 22799 32493
rect 22741 32484 22753 32487
rect 22152 32456 22753 32484
rect 22152 32444 22158 32456
rect 22741 32453 22753 32456
rect 22787 32453 22799 32487
rect 28169 32487 28227 32493
rect 28169 32484 28181 32487
rect 22741 32447 22799 32453
rect 25884 32456 28181 32484
rect 25884 32428 25912 32456
rect 3510 32376 3516 32428
rect 3568 32416 3574 32428
rect 3970 32416 3976 32428
rect 3568 32388 3976 32416
rect 3568 32376 3574 32388
rect 3970 32376 3976 32388
rect 4028 32416 4034 32428
rect 4617 32419 4675 32425
rect 4617 32416 4629 32419
rect 4028 32388 4629 32416
rect 4028 32376 4034 32388
rect 4617 32385 4629 32388
rect 4663 32416 4675 32419
rect 5166 32416 5172 32428
rect 4663 32388 5172 32416
rect 4663 32385 4675 32388
rect 4617 32379 4675 32385
rect 5166 32376 5172 32388
rect 5224 32376 5230 32428
rect 7374 32416 7380 32428
rect 7335 32388 7380 32416
rect 7374 32376 7380 32388
rect 7432 32376 7438 32428
rect 8662 32376 8668 32428
rect 8720 32416 8726 32428
rect 8941 32419 8999 32425
rect 8941 32416 8953 32419
rect 8720 32388 8953 32416
rect 8720 32376 8726 32388
rect 8941 32385 8953 32388
rect 8987 32385 8999 32419
rect 8941 32379 8999 32385
rect 13725 32419 13783 32425
rect 13725 32385 13737 32419
rect 13771 32416 13783 32419
rect 14090 32416 14096 32428
rect 13771 32388 14096 32416
rect 13771 32385 13783 32388
rect 13725 32379 13783 32385
rect 14090 32376 14096 32388
rect 14148 32376 14154 32428
rect 14918 32416 14924 32428
rect 14879 32388 14924 32416
rect 14918 32376 14924 32388
rect 14976 32376 14982 32428
rect 16945 32419 17003 32425
rect 16945 32385 16957 32419
rect 16991 32416 17003 32419
rect 17678 32416 17684 32428
rect 16991 32388 17684 32416
rect 16991 32385 17003 32388
rect 16945 32379 17003 32385
rect 17678 32376 17684 32388
rect 17736 32376 17742 32428
rect 21082 32416 21088 32428
rect 21043 32388 21088 32416
rect 21082 32376 21088 32388
rect 21140 32376 21146 32428
rect 24210 32416 24216 32428
rect 24171 32388 24216 32416
rect 24210 32376 24216 32388
rect 24268 32376 24274 32428
rect 25038 32376 25044 32428
rect 25096 32416 25102 32428
rect 25777 32419 25835 32425
rect 25777 32416 25789 32419
rect 25096 32388 25789 32416
rect 25096 32376 25102 32388
rect 25777 32385 25789 32388
rect 25823 32416 25835 32419
rect 25866 32416 25872 32428
rect 25823 32388 25872 32416
rect 25823 32385 25835 32388
rect 25777 32379 25835 32385
rect 25866 32376 25872 32388
rect 25924 32376 25930 32428
rect 26697 32419 26755 32425
rect 26697 32385 26709 32419
rect 26743 32416 26755 32419
rect 27062 32416 27068 32428
rect 26743 32388 27068 32416
rect 26743 32385 26755 32388
rect 26697 32379 26755 32385
rect 27062 32376 27068 32388
rect 27120 32416 27126 32428
rect 27356 32425 27384 32456
rect 28169 32453 28181 32456
rect 28215 32453 28227 32487
rect 28169 32447 28227 32453
rect 27249 32419 27307 32425
rect 27249 32416 27261 32419
rect 27120 32388 27261 32416
rect 27120 32376 27126 32388
rect 27249 32385 27261 32388
rect 27295 32385 27307 32419
rect 27249 32379 27307 32385
rect 27341 32419 27399 32425
rect 27341 32385 27353 32419
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 1394 32308 1400 32360
rect 1452 32348 1458 32360
rect 1857 32351 1915 32357
rect 1857 32348 1869 32351
rect 1452 32320 1869 32348
rect 1452 32308 1458 32320
rect 1857 32317 1869 32320
rect 1903 32348 1915 32351
rect 3234 32348 3240 32360
rect 1903 32320 3240 32348
rect 1903 32317 1915 32320
rect 1857 32311 1915 32317
rect 3234 32308 3240 32320
rect 3292 32348 3298 32360
rect 3694 32348 3700 32360
rect 3292 32320 3700 32348
rect 3292 32308 3298 32320
rect 3694 32308 3700 32320
rect 3752 32308 3758 32360
rect 3786 32308 3792 32360
rect 3844 32348 3850 32360
rect 4433 32351 4491 32357
rect 4433 32348 4445 32351
rect 3844 32320 4445 32348
rect 3844 32308 3850 32320
rect 4433 32317 4445 32320
rect 4479 32317 4491 32351
rect 4433 32311 4491 32317
rect 5534 32308 5540 32360
rect 5592 32348 5598 32360
rect 5629 32351 5687 32357
rect 5629 32348 5641 32351
rect 5592 32320 5641 32348
rect 5592 32308 5598 32320
rect 5629 32317 5641 32320
rect 5675 32317 5687 32351
rect 5629 32311 5687 32317
rect 7834 32308 7840 32360
rect 7892 32348 7898 32360
rect 8757 32351 8815 32357
rect 8757 32348 8769 32351
rect 7892 32320 8769 32348
rect 7892 32308 7898 32320
rect 8757 32317 8769 32320
rect 8803 32348 8815 32351
rect 9674 32348 9680 32360
rect 8803 32320 9680 32348
rect 8803 32317 8815 32320
rect 8757 32311 8815 32317
rect 9674 32308 9680 32320
rect 9732 32308 9738 32360
rect 14182 32308 14188 32360
rect 14240 32348 14246 32360
rect 14737 32351 14795 32357
rect 14737 32348 14749 32351
rect 14240 32320 14749 32348
rect 14240 32308 14246 32320
rect 14737 32317 14749 32320
rect 14783 32317 14795 32351
rect 14737 32311 14795 32317
rect 14829 32351 14887 32357
rect 14829 32317 14841 32351
rect 14875 32348 14887 32351
rect 15102 32348 15108 32360
rect 14875 32320 15108 32348
rect 14875 32317 14887 32320
rect 14829 32311 14887 32317
rect 15102 32308 15108 32320
rect 15160 32308 15166 32360
rect 16393 32351 16451 32357
rect 16393 32317 16405 32351
rect 16439 32348 16451 32351
rect 16574 32348 16580 32360
rect 16439 32320 16580 32348
rect 16439 32317 16451 32320
rect 16393 32311 16451 32317
rect 16574 32308 16580 32320
rect 16632 32348 16638 32360
rect 16669 32351 16727 32357
rect 16669 32348 16681 32351
rect 16632 32320 16681 32348
rect 16632 32308 16638 32320
rect 16669 32317 16681 32320
rect 16715 32317 16727 32351
rect 16669 32311 16727 32317
rect 18049 32351 18107 32357
rect 18049 32317 18061 32351
rect 18095 32348 18107 32351
rect 18138 32348 18144 32360
rect 18095 32320 18144 32348
rect 18095 32317 18107 32320
rect 18049 32311 18107 32317
rect 18138 32308 18144 32320
rect 18196 32348 18202 32360
rect 18874 32348 18880 32360
rect 18196 32320 18880 32348
rect 18196 32308 18202 32320
rect 18874 32308 18880 32320
rect 18932 32348 18938 32360
rect 19797 32351 19855 32357
rect 19797 32348 19809 32351
rect 18932 32320 19809 32348
rect 18932 32308 18938 32320
rect 19797 32317 19809 32320
rect 19843 32348 19855 32351
rect 19978 32348 19984 32360
rect 19843 32320 19984 32348
rect 19843 32317 19855 32320
rect 19797 32311 19855 32317
rect 19978 32308 19984 32320
rect 20036 32348 20042 32360
rect 20898 32348 20904 32360
rect 20036 32320 20904 32348
rect 20036 32308 20042 32320
rect 20898 32308 20904 32320
rect 20956 32308 20962 32360
rect 23290 32308 23296 32360
rect 23348 32348 23354 32360
rect 24029 32351 24087 32357
rect 24029 32348 24041 32351
rect 23348 32320 24041 32348
rect 23348 32308 23354 32320
rect 24029 32317 24041 32320
rect 24075 32348 24087 32351
rect 24118 32348 24124 32360
rect 24075 32320 24124 32348
rect 24075 32317 24087 32320
rect 24029 32311 24087 32317
rect 24118 32308 24124 32320
rect 24176 32308 24182 32360
rect 26878 32308 26884 32360
rect 26936 32348 26942 32360
rect 27157 32351 27215 32357
rect 27157 32348 27169 32351
rect 26936 32320 27169 32348
rect 26936 32308 26942 32320
rect 27157 32317 27169 32320
rect 27203 32348 27215 32351
rect 27798 32348 27804 32360
rect 27203 32320 27804 32348
rect 27203 32317 27215 32320
rect 27157 32311 27215 32317
rect 27798 32308 27804 32320
rect 27856 32308 27862 32360
rect 2124 32283 2182 32289
rect 2124 32249 2136 32283
rect 2170 32280 2182 32283
rect 2774 32280 2780 32292
rect 2170 32252 2780 32280
rect 2170 32249 2182 32252
rect 2124 32243 2182 32249
rect 2774 32240 2780 32252
rect 2832 32240 2838 32292
rect 7285 32283 7343 32289
rect 7285 32280 7297 32283
rect 6564 32252 7297 32280
rect 3605 32215 3663 32221
rect 3605 32181 3617 32215
rect 3651 32212 3663 32215
rect 3694 32212 3700 32224
rect 3651 32184 3700 32212
rect 3651 32181 3663 32184
rect 3605 32175 3663 32181
rect 3694 32172 3700 32184
rect 3752 32172 3758 32224
rect 4062 32212 4068 32224
rect 4023 32184 4068 32212
rect 4062 32172 4068 32184
rect 4120 32172 4126 32224
rect 4522 32172 4528 32224
rect 4580 32212 4586 32224
rect 5077 32215 5135 32221
rect 5077 32212 5089 32215
rect 4580 32184 5089 32212
rect 4580 32172 4586 32184
rect 5077 32181 5089 32184
rect 5123 32181 5135 32215
rect 5077 32175 5135 32181
rect 5534 32172 5540 32224
rect 5592 32212 5598 32224
rect 6564 32221 6592 32252
rect 7285 32249 7297 32252
rect 7331 32249 7343 32283
rect 7285 32243 7343 32249
rect 8478 32240 8484 32292
rect 8536 32280 8542 32292
rect 8849 32283 8907 32289
rect 8849 32280 8861 32283
rect 8536 32252 8861 32280
rect 8536 32240 8542 32252
rect 8849 32249 8861 32252
rect 8895 32249 8907 32283
rect 8849 32243 8907 32249
rect 17497 32283 17555 32289
rect 17497 32249 17509 32283
rect 17543 32280 17555 32283
rect 18294 32283 18352 32289
rect 18294 32280 18306 32283
rect 17543 32252 18306 32280
rect 17543 32249 17555 32252
rect 17497 32243 17555 32249
rect 18294 32249 18306 32252
rect 18340 32280 18352 32283
rect 19150 32280 19156 32292
rect 18340 32252 19156 32280
rect 18340 32249 18352 32252
rect 18294 32243 18352 32249
rect 19150 32240 19156 32252
rect 19208 32240 19214 32292
rect 21330 32283 21388 32289
rect 21330 32280 21342 32283
rect 20916 32252 21342 32280
rect 6549 32215 6607 32221
rect 6549 32212 6561 32215
rect 5592 32184 6561 32212
rect 5592 32172 5598 32184
rect 6549 32181 6561 32184
rect 6595 32181 6607 32215
rect 7190 32212 7196 32224
rect 7151 32184 7196 32212
rect 6549 32175 6607 32181
rect 7190 32172 7196 32184
rect 7248 32172 7254 32224
rect 8386 32212 8392 32224
rect 8347 32184 8392 32212
rect 8386 32172 8392 32184
rect 8444 32172 8450 32224
rect 17865 32215 17923 32221
rect 17865 32181 17877 32215
rect 17911 32212 17923 32215
rect 18138 32212 18144 32224
rect 17911 32184 18144 32212
rect 17911 32181 17923 32184
rect 17865 32175 17923 32181
rect 18138 32172 18144 32184
rect 18196 32172 18202 32224
rect 19426 32212 19432 32224
rect 19387 32184 19432 32212
rect 19426 32172 19432 32184
rect 19484 32172 19490 32224
rect 20806 32172 20812 32224
rect 20864 32212 20870 32224
rect 20916 32221 20944 32252
rect 21330 32249 21342 32252
rect 21376 32249 21388 32283
rect 21330 32243 21388 32249
rect 24765 32283 24823 32289
rect 24765 32249 24777 32283
rect 24811 32280 24823 32283
rect 25593 32283 25651 32289
rect 25593 32280 25605 32283
rect 24811 32252 25605 32280
rect 24811 32249 24823 32252
rect 24765 32243 24823 32249
rect 25593 32249 25605 32252
rect 25639 32280 25651 32283
rect 26234 32280 26240 32292
rect 25639 32252 26240 32280
rect 25639 32249 25651 32252
rect 25593 32243 25651 32249
rect 26234 32240 26240 32252
rect 26292 32240 26298 32292
rect 20901 32215 20959 32221
rect 20901 32212 20913 32215
rect 20864 32184 20913 32212
rect 20864 32172 20870 32184
rect 20901 32181 20913 32184
rect 20947 32181 20959 32215
rect 23658 32212 23664 32224
rect 23619 32184 23664 32212
rect 20901 32175 20959 32181
rect 23658 32172 23664 32184
rect 23716 32172 23722 32224
rect 24118 32212 24124 32224
rect 24079 32184 24124 32212
rect 24118 32172 24124 32184
rect 24176 32172 24182 32224
rect 25133 32215 25191 32221
rect 25133 32181 25145 32215
rect 25179 32212 25191 32215
rect 25685 32215 25743 32221
rect 25685 32212 25697 32215
rect 25179 32184 25697 32212
rect 25179 32181 25191 32184
rect 25133 32175 25191 32181
rect 25685 32181 25697 32184
rect 25731 32212 25743 32215
rect 26694 32212 26700 32224
rect 25731 32184 26700 32212
rect 25731 32181 25743 32184
rect 25685 32175 25743 32181
rect 26694 32172 26700 32184
rect 26752 32172 26758 32224
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 2774 31968 2780 32020
rect 2832 32008 2838 32020
rect 3234 32008 3240 32020
rect 2832 31980 2925 32008
rect 3195 31980 3240 32008
rect 2832 31968 2838 31980
rect 3234 31968 3240 31980
rect 3292 31968 3298 32020
rect 4065 32011 4123 32017
rect 4065 31977 4077 32011
rect 4111 32008 4123 32011
rect 4522 32008 4528 32020
rect 4111 31980 4528 32008
rect 4111 31977 4123 31980
rect 4065 31971 4123 31977
rect 4522 31968 4528 31980
rect 4580 31968 4586 32020
rect 5166 32008 5172 32020
rect 5127 31980 5172 32008
rect 5166 31968 5172 31980
rect 5224 31968 5230 32020
rect 5813 32011 5871 32017
rect 5813 31977 5825 32011
rect 5859 32008 5871 32011
rect 6270 32008 6276 32020
rect 5859 31980 6276 32008
rect 5859 31977 5871 31980
rect 5813 31971 5871 31977
rect 6270 31968 6276 31980
rect 6328 31968 6334 32020
rect 6917 32011 6975 32017
rect 6917 31977 6929 32011
rect 6963 32008 6975 32011
rect 7190 32008 7196 32020
rect 6963 31980 7196 32008
rect 6963 31977 6975 31980
rect 6917 31971 6975 31977
rect 7190 31968 7196 31980
rect 7248 31968 7254 32020
rect 7282 31968 7288 32020
rect 7340 32008 7346 32020
rect 7340 31980 7385 32008
rect 7340 31968 7346 31980
rect 8386 31968 8392 32020
rect 8444 32008 8450 32020
rect 9033 32011 9091 32017
rect 9033 32008 9045 32011
rect 8444 31980 9045 32008
rect 8444 31968 8450 31980
rect 9033 31977 9045 31980
rect 9079 31977 9091 32011
rect 9033 31971 9091 31977
rect 13725 32011 13783 32017
rect 13725 31977 13737 32011
rect 13771 32008 13783 32011
rect 14274 32008 14280 32020
rect 13771 31980 14280 32008
rect 13771 31977 13783 31980
rect 13725 31971 13783 31977
rect 14274 31968 14280 31980
rect 14332 31968 14338 32020
rect 14829 32011 14887 32017
rect 14829 31977 14841 32011
rect 14875 32008 14887 32011
rect 15102 32008 15108 32020
rect 14875 31980 15108 32008
rect 14875 31977 14887 31980
rect 14829 31971 14887 31977
rect 15102 31968 15108 31980
rect 15160 31968 15166 32020
rect 15562 31968 15568 32020
rect 15620 32008 15626 32020
rect 16117 32011 16175 32017
rect 16117 32008 16129 32011
rect 15620 31980 16129 32008
rect 15620 31968 15626 31980
rect 16117 31977 16129 31980
rect 16163 31977 16175 32011
rect 16117 31971 16175 31977
rect 17773 32011 17831 32017
rect 17773 31977 17785 32011
rect 17819 32008 17831 32011
rect 17862 32008 17868 32020
rect 17819 31980 17868 32008
rect 17819 31977 17831 31980
rect 17773 31971 17831 31977
rect 17862 31968 17868 31980
rect 17920 31968 17926 32020
rect 18874 32008 18880 32020
rect 18835 31980 18880 32008
rect 18874 31968 18880 31980
rect 18932 31968 18938 32020
rect 20806 31968 20812 32020
rect 20864 32008 20870 32020
rect 22465 32011 22523 32017
rect 22465 32008 22477 32011
rect 20864 31980 22477 32008
rect 20864 31968 20870 31980
rect 22465 31977 22477 31980
rect 22511 31977 22523 32011
rect 22465 31971 22523 31977
rect 22922 31968 22928 32020
rect 22980 32008 22986 32020
rect 23109 32011 23167 32017
rect 23109 32008 23121 32011
rect 22980 31980 23121 32008
rect 22980 31968 22986 31980
rect 23109 31977 23121 31980
rect 23155 31977 23167 32011
rect 23109 31971 23167 31977
rect 23477 32011 23535 32017
rect 23477 31977 23489 32011
rect 23523 32008 23535 32011
rect 23937 32011 23995 32017
rect 23937 32008 23949 32011
rect 23523 31980 23949 32008
rect 23523 31977 23535 31980
rect 23477 31971 23535 31977
rect 23937 31977 23949 31980
rect 23983 32008 23995 32011
rect 24118 32008 24124 32020
rect 23983 31980 24124 32008
rect 23983 31977 23995 31980
rect 23937 31971 23995 31977
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 24210 31968 24216 32020
rect 24268 32008 24274 32020
rect 24765 32011 24823 32017
rect 24268 31980 24313 32008
rect 24268 31968 24274 31980
rect 24765 31977 24777 32011
rect 24811 32008 24823 32011
rect 25222 32008 25228 32020
rect 24811 31980 25228 32008
rect 24811 31977 24823 31980
rect 24765 31971 24823 31977
rect 25222 31968 25228 31980
rect 25280 31968 25286 32020
rect 25866 32008 25872 32020
rect 25827 31980 25872 32008
rect 25866 31968 25872 31980
rect 25924 31968 25930 32020
rect 26878 32008 26884 32020
rect 26839 31980 26884 32008
rect 26878 31968 26884 31980
rect 26936 31968 26942 32020
rect 35621 32011 35679 32017
rect 35621 31977 35633 32011
rect 35667 32008 35679 32011
rect 35802 32008 35808 32020
rect 35667 31980 35808 32008
rect 35667 31977 35679 31980
rect 35621 31971 35679 31977
rect 35802 31968 35808 31980
rect 35860 31968 35866 32020
rect 2792 31940 2820 31968
rect 3418 31940 3424 31952
rect 2792 31912 3424 31940
rect 3418 31900 3424 31912
rect 3476 31940 3482 31952
rect 3694 31940 3700 31952
rect 3476 31912 3700 31940
rect 3476 31900 3482 31912
rect 3694 31900 3700 31912
rect 3752 31940 3758 31952
rect 4433 31943 4491 31949
rect 4433 31940 4445 31943
rect 3752 31912 4445 31940
rect 3752 31900 3758 31912
rect 4433 31909 4445 31912
rect 4479 31909 4491 31943
rect 4433 31903 4491 31909
rect 6549 31943 6607 31949
rect 6549 31909 6561 31943
rect 6595 31940 6607 31943
rect 7374 31940 7380 31952
rect 6595 31912 7380 31940
rect 6595 31909 6607 31912
rect 6549 31903 6607 31909
rect 7374 31900 7380 31912
rect 7432 31940 7438 31952
rect 7561 31943 7619 31949
rect 7561 31940 7573 31943
rect 7432 31912 7573 31940
rect 7432 31900 7438 31912
rect 7561 31909 7573 31912
rect 7607 31909 7619 31943
rect 7561 31903 7619 31909
rect 11054 31900 11060 31952
rect 11112 31940 11118 31952
rect 11232 31943 11290 31949
rect 11232 31940 11244 31943
rect 11112 31912 11244 31940
rect 11112 31900 11118 31912
rect 11232 31909 11244 31912
rect 11278 31940 11290 31943
rect 14461 31943 14519 31949
rect 14461 31940 14473 31943
rect 11278 31912 14473 31940
rect 11278 31909 11290 31912
rect 11232 31903 11290 31909
rect 14461 31909 14473 31912
rect 14507 31940 14519 31943
rect 14918 31940 14924 31952
rect 14507 31912 14924 31940
rect 14507 31909 14519 31912
rect 14461 31903 14519 31909
rect 14918 31900 14924 31912
rect 14976 31900 14982 31952
rect 15841 31943 15899 31949
rect 15841 31909 15853 31943
rect 15887 31940 15899 31943
rect 16022 31940 16028 31952
rect 15887 31912 16028 31940
rect 15887 31909 15899 31912
rect 15841 31903 15899 31909
rect 16022 31900 16028 31912
rect 16080 31900 16086 31952
rect 20717 31943 20775 31949
rect 20717 31909 20729 31943
rect 20763 31940 20775 31943
rect 21082 31940 21088 31952
rect 20763 31912 21088 31940
rect 20763 31909 20775 31912
rect 20717 31903 20775 31909
rect 21082 31900 21088 31912
rect 21140 31900 21146 31952
rect 22002 31900 22008 31952
rect 22060 31940 22066 31952
rect 22940 31940 22968 31968
rect 22060 31912 22968 31940
rect 22060 31900 22066 31912
rect 25130 31900 25136 31952
rect 25188 31940 25194 31952
rect 25317 31943 25375 31949
rect 25317 31940 25329 31943
rect 25188 31912 25329 31940
rect 25188 31900 25194 31912
rect 25317 31909 25329 31912
rect 25363 31909 25375 31943
rect 25317 31903 25375 31909
rect 26694 31900 26700 31952
rect 26752 31940 26758 31952
rect 27332 31943 27390 31949
rect 27332 31940 27344 31943
rect 26752 31912 27344 31940
rect 26752 31900 26758 31912
rect 27332 31909 27344 31912
rect 27378 31940 27390 31943
rect 28534 31940 28540 31952
rect 27378 31912 28540 31940
rect 27378 31909 27390 31912
rect 27332 31903 27390 31909
rect 28534 31900 28540 31912
rect 28592 31900 28598 31952
rect 1664 31875 1722 31881
rect 1664 31841 1676 31875
rect 1710 31872 1722 31875
rect 2498 31872 2504 31884
rect 1710 31844 2504 31872
rect 1710 31841 1722 31844
rect 1664 31835 1722 31841
rect 2498 31832 2504 31844
rect 2556 31832 2562 31884
rect 4525 31875 4583 31881
rect 4525 31841 4537 31875
rect 4571 31872 4583 31875
rect 4706 31872 4712 31884
rect 4571 31844 4712 31872
rect 4571 31841 4583 31844
rect 4525 31835 4583 31841
rect 4706 31832 4712 31844
rect 4764 31832 4770 31884
rect 5626 31872 5632 31884
rect 5587 31844 5632 31872
rect 5626 31832 5632 31844
rect 5684 31832 5690 31884
rect 8478 31872 8484 31884
rect 8439 31844 8484 31872
rect 8478 31832 8484 31844
rect 8536 31832 8542 31884
rect 9398 31832 9404 31884
rect 9456 31872 9462 31884
rect 10965 31875 11023 31881
rect 10965 31872 10977 31875
rect 9456 31844 10977 31872
rect 9456 31832 9462 31844
rect 10965 31841 10977 31844
rect 11011 31872 11023 31875
rect 11514 31872 11520 31884
rect 11011 31844 11520 31872
rect 11011 31841 11023 31844
rect 10965 31835 11023 31841
rect 11514 31832 11520 31844
rect 11572 31832 11578 31884
rect 18138 31872 18144 31884
rect 18099 31844 18144 31872
rect 18138 31832 18144 31844
rect 18196 31832 18202 31884
rect 18414 31872 18420 31884
rect 18248 31844 18420 31872
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 4617 31807 4675 31813
rect 4617 31773 4629 31807
rect 4663 31773 4675 31807
rect 4617 31767 4675 31773
rect 4632 31736 4660 31767
rect 5166 31764 5172 31816
rect 5224 31804 5230 31816
rect 9306 31804 9312 31816
rect 5224 31776 5488 31804
rect 5224 31764 5230 31776
rect 4890 31736 4896 31748
rect 4632 31708 4896 31736
rect 4890 31696 4896 31708
rect 4948 31696 4954 31748
rect 5460 31736 5488 31776
rect 8680 31776 9312 31804
rect 8680 31745 8708 31776
rect 9306 31764 9312 31776
rect 9364 31764 9370 31816
rect 9493 31807 9551 31813
rect 9493 31773 9505 31807
rect 9539 31804 9551 31807
rect 9582 31804 9588 31816
rect 9539 31776 9588 31804
rect 9539 31773 9551 31776
rect 9493 31767 9551 31773
rect 9582 31764 9588 31776
rect 9640 31764 9646 31816
rect 15286 31804 15292 31816
rect 15247 31776 15292 31804
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 18248 31813 18276 31844
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 21352 31875 21410 31881
rect 21352 31841 21364 31875
rect 21398 31872 21410 31875
rect 21634 31872 21640 31884
rect 21398 31844 21640 31872
rect 21398 31841 21410 31844
rect 21352 31835 21410 31841
rect 21634 31832 21640 31844
rect 21692 31832 21698 31884
rect 23293 31875 23351 31881
rect 23293 31841 23305 31875
rect 23339 31872 23351 31875
rect 23382 31872 23388 31884
rect 23339 31844 23388 31872
rect 23339 31841 23351 31844
rect 23293 31835 23351 31841
rect 23382 31832 23388 31844
rect 23440 31832 23446 31884
rect 24762 31832 24768 31884
rect 24820 31872 24826 31884
rect 25222 31872 25228 31884
rect 24820 31844 25228 31872
rect 24820 31832 24826 31844
rect 25222 31832 25228 31844
rect 25280 31832 25286 31884
rect 25332 31844 25544 31872
rect 18233 31807 18291 31813
rect 18233 31804 18245 31807
rect 17972 31776 18245 31804
rect 8665 31739 8723 31745
rect 5460 31708 5580 31736
rect 3694 31668 3700 31680
rect 3655 31640 3700 31668
rect 3694 31628 3700 31640
rect 3752 31628 3758 31680
rect 5552 31668 5580 31708
rect 8665 31705 8677 31739
rect 8711 31736 8723 31739
rect 8711 31708 8745 31736
rect 8711 31705 8723 31708
rect 8665 31699 8723 31705
rect 17862 31696 17868 31748
rect 17920 31736 17926 31748
rect 17972 31736 18000 31776
rect 18233 31773 18245 31776
rect 18279 31773 18291 31807
rect 18233 31767 18291 31773
rect 18325 31807 18383 31813
rect 18325 31773 18337 31807
rect 18371 31804 18383 31807
rect 18371 31776 18405 31804
rect 18371 31773 18383 31776
rect 18325 31767 18383 31773
rect 17920 31708 18000 31736
rect 17920 31696 17926 31708
rect 18046 31696 18052 31748
rect 18104 31736 18110 31748
rect 18340 31736 18368 31767
rect 20898 31764 20904 31816
rect 20956 31804 20962 31816
rect 21085 31807 21143 31813
rect 21085 31804 21097 31807
rect 20956 31776 21097 31804
rect 20956 31764 20962 31776
rect 21085 31773 21097 31776
rect 21131 31773 21143 31807
rect 21085 31767 21143 31773
rect 24210 31764 24216 31816
rect 24268 31804 24274 31816
rect 25332 31804 25360 31844
rect 25516 31816 25544 31844
rect 26786 31832 26792 31884
rect 26844 31872 26850 31884
rect 27065 31875 27123 31881
rect 27065 31872 27077 31875
rect 26844 31844 27077 31872
rect 26844 31832 26850 31844
rect 27065 31841 27077 31844
rect 27111 31872 27123 31875
rect 27154 31872 27160 31884
rect 27111 31844 27160 31872
rect 27111 31841 27123 31844
rect 27065 31835 27123 31841
rect 27154 31832 27160 31844
rect 27212 31832 27218 31884
rect 35434 31872 35440 31884
rect 35395 31844 35440 31872
rect 35434 31832 35440 31844
rect 35492 31832 35498 31884
rect 24268 31776 25360 31804
rect 24268 31764 24274 31776
rect 25498 31764 25504 31816
rect 25556 31804 25562 31816
rect 25556 31776 25649 31804
rect 25556 31764 25562 31776
rect 18598 31736 18604 31748
rect 18104 31708 18604 31736
rect 18104 31696 18110 31708
rect 18598 31696 18604 31708
rect 18656 31696 18662 31748
rect 5718 31668 5724 31680
rect 5552 31640 5724 31668
rect 5718 31628 5724 31640
rect 5776 31668 5782 31680
rect 5902 31668 5908 31680
rect 5776 31640 5908 31668
rect 5776 31628 5782 31640
rect 5902 31628 5908 31640
rect 5960 31628 5966 31680
rect 12342 31668 12348 31680
rect 12303 31640 12348 31668
rect 12342 31628 12348 31640
rect 12400 31628 12406 31680
rect 24854 31668 24860 31680
rect 24815 31640 24860 31668
rect 24854 31628 24860 31640
rect 24912 31628 24918 31680
rect 28442 31668 28448 31680
rect 28403 31640 28448 31668
rect 28442 31628 28448 31640
rect 28500 31628 28506 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 3418 31464 3424 31476
rect 3379 31436 3424 31464
rect 3418 31424 3424 31436
rect 3476 31424 3482 31476
rect 4706 31464 4712 31476
rect 4667 31436 4712 31464
rect 4706 31424 4712 31436
rect 4764 31424 4770 31476
rect 5626 31424 5632 31476
rect 5684 31464 5690 31476
rect 6181 31467 6239 31473
rect 6181 31464 6193 31467
rect 5684 31436 6193 31464
rect 5684 31424 5690 31436
rect 6181 31433 6193 31436
rect 6227 31433 6239 31467
rect 6181 31427 6239 31433
rect 7009 31467 7067 31473
rect 7009 31433 7021 31467
rect 7055 31464 7067 31467
rect 7190 31464 7196 31476
rect 7055 31436 7196 31464
rect 7055 31433 7067 31436
rect 7009 31427 7067 31433
rect 7190 31424 7196 31436
rect 7248 31424 7254 31476
rect 8478 31464 8484 31476
rect 8439 31436 8484 31464
rect 8478 31424 8484 31436
rect 8536 31424 8542 31476
rect 8570 31424 8576 31476
rect 8628 31464 8634 31476
rect 8757 31467 8815 31473
rect 8757 31464 8769 31467
rect 8628 31436 8769 31464
rect 8628 31424 8634 31436
rect 8757 31433 8769 31436
rect 8803 31464 8815 31467
rect 9398 31464 9404 31476
rect 8803 31436 9404 31464
rect 8803 31433 8815 31436
rect 8757 31427 8815 31433
rect 9398 31424 9404 31436
rect 9456 31424 9462 31476
rect 10873 31467 10931 31473
rect 10873 31433 10885 31467
rect 10919 31464 10931 31467
rect 10962 31464 10968 31476
rect 10919 31436 10968 31464
rect 10919 31433 10931 31436
rect 10873 31427 10931 31433
rect 10962 31424 10968 31436
rect 11020 31424 11026 31476
rect 11882 31464 11888 31476
rect 11843 31436 11888 31464
rect 11882 31424 11888 31436
rect 11940 31424 11946 31476
rect 12621 31467 12679 31473
rect 12621 31433 12633 31467
rect 12667 31464 12679 31467
rect 13081 31467 13139 31473
rect 12667 31436 12756 31464
rect 12667 31433 12679 31436
rect 12621 31427 12679 31433
rect 2498 31356 2504 31408
rect 2556 31396 2562 31408
rect 2777 31399 2835 31405
rect 2777 31396 2789 31399
rect 2556 31368 2789 31396
rect 2556 31356 2562 31368
rect 2777 31365 2789 31368
rect 2823 31396 2835 31399
rect 4724 31396 4752 31424
rect 2823 31368 4752 31396
rect 2823 31365 2835 31368
rect 2777 31359 2835 31365
rect 11514 31356 11520 31408
rect 11572 31396 11578 31408
rect 12161 31399 12219 31405
rect 12161 31396 12173 31399
rect 11572 31368 12173 31396
rect 11572 31356 11578 31368
rect 12161 31365 12173 31368
rect 12207 31365 12219 31399
rect 12161 31359 12219 31365
rect 1394 31328 1400 31340
rect 1355 31300 1400 31328
rect 1394 31288 1400 31300
rect 1452 31288 1458 31340
rect 3145 31331 3203 31337
rect 3145 31297 3157 31331
rect 3191 31328 3203 31331
rect 3970 31328 3976 31340
rect 3191 31300 3976 31328
rect 3191 31297 3203 31300
rect 3145 31291 3203 31297
rect 3970 31288 3976 31300
rect 4028 31328 4034 31340
rect 4157 31331 4215 31337
rect 4157 31328 4169 31331
rect 4028 31300 4169 31328
rect 4028 31288 4034 31300
rect 4157 31297 4169 31300
rect 4203 31297 4215 31331
rect 5718 31328 5724 31340
rect 5679 31300 5724 31328
rect 4157 31291 4215 31297
rect 5718 31288 5724 31300
rect 5776 31288 5782 31340
rect 9214 31288 9220 31340
rect 9272 31328 9278 31340
rect 9582 31328 9588 31340
rect 9272 31300 9588 31328
rect 9272 31288 9278 31300
rect 9582 31288 9588 31300
rect 9640 31328 9646 31340
rect 9953 31331 10011 31337
rect 9953 31328 9965 31331
rect 9640 31300 9965 31328
rect 9640 31288 9646 31300
rect 9953 31297 9965 31300
rect 9999 31328 10011 31331
rect 12728 31328 12756 31436
rect 13081 31433 13093 31467
rect 13127 31464 13139 31467
rect 13906 31464 13912 31476
rect 13127 31436 13912 31464
rect 13127 31433 13139 31436
rect 13081 31427 13139 31433
rect 9999 31300 12756 31328
rect 9999 31297 10011 31300
rect 9953 31291 10011 31297
rect 6825 31263 6883 31269
rect 6825 31260 6837 31263
rect 5184 31232 6837 31260
rect 1670 31201 1676 31204
rect 1664 31192 1676 31201
rect 1631 31164 1676 31192
rect 1664 31155 1676 31164
rect 1670 31152 1676 31155
rect 1728 31152 1734 31204
rect 2958 31152 2964 31204
rect 3016 31192 3022 31204
rect 3694 31192 3700 31204
rect 3016 31164 3700 31192
rect 3016 31152 3022 31164
rect 3694 31152 3700 31164
rect 3752 31192 3758 31204
rect 3973 31195 4031 31201
rect 3973 31192 3985 31195
rect 3752 31164 3985 31192
rect 3752 31152 3758 31164
rect 3973 31161 3985 31164
rect 4019 31161 4031 31195
rect 3973 31155 4031 31161
rect 3602 31124 3608 31136
rect 3563 31096 3608 31124
rect 3602 31084 3608 31096
rect 3660 31084 3666 31136
rect 4062 31124 4068 31136
rect 4023 31096 4068 31124
rect 4062 31084 4068 31096
rect 4120 31084 4126 31136
rect 5074 31124 5080 31136
rect 5035 31096 5080 31124
rect 5074 31084 5080 31096
rect 5132 31084 5138 31136
rect 5184 31133 5212 31232
rect 6825 31229 6837 31232
rect 6871 31260 6883 31263
rect 7377 31263 7435 31269
rect 7377 31260 7389 31263
rect 6871 31232 7389 31260
rect 6871 31229 6883 31232
rect 6825 31223 6883 31229
rect 7377 31229 7389 31232
rect 7423 31229 7435 31263
rect 7377 31223 7435 31229
rect 8205 31263 8263 31269
rect 8205 31229 8217 31263
rect 8251 31260 8263 31263
rect 8662 31260 8668 31272
rect 8251 31232 8668 31260
rect 8251 31229 8263 31232
rect 8205 31223 8263 31229
rect 8662 31220 8668 31232
rect 8720 31260 8726 31272
rect 8941 31263 8999 31269
rect 8941 31260 8953 31263
rect 8720 31232 8953 31260
rect 8720 31220 8726 31232
rect 8941 31229 8953 31232
rect 8987 31260 8999 31263
rect 10505 31263 10563 31269
rect 8987 31232 9996 31260
rect 8987 31229 8999 31232
rect 8941 31223 8999 31229
rect 5258 31152 5264 31204
rect 5316 31192 5322 31204
rect 5629 31195 5687 31201
rect 5629 31192 5641 31195
rect 5316 31164 5641 31192
rect 5316 31152 5322 31164
rect 5629 31161 5641 31164
rect 5675 31161 5687 31195
rect 5629 31155 5687 31161
rect 9309 31195 9367 31201
rect 9309 31161 9321 31195
rect 9355 31192 9367 31195
rect 9858 31192 9864 31204
rect 9355 31164 9864 31192
rect 9355 31161 9367 31164
rect 9309 31155 9367 31161
rect 9858 31152 9864 31164
rect 9916 31152 9922 31204
rect 9968 31192 9996 31232
rect 10505 31229 10517 31263
rect 10551 31260 10563 31263
rect 11146 31260 11152 31272
rect 10551 31232 11152 31260
rect 10551 31229 10563 31232
rect 10505 31223 10563 31229
rect 11146 31220 11152 31232
rect 11204 31220 11210 31272
rect 11241 31263 11299 31269
rect 11241 31229 11253 31263
rect 11287 31260 11299 31263
rect 11882 31260 11888 31272
rect 11287 31232 11888 31260
rect 11287 31229 11299 31232
rect 11241 31223 11299 31229
rect 11882 31220 11888 31232
rect 11940 31220 11946 31272
rect 12437 31263 12495 31269
rect 12437 31229 12449 31263
rect 12483 31260 12495 31263
rect 13096 31260 13124 31427
rect 13906 31424 13912 31436
rect 13964 31424 13970 31476
rect 16482 31464 16488 31476
rect 16443 31436 16488 31464
rect 16482 31424 16488 31436
rect 16540 31424 16546 31476
rect 17034 31464 17040 31476
rect 16995 31436 17040 31464
rect 17034 31424 17040 31436
rect 17092 31424 17098 31476
rect 17862 31464 17868 31476
rect 17823 31436 17868 31464
rect 17862 31424 17868 31436
rect 17920 31424 17926 31476
rect 18598 31464 18604 31476
rect 18559 31436 18604 31464
rect 18598 31424 18604 31436
rect 18656 31424 18662 31476
rect 20806 31464 20812 31476
rect 20767 31436 20812 31464
rect 20806 31424 20812 31436
rect 20864 31424 20870 31476
rect 21453 31467 21511 31473
rect 21453 31433 21465 31467
rect 21499 31464 21511 31467
rect 21818 31464 21824 31476
rect 21499 31436 21824 31464
rect 21499 31433 21511 31436
rect 21453 31427 21511 31433
rect 21818 31424 21824 31436
rect 21876 31424 21882 31476
rect 23382 31464 23388 31476
rect 23343 31436 23388 31464
rect 23382 31424 23388 31436
rect 23440 31424 23446 31476
rect 24121 31467 24179 31473
rect 24121 31433 24133 31467
rect 24167 31464 24179 31467
rect 24762 31464 24768 31476
rect 24167 31436 24768 31464
rect 24167 31433 24179 31436
rect 24121 31427 24179 31433
rect 24762 31424 24768 31436
rect 24820 31424 24826 31476
rect 25130 31424 25136 31476
rect 25188 31464 25194 31476
rect 25593 31467 25651 31473
rect 25593 31464 25605 31467
rect 25188 31436 25605 31464
rect 25188 31424 25194 31436
rect 25593 31433 25605 31436
rect 25639 31433 25651 31467
rect 26234 31464 26240 31476
rect 26195 31436 26240 31464
rect 25593 31427 25651 31433
rect 26234 31424 26240 31436
rect 26292 31424 26298 31476
rect 26694 31464 26700 31476
rect 26655 31436 26700 31464
rect 26694 31424 26700 31436
rect 26752 31424 26758 31476
rect 14737 31399 14795 31405
rect 14737 31365 14749 31399
rect 14783 31396 14795 31399
rect 16574 31396 16580 31408
rect 14783 31368 16580 31396
rect 14783 31365 14795 31368
rect 14737 31359 14795 31365
rect 16574 31356 16580 31368
rect 16632 31396 16638 31408
rect 16853 31399 16911 31405
rect 16853 31396 16865 31399
rect 16632 31368 16865 31396
rect 16632 31356 16638 31368
rect 16853 31365 16865 31368
rect 16899 31365 16911 31399
rect 16853 31359 16911 31365
rect 25317 31399 25375 31405
rect 25317 31365 25329 31399
rect 25363 31396 25375 31399
rect 26050 31396 26056 31408
rect 25363 31368 26056 31396
rect 25363 31365 25375 31368
rect 25317 31359 25375 31365
rect 13538 31260 13544 31272
rect 12483 31232 13124 31260
rect 13451 31232 13544 31260
rect 12483 31229 12495 31232
rect 12437 31223 12495 31229
rect 13538 31220 13544 31232
rect 13596 31260 13602 31272
rect 14093 31263 14151 31269
rect 14093 31260 14105 31263
rect 13596 31232 14105 31260
rect 13596 31220 13602 31232
rect 14093 31229 14105 31232
rect 14139 31229 14151 31263
rect 14093 31223 14151 31229
rect 14366 31220 14372 31272
rect 14424 31260 14430 31272
rect 14921 31263 14979 31269
rect 14921 31260 14933 31263
rect 14424 31232 14933 31260
rect 14424 31220 14430 31232
rect 14921 31229 14933 31232
rect 14967 31260 14979 31263
rect 15197 31263 15255 31269
rect 15197 31260 15209 31263
rect 14967 31232 15209 31260
rect 14967 31229 14979 31232
rect 14921 31223 14979 31229
rect 15197 31229 15209 31232
rect 15243 31229 15255 31263
rect 15470 31260 15476 31272
rect 15383 31232 15476 31260
rect 15197 31223 15255 31229
rect 15470 31220 15476 31232
rect 15528 31260 15534 31272
rect 16025 31263 16083 31269
rect 16025 31260 16037 31263
rect 15528 31232 16037 31260
rect 15528 31220 15534 31232
rect 16025 31229 16037 31232
rect 16071 31229 16083 31263
rect 16868 31260 16896 31359
rect 22002 31328 22008 31340
rect 21963 31300 22008 31328
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 17221 31263 17279 31269
rect 17221 31260 17233 31263
rect 16868 31232 17233 31260
rect 16025 31223 16083 31229
rect 17221 31229 17233 31232
rect 17267 31229 17279 31263
rect 17221 31223 17279 31229
rect 20806 31220 20812 31272
rect 20864 31260 20870 31272
rect 21821 31263 21879 31269
rect 21821 31260 21833 31263
rect 20864 31232 21833 31260
rect 20864 31220 20870 31232
rect 21821 31229 21833 31232
rect 21867 31229 21879 31263
rect 21821 31223 21879 31229
rect 24581 31263 24639 31269
rect 24581 31229 24593 31263
rect 24627 31260 24639 31263
rect 25332 31260 25360 31359
rect 26050 31356 26056 31368
rect 26108 31356 26114 31408
rect 26252 31328 26280 31424
rect 26252 31300 26924 31328
rect 24627 31232 25360 31260
rect 24627 31229 24639 31232
rect 24581 31223 24639 31229
rect 26602 31220 26608 31272
rect 26660 31260 26666 31272
rect 26786 31260 26792 31272
rect 26660 31232 26792 31260
rect 26660 31220 26666 31232
rect 26786 31220 26792 31232
rect 26844 31220 26850 31272
rect 26896 31260 26924 31300
rect 27045 31263 27103 31269
rect 27045 31260 27057 31263
rect 26896 31232 27057 31260
rect 27045 31229 27057 31232
rect 27091 31260 27103 31263
rect 28442 31260 28448 31272
rect 27091 31232 28448 31260
rect 27091 31229 27103 31232
rect 27045 31223 27103 31229
rect 28442 31220 28448 31232
rect 28500 31220 28506 31272
rect 18138 31192 18144 31204
rect 9968 31164 11008 31192
rect 5169 31127 5227 31133
rect 5169 31093 5181 31127
rect 5215 31093 5227 31127
rect 5169 31087 5227 31093
rect 5350 31084 5356 31136
rect 5408 31124 5414 31136
rect 5537 31127 5595 31133
rect 5537 31124 5549 31127
rect 5408 31096 5549 31124
rect 5408 31084 5414 31096
rect 5537 31093 5549 31096
rect 5583 31093 5595 31127
rect 5537 31087 5595 31093
rect 9401 31127 9459 31133
rect 9401 31093 9413 31127
rect 9447 31124 9459 31127
rect 9582 31124 9588 31136
rect 9447 31096 9588 31124
rect 9447 31093 9459 31096
rect 9401 31087 9459 31093
rect 9582 31084 9588 31096
rect 9640 31084 9646 31136
rect 9766 31124 9772 31136
rect 9727 31096 9772 31124
rect 9766 31084 9772 31096
rect 9824 31084 9830 31136
rect 10980 31133 11008 31164
rect 15672 31164 18144 31192
rect 10965 31127 11023 31133
rect 10965 31093 10977 31127
rect 11011 31093 11023 31127
rect 10965 31087 11023 31093
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 11425 31127 11483 31133
rect 11425 31124 11437 31127
rect 11388 31096 11437 31124
rect 11388 31084 11394 31096
rect 11425 31093 11437 31096
rect 11471 31093 11483 31127
rect 11425 31087 11483 31093
rect 13078 31084 13084 31136
rect 13136 31124 13142 31136
rect 15672 31133 15700 31164
rect 18138 31152 18144 31164
rect 18196 31192 18202 31204
rect 18233 31195 18291 31201
rect 18233 31192 18245 31195
rect 18196 31164 18245 31192
rect 18196 31152 18202 31164
rect 18233 31161 18245 31164
rect 18279 31161 18291 31195
rect 18233 31155 18291 31161
rect 21177 31195 21235 31201
rect 21177 31161 21189 31195
rect 21223 31192 21235 31195
rect 21634 31192 21640 31204
rect 21223 31164 21640 31192
rect 21223 31161 21235 31164
rect 21177 31155 21235 31161
rect 21634 31152 21640 31164
rect 21692 31192 21698 31204
rect 21913 31195 21971 31201
rect 21913 31192 21925 31195
rect 21692 31164 21925 31192
rect 21692 31152 21698 31164
rect 21913 31161 21925 31164
rect 21959 31161 21971 31195
rect 21913 31155 21971 31161
rect 24489 31195 24547 31201
rect 24489 31161 24501 31195
rect 24535 31192 24547 31195
rect 24762 31192 24768 31204
rect 24535 31164 24768 31192
rect 24535 31161 24547 31164
rect 24489 31155 24547 31161
rect 24762 31152 24768 31164
rect 24820 31152 24826 31204
rect 13725 31127 13783 31133
rect 13725 31124 13737 31127
rect 13136 31096 13737 31124
rect 13136 31084 13142 31096
rect 13725 31093 13737 31096
rect 13771 31093 13783 31127
rect 13725 31087 13783 31093
rect 15657 31127 15715 31133
rect 15657 31093 15669 31127
rect 15703 31093 15715 31127
rect 15657 31087 15715 31093
rect 24949 31127 25007 31133
rect 24949 31093 24961 31127
rect 24995 31124 25007 31127
rect 25130 31124 25136 31136
rect 24995 31096 25136 31124
rect 24995 31093 25007 31096
rect 24949 31087 25007 31093
rect 25130 31084 25136 31096
rect 25188 31084 25194 31136
rect 28166 31124 28172 31136
rect 28127 31096 28172 31124
rect 28166 31084 28172 31096
rect 28224 31084 28230 31136
rect 35434 31124 35440 31136
rect 35395 31096 35440 31124
rect 35434 31084 35440 31096
rect 35492 31084 35498 31136
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 2041 30923 2099 30929
rect 2041 30889 2053 30923
rect 2087 30920 2099 30923
rect 2498 30920 2504 30932
rect 2087 30892 2504 30920
rect 2087 30889 2099 30892
rect 2041 30883 2099 30889
rect 2498 30880 2504 30892
rect 2556 30880 2562 30932
rect 2774 30880 2780 30932
rect 2832 30920 2838 30932
rect 3697 30923 3755 30929
rect 3697 30920 3709 30923
rect 2832 30892 3709 30920
rect 2832 30880 2838 30892
rect 3697 30889 3709 30892
rect 3743 30920 3755 30923
rect 4062 30920 4068 30932
rect 3743 30892 4068 30920
rect 3743 30889 3755 30892
rect 3697 30883 3755 30889
rect 4062 30880 4068 30892
rect 4120 30880 4126 30932
rect 4433 30923 4491 30929
rect 4433 30889 4445 30923
rect 4479 30920 4491 30923
rect 5442 30920 5448 30932
rect 4479 30892 5448 30920
rect 4479 30889 4491 30892
rect 4433 30883 4491 30889
rect 5442 30880 5448 30892
rect 5500 30880 5506 30932
rect 10689 30923 10747 30929
rect 10689 30889 10701 30923
rect 10735 30920 10747 30923
rect 11514 30920 11520 30932
rect 10735 30892 11520 30920
rect 10735 30889 10747 30892
rect 10689 30883 10747 30889
rect 1394 30812 1400 30864
rect 1452 30852 1458 30864
rect 2317 30855 2375 30861
rect 2317 30852 2329 30855
rect 1452 30824 2329 30852
rect 1452 30812 1458 30824
rect 2317 30821 2329 30824
rect 2363 30821 2375 30855
rect 2317 30815 2375 30821
rect 5620 30855 5678 30861
rect 5620 30821 5632 30855
rect 5666 30852 5678 30855
rect 6270 30852 6276 30864
rect 5666 30824 6276 30852
rect 5666 30821 5678 30824
rect 5620 30815 5678 30821
rect 6270 30812 6276 30824
rect 6328 30812 6334 30864
rect 3602 30744 3608 30796
rect 3660 30784 3666 30796
rect 3970 30784 3976 30796
rect 3660 30756 3976 30784
rect 3660 30744 3666 30756
rect 3970 30744 3976 30756
rect 4028 30784 4034 30796
rect 4249 30787 4307 30793
rect 4249 30784 4261 30787
rect 4028 30756 4261 30784
rect 4028 30744 4034 30756
rect 4249 30753 4261 30756
rect 4295 30753 4307 30787
rect 4890 30784 4896 30796
rect 4803 30756 4896 30784
rect 4249 30747 4307 30753
rect 4890 30744 4896 30756
rect 4948 30784 4954 30796
rect 5442 30784 5448 30796
rect 4948 30756 5448 30784
rect 4948 30744 4954 30756
rect 5442 30744 5448 30756
rect 5500 30744 5506 30796
rect 8662 30784 8668 30796
rect 8623 30756 8668 30784
rect 8662 30744 8668 30756
rect 8720 30744 8726 30796
rect 9677 30787 9735 30793
rect 9677 30753 9689 30787
rect 9723 30784 9735 30787
rect 9950 30784 9956 30796
rect 9723 30756 9956 30784
rect 9723 30753 9735 30756
rect 9677 30747 9735 30753
rect 9950 30744 9956 30756
rect 10008 30784 10014 30796
rect 10796 30793 10824 30892
rect 11514 30880 11520 30892
rect 11572 30880 11578 30932
rect 12710 30920 12716 30932
rect 12671 30892 12716 30920
rect 12710 30880 12716 30892
rect 12768 30880 12774 30932
rect 13078 30920 13084 30932
rect 13039 30892 13084 30920
rect 13078 30880 13084 30892
rect 13136 30880 13142 30932
rect 13538 30920 13544 30932
rect 13499 30892 13544 30920
rect 13538 30880 13544 30892
rect 13596 30880 13602 30932
rect 14366 30920 14372 30932
rect 14327 30892 14372 30920
rect 14366 30880 14372 30892
rect 14424 30880 14430 30932
rect 17770 30920 17776 30932
rect 17731 30892 17776 30920
rect 17770 30880 17776 30892
rect 17828 30880 17834 30932
rect 20898 30880 20904 30932
rect 20956 30920 20962 30932
rect 21085 30923 21143 30929
rect 21085 30920 21097 30923
rect 20956 30892 21097 30920
rect 20956 30880 20962 30892
rect 21085 30889 21097 30892
rect 21131 30889 21143 30923
rect 21085 30883 21143 30889
rect 21545 30923 21603 30929
rect 21545 30889 21557 30923
rect 21591 30920 21603 30923
rect 21634 30920 21640 30932
rect 21591 30892 21640 30920
rect 21591 30889 21603 30892
rect 21545 30883 21603 30889
rect 21634 30880 21640 30892
rect 21692 30880 21698 30932
rect 21913 30923 21971 30929
rect 21913 30889 21925 30923
rect 21959 30920 21971 30923
rect 22002 30920 22008 30932
rect 21959 30892 22008 30920
rect 21959 30889 21971 30892
rect 21913 30883 21971 30889
rect 22002 30880 22008 30892
rect 22060 30880 22066 30932
rect 22741 30923 22799 30929
rect 22741 30889 22753 30923
rect 22787 30920 22799 30923
rect 23290 30920 23296 30932
rect 22787 30892 23296 30920
rect 22787 30889 22799 30892
rect 22741 30883 22799 30889
rect 23290 30880 23296 30892
rect 23348 30880 23354 30932
rect 23934 30880 23940 30932
rect 23992 30920 23998 30932
rect 24305 30923 24363 30929
rect 24305 30920 24317 30923
rect 23992 30892 24317 30920
rect 23992 30880 23998 30892
rect 24305 30889 24317 30892
rect 24351 30920 24363 30923
rect 24762 30920 24768 30932
rect 24351 30892 24768 30920
rect 24351 30889 24363 30892
rect 24305 30883 24363 30889
rect 24762 30880 24768 30892
rect 24820 30880 24826 30932
rect 25498 30920 25504 30932
rect 25459 30892 25504 30920
rect 25498 30880 25504 30892
rect 25556 30880 25562 30932
rect 35618 30920 35624 30932
rect 35579 30892 35624 30920
rect 35618 30880 35624 30892
rect 35676 30880 35682 30932
rect 12897 30855 12955 30861
rect 12897 30821 12909 30855
rect 12943 30852 12955 30855
rect 13357 30855 13415 30861
rect 13357 30852 13369 30855
rect 12943 30824 13369 30852
rect 12943 30821 12955 30824
rect 12897 30815 12955 30821
rect 13357 30821 13369 30824
rect 13403 30821 13415 30855
rect 13357 30815 13415 30821
rect 15562 30812 15568 30864
rect 15620 30852 15626 30864
rect 15810 30855 15868 30861
rect 15810 30852 15822 30855
rect 15620 30824 15822 30852
rect 15620 30812 15626 30824
rect 15810 30821 15822 30824
rect 15856 30821 15868 30855
rect 15810 30815 15868 30821
rect 10229 30787 10287 30793
rect 10229 30784 10241 30787
rect 10008 30756 10241 30784
rect 10008 30744 10014 30756
rect 10229 30753 10241 30756
rect 10275 30753 10287 30787
rect 10229 30747 10287 30753
rect 10781 30787 10839 30793
rect 10781 30753 10793 30787
rect 10827 30753 10839 30787
rect 11037 30787 11095 30793
rect 11037 30784 11049 30787
rect 10781 30747 10839 30753
rect 10888 30756 11049 30784
rect 5350 30716 5356 30728
rect 5311 30688 5356 30716
rect 5350 30676 5356 30688
rect 5408 30676 5414 30728
rect 9493 30719 9551 30725
rect 9493 30685 9505 30719
rect 9539 30716 9551 30719
rect 9766 30716 9772 30728
rect 9539 30688 9772 30716
rect 9539 30685 9551 30688
rect 9493 30679 9551 30685
rect 9766 30676 9772 30688
rect 9824 30716 9830 30728
rect 10686 30716 10692 30728
rect 9824 30688 10692 30716
rect 9824 30676 9830 30688
rect 10686 30676 10692 30688
rect 10744 30716 10750 30728
rect 10888 30716 10916 30756
rect 11037 30753 11049 30756
rect 11083 30753 11095 30787
rect 11037 30747 11095 30753
rect 13173 30787 13231 30793
rect 13173 30753 13185 30787
rect 13219 30784 13231 30787
rect 13722 30784 13728 30796
rect 13219 30756 13728 30784
rect 13219 30753 13231 30756
rect 13173 30747 13231 30753
rect 13722 30744 13728 30756
rect 13780 30744 13786 30796
rect 14550 30784 14556 30796
rect 14511 30756 14556 30784
rect 14550 30744 14556 30756
rect 14608 30744 14614 30796
rect 15105 30787 15163 30793
rect 15105 30753 15117 30787
rect 15151 30784 15163 30787
rect 17034 30784 17040 30796
rect 15151 30756 17040 30784
rect 15151 30753 15163 30756
rect 15105 30747 15163 30753
rect 15580 30725 15608 30756
rect 17034 30744 17040 30756
rect 17092 30744 17098 30796
rect 17497 30787 17555 30793
rect 17497 30753 17509 30787
rect 17543 30784 17555 30787
rect 18141 30787 18199 30793
rect 18141 30784 18153 30787
rect 17543 30756 18153 30784
rect 17543 30753 17555 30756
rect 17497 30747 17555 30753
rect 18141 30753 18153 30756
rect 18187 30753 18199 30787
rect 18141 30747 18199 30753
rect 18233 30787 18291 30793
rect 18233 30753 18245 30787
rect 18279 30784 18291 30787
rect 18782 30784 18788 30796
rect 18279 30756 18788 30784
rect 18279 30753 18291 30756
rect 18233 30747 18291 30753
rect 18782 30744 18788 30756
rect 18840 30744 18846 30796
rect 22554 30784 22560 30796
rect 22515 30756 22560 30784
rect 22554 30744 22560 30756
rect 22612 30744 22618 30796
rect 25130 30744 25136 30796
rect 25188 30784 25194 30796
rect 26510 30784 26516 30796
rect 25188 30756 26516 30784
rect 25188 30744 25194 30756
rect 26510 30744 26516 30756
rect 26568 30744 26574 30796
rect 35437 30787 35495 30793
rect 35437 30753 35449 30787
rect 35483 30784 35495 30787
rect 35618 30784 35624 30796
rect 35483 30756 35624 30784
rect 35483 30753 35495 30756
rect 35437 30747 35495 30753
rect 35618 30744 35624 30756
rect 35676 30744 35682 30796
rect 10744 30688 10916 30716
rect 15565 30719 15623 30725
rect 10744 30676 10750 30688
rect 15565 30685 15577 30719
rect 15611 30685 15623 30719
rect 17770 30716 17776 30728
rect 15565 30679 15623 30685
rect 16960 30688 17776 30716
rect 1670 30648 1676 30660
rect 1631 30620 1676 30648
rect 1670 30608 1676 30620
rect 1728 30608 1734 30660
rect 7006 30648 7012 30660
rect 6967 30620 7012 30648
rect 7006 30608 7012 30620
rect 7064 30608 7070 30660
rect 9861 30651 9919 30657
rect 9861 30617 9873 30651
rect 9907 30648 9919 30651
rect 12161 30651 12219 30657
rect 9907 30620 10824 30648
rect 9907 30617 9919 30620
rect 9861 30611 9919 30617
rect 3050 30580 3056 30592
rect 3011 30552 3056 30580
rect 3050 30540 3056 30552
rect 3108 30540 3114 30592
rect 5258 30580 5264 30592
rect 5219 30552 5264 30580
rect 5258 30540 5264 30552
rect 5316 30540 5322 30592
rect 6730 30580 6736 30592
rect 6691 30552 6736 30580
rect 6730 30540 6736 30552
rect 6788 30540 6794 30592
rect 8478 30580 8484 30592
rect 8439 30552 8484 30580
rect 8478 30540 8484 30552
rect 8536 30540 8542 30592
rect 10796 30580 10824 30620
rect 12161 30617 12173 30651
rect 12207 30648 12219 30651
rect 12894 30648 12900 30660
rect 12207 30620 12900 30648
rect 12207 30617 12219 30620
rect 12161 30611 12219 30617
rect 12894 30608 12900 30620
rect 12952 30608 12958 30660
rect 16960 30657 16988 30688
rect 17770 30676 17776 30688
rect 17828 30716 17834 30728
rect 18322 30716 18328 30728
rect 17828 30688 18328 30716
rect 17828 30676 17834 30688
rect 18322 30676 18328 30688
rect 18380 30676 18386 30728
rect 23658 30676 23664 30728
rect 23716 30716 23722 30728
rect 24857 30719 24915 30725
rect 24857 30716 24869 30719
rect 23716 30688 24869 30716
rect 23716 30676 23722 30688
rect 24857 30685 24869 30688
rect 24903 30685 24915 30719
rect 24857 30679 24915 30685
rect 25041 30719 25099 30725
rect 25041 30685 25053 30719
rect 25087 30716 25099 30719
rect 25087 30688 26740 30716
rect 25087 30685 25099 30688
rect 25041 30679 25099 30685
rect 16945 30651 17003 30657
rect 16945 30617 16957 30651
rect 16991 30617 17003 30651
rect 16945 30611 17003 30617
rect 24118 30608 24124 30660
rect 24176 30648 24182 30660
rect 25056 30648 25084 30679
rect 26712 30657 26740 30688
rect 24176 30620 25084 30648
rect 26697 30651 26755 30657
rect 24176 30608 24182 30620
rect 26697 30617 26709 30651
rect 26743 30617 26755 30651
rect 26697 30611 26755 30617
rect 11054 30580 11060 30592
rect 10796 30552 11060 30580
rect 11054 30540 11060 30552
rect 11112 30540 11118 30592
rect 14274 30580 14280 30592
rect 14235 30552 14280 30580
rect 14274 30540 14280 30552
rect 14332 30540 14338 30592
rect 16574 30540 16580 30592
rect 16632 30580 16638 30592
rect 17221 30583 17279 30589
rect 17221 30580 17233 30583
rect 16632 30552 17233 30580
rect 16632 30540 16638 30552
rect 17221 30549 17233 30552
rect 17267 30580 17279 30583
rect 17497 30583 17555 30589
rect 17497 30580 17509 30583
rect 17267 30552 17509 30580
rect 17267 30549 17279 30552
rect 17221 30543 17279 30549
rect 17497 30549 17509 30552
rect 17543 30580 17555 30583
rect 17589 30583 17647 30589
rect 17589 30580 17601 30583
rect 17543 30552 17601 30580
rect 17543 30549 17555 30552
rect 17497 30543 17555 30549
rect 17589 30549 17601 30552
rect 17635 30549 17647 30583
rect 18874 30580 18880 30592
rect 18835 30552 18880 30580
rect 17589 30543 17647 30549
rect 18874 30540 18880 30552
rect 18932 30540 18938 30592
rect 24394 30580 24400 30592
rect 24355 30552 24400 30580
rect 24394 30540 24400 30552
rect 24452 30540 24458 30592
rect 26602 30540 26608 30592
rect 26660 30580 26666 30592
rect 27065 30583 27123 30589
rect 27065 30580 27077 30583
rect 26660 30552 27077 30580
rect 26660 30540 26666 30552
rect 27065 30549 27077 30552
rect 27111 30580 27123 30583
rect 27433 30583 27491 30589
rect 27433 30580 27445 30583
rect 27111 30552 27445 30580
rect 27111 30549 27123 30552
rect 27065 30543 27123 30549
rect 27433 30549 27445 30552
rect 27479 30549 27491 30583
rect 27433 30543 27491 30549
rect 32493 30583 32551 30589
rect 32493 30549 32505 30583
rect 32539 30580 32551 30583
rect 33042 30580 33048 30592
rect 32539 30552 33048 30580
rect 32539 30549 32551 30552
rect 32493 30543 32551 30549
rect 33042 30540 33048 30552
rect 33100 30540 33106 30592
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 1394 30336 1400 30388
rect 1452 30376 1458 30388
rect 1581 30379 1639 30385
rect 1581 30376 1593 30379
rect 1452 30348 1593 30376
rect 1452 30336 1458 30348
rect 1581 30345 1593 30348
rect 1627 30345 1639 30379
rect 2958 30376 2964 30388
rect 2919 30348 2964 30376
rect 1581 30339 1639 30345
rect 2958 30336 2964 30348
rect 3016 30336 3022 30388
rect 3970 30376 3976 30388
rect 3931 30348 3976 30376
rect 3970 30336 3976 30348
rect 4028 30336 4034 30388
rect 4890 30376 4896 30388
rect 4080 30348 4896 30376
rect 2314 30268 2320 30320
rect 2372 30308 2378 30320
rect 2501 30311 2559 30317
rect 2501 30308 2513 30311
rect 2372 30280 2513 30308
rect 2372 30268 2378 30280
rect 2501 30277 2513 30280
rect 2547 30308 2559 30311
rect 4080 30308 4108 30348
rect 4890 30336 4896 30348
rect 4948 30336 4954 30388
rect 5258 30336 5264 30388
rect 5316 30376 5322 30388
rect 6825 30379 6883 30385
rect 6825 30376 6837 30379
rect 5316 30348 6837 30376
rect 5316 30336 5322 30348
rect 6825 30345 6837 30348
rect 6871 30345 6883 30379
rect 9858 30376 9864 30388
rect 9819 30348 9864 30376
rect 6825 30339 6883 30345
rect 9858 30336 9864 30348
rect 9916 30336 9922 30388
rect 13722 30376 13728 30388
rect 13683 30348 13728 30376
rect 13722 30336 13728 30348
rect 13780 30336 13786 30388
rect 18874 30376 18880 30388
rect 18064 30348 18880 30376
rect 5902 30308 5908 30320
rect 2547 30280 4108 30308
rect 5863 30280 5908 30308
rect 2547 30277 2559 30280
rect 2501 30271 2559 30277
rect 3528 30249 3556 30280
rect 5902 30268 5908 30280
rect 5960 30268 5966 30320
rect 10778 30308 10784 30320
rect 10739 30280 10784 30308
rect 10778 30268 10784 30280
rect 10836 30268 10842 30320
rect 3513 30243 3571 30249
rect 3513 30209 3525 30243
rect 3559 30209 3571 30243
rect 3513 30203 3571 30209
rect 5534 30200 5540 30252
rect 5592 30240 5598 30252
rect 5994 30240 6000 30252
rect 5592 30212 6000 30240
rect 5592 30200 5598 30212
rect 5994 30200 6000 30212
rect 6052 30240 6058 30252
rect 7469 30243 7527 30249
rect 7469 30240 7481 30243
rect 6052 30212 7481 30240
rect 6052 30200 6058 30212
rect 7469 30209 7481 30212
rect 7515 30240 7527 30243
rect 7837 30243 7895 30249
rect 7837 30240 7849 30243
rect 7515 30212 7849 30240
rect 7515 30209 7527 30212
rect 7469 30203 7527 30209
rect 7837 30209 7849 30212
rect 7883 30209 7895 30243
rect 11422 30240 11428 30252
rect 11383 30212 11428 30240
rect 7837 30203 7895 30209
rect 11422 30200 11428 30212
rect 11480 30200 11486 30252
rect 13078 30200 13084 30252
rect 13136 30240 13142 30252
rect 13173 30243 13231 30249
rect 13173 30240 13185 30243
rect 13136 30212 13185 30240
rect 13136 30200 13142 30212
rect 13173 30209 13185 30212
rect 13219 30209 13231 30243
rect 13173 30203 13231 30209
rect 16482 30200 16488 30252
rect 16540 30240 16546 30252
rect 16945 30243 17003 30249
rect 16945 30240 16957 30243
rect 16540 30212 16957 30240
rect 16540 30200 16546 30212
rect 16945 30209 16957 30212
rect 16991 30240 17003 30243
rect 17310 30240 17316 30252
rect 16991 30212 17316 30240
rect 16991 30209 17003 30212
rect 16945 30203 17003 30209
rect 17310 30200 17316 30212
rect 17368 30200 17374 30252
rect 18064 30249 18092 30348
rect 18874 30336 18880 30348
rect 18932 30336 18938 30388
rect 21634 30336 21640 30388
rect 21692 30376 21698 30388
rect 22554 30376 22560 30388
rect 21692 30348 22048 30376
rect 22515 30348 22560 30376
rect 21692 30336 21698 30348
rect 22020 30308 22048 30348
rect 22554 30336 22560 30348
rect 22612 30336 22618 30388
rect 24670 30376 24676 30388
rect 24631 30348 24676 30376
rect 24670 30336 24676 30348
rect 24728 30336 24734 30388
rect 26510 30376 26516 30388
rect 26471 30348 26516 30376
rect 26510 30336 26516 30348
rect 26568 30336 26574 30388
rect 22097 30311 22155 30317
rect 22097 30308 22109 30311
rect 22020 30280 22109 30308
rect 22097 30277 22109 30280
rect 22143 30277 22155 30311
rect 22097 30271 22155 30277
rect 18049 30243 18107 30249
rect 18049 30209 18061 30243
rect 18095 30209 18107 30243
rect 18049 30203 18107 30209
rect 18230 30200 18236 30252
rect 18288 30240 18294 30252
rect 18512 30243 18570 30249
rect 18512 30240 18524 30243
rect 18288 30212 18524 30240
rect 18288 30200 18294 30212
rect 18512 30209 18524 30212
rect 18558 30209 18570 30243
rect 18782 30240 18788 30252
rect 18743 30212 18788 30240
rect 18512 30203 18570 30209
rect 18782 30200 18788 30212
rect 18840 30200 18846 30252
rect 24688 30240 24716 30336
rect 35621 30311 35679 30317
rect 35621 30277 35633 30311
rect 35667 30308 35679 30311
rect 35710 30308 35716 30320
rect 35667 30280 35716 30308
rect 35667 30277 35679 30280
rect 35621 30271 35679 30277
rect 35710 30268 35716 30280
rect 35768 30268 35774 30320
rect 33042 30240 33048 30252
rect 24688 30212 24900 30240
rect 33003 30212 33048 30240
rect 3050 30132 3056 30184
rect 3108 30172 3114 30184
rect 3329 30175 3387 30181
rect 3329 30172 3341 30175
rect 3108 30144 3341 30172
rect 3108 30132 3114 30144
rect 3329 30141 3341 30144
rect 3375 30141 3387 30175
rect 3329 30135 3387 30141
rect 4525 30175 4583 30181
rect 4525 30141 4537 30175
rect 4571 30172 4583 30175
rect 5350 30172 5356 30184
rect 4571 30144 5356 30172
rect 4571 30141 4583 30144
rect 4525 30135 4583 30141
rect 5350 30132 5356 30144
rect 5408 30172 5414 30184
rect 6454 30172 6460 30184
rect 5408 30144 6460 30172
rect 5408 30132 5414 30144
rect 6454 30132 6460 30144
rect 6512 30132 6518 30184
rect 7006 30132 7012 30184
rect 7064 30172 7070 30184
rect 7193 30175 7251 30181
rect 7193 30172 7205 30175
rect 7064 30144 7205 30172
rect 7064 30132 7070 30144
rect 7193 30141 7205 30144
rect 7239 30141 7251 30175
rect 7193 30135 7251 30141
rect 8481 30175 8539 30181
rect 8481 30141 8493 30175
rect 8527 30172 8539 30175
rect 8570 30172 8576 30184
rect 8527 30144 8576 30172
rect 8527 30141 8539 30144
rect 8481 30135 8539 30141
rect 8570 30132 8576 30144
rect 8628 30132 8634 30184
rect 11054 30132 11060 30184
rect 11112 30172 11118 30184
rect 11149 30175 11207 30181
rect 11149 30172 11161 30175
rect 11112 30144 11161 30172
rect 11112 30132 11118 30144
rect 11149 30141 11161 30144
rect 11195 30172 11207 30175
rect 11793 30175 11851 30181
rect 11793 30172 11805 30175
rect 11195 30144 11805 30172
rect 11195 30141 11207 30144
rect 11149 30135 11207 30141
rect 11793 30141 11805 30144
rect 11839 30141 11851 30175
rect 11793 30135 11851 30141
rect 12894 30132 12900 30184
rect 12952 30172 12958 30184
rect 14001 30175 14059 30181
rect 14001 30172 14013 30175
rect 12952 30144 14013 30172
rect 12952 30132 12958 30144
rect 14001 30141 14013 30144
rect 14047 30141 14059 30175
rect 14182 30172 14188 30184
rect 14143 30144 14188 30172
rect 14001 30135 14059 30141
rect 14182 30132 14188 30144
rect 14240 30132 14246 30184
rect 14274 30132 14280 30184
rect 14332 30172 14338 30184
rect 14441 30175 14499 30181
rect 14441 30172 14453 30175
rect 14332 30144 14453 30172
rect 14332 30132 14338 30144
rect 14441 30141 14453 30144
rect 14487 30141 14499 30175
rect 14441 30135 14499 30141
rect 16301 30175 16359 30181
rect 16301 30141 16313 30175
rect 16347 30172 16359 30175
rect 16758 30172 16764 30184
rect 16347 30144 16764 30172
rect 16347 30141 16359 30144
rect 16301 30135 16359 30141
rect 16758 30132 16764 30144
rect 16816 30132 16822 30184
rect 18414 30132 18420 30184
rect 18472 30172 18478 30184
rect 20257 30175 20315 30181
rect 18472 30144 19932 30172
rect 18472 30132 18478 30144
rect 2869 30107 2927 30113
rect 2869 30073 2881 30107
rect 2915 30104 2927 30107
rect 3421 30107 3479 30113
rect 3421 30104 3433 30107
rect 2915 30076 3433 30104
rect 2915 30073 2927 30076
rect 2869 30067 2927 30073
rect 3421 30073 3433 30076
rect 3467 30104 3479 30107
rect 4062 30104 4068 30116
rect 3467 30076 4068 30104
rect 3467 30073 3479 30076
rect 3421 30067 3479 30073
rect 4062 30064 4068 30076
rect 4120 30064 4126 30116
rect 4433 30107 4491 30113
rect 4433 30073 4445 30107
rect 4479 30104 4491 30107
rect 4770 30107 4828 30113
rect 4770 30104 4782 30107
rect 4479 30076 4782 30104
rect 4479 30073 4491 30076
rect 4433 30067 4491 30073
rect 4770 30073 4782 30076
rect 4816 30104 4828 30107
rect 6549 30107 6607 30113
rect 6549 30104 6561 30107
rect 4816 30076 6561 30104
rect 4816 30073 4828 30076
rect 4770 30067 4828 30073
rect 6549 30073 6561 30076
rect 6595 30104 6607 30107
rect 6730 30104 6736 30116
rect 6595 30076 6736 30104
rect 6595 30073 6607 30076
rect 6549 30067 6607 30073
rect 6730 30064 6736 30076
rect 6788 30104 6794 30116
rect 7285 30107 7343 30113
rect 7285 30104 7297 30107
rect 6788 30076 7297 30104
rect 6788 30064 6794 30076
rect 7285 30073 7297 30076
rect 7331 30073 7343 30107
rect 8726 30107 8784 30113
rect 8726 30104 8738 30107
rect 7285 30067 7343 30073
rect 8404 30076 8738 30104
rect 8404 30048 8432 30076
rect 8726 30073 8738 30076
rect 8772 30073 8784 30107
rect 11241 30107 11299 30113
rect 11241 30104 11253 30107
rect 8726 30067 8784 30073
rect 10244 30076 11253 30104
rect 10244 30048 10272 30076
rect 11241 30073 11253 30076
rect 11287 30073 11299 30107
rect 11241 30067 11299 30073
rect 12253 30107 12311 30113
rect 12253 30073 12265 30107
rect 12299 30104 12311 30107
rect 12434 30104 12440 30116
rect 12299 30076 12440 30104
rect 12299 30073 12311 30076
rect 12253 30067 12311 30073
rect 12434 30064 12440 30076
rect 12492 30104 12498 30116
rect 13081 30107 13139 30113
rect 13081 30104 13093 30107
rect 12492 30076 13093 30104
rect 12492 30064 12498 30076
rect 13081 30073 13093 30076
rect 13127 30073 13139 30107
rect 13081 30067 13139 30073
rect 15654 30064 15660 30116
rect 15712 30104 15718 30116
rect 17773 30107 17831 30113
rect 17773 30104 17785 30107
rect 15712 30076 17785 30104
rect 15712 30064 15718 30076
rect 17773 30073 17785 30076
rect 17819 30073 17831 30107
rect 17773 30067 17831 30073
rect 6270 30036 6276 30048
rect 6231 30008 6276 30036
rect 6270 29996 6276 30008
rect 6328 29996 6334 30048
rect 8386 30036 8392 30048
rect 8347 30008 8392 30036
rect 8386 29996 8392 30008
rect 8444 29996 8450 30048
rect 10226 30036 10232 30048
rect 10187 30008 10232 30036
rect 10226 29996 10232 30008
rect 10284 29996 10290 30048
rect 10686 30036 10692 30048
rect 10647 30008 10692 30036
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 12618 30036 12624 30048
rect 12579 30008 12624 30036
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 12710 29996 12716 30048
rect 12768 30036 12774 30048
rect 12989 30039 13047 30045
rect 12989 30036 13001 30039
rect 12768 30008 13001 30036
rect 12768 29996 12774 30008
rect 12989 30005 13001 30008
rect 13035 30005 13047 30039
rect 15562 30036 15568 30048
rect 15523 30008 15568 30036
rect 12989 29999 13047 30005
rect 15562 29996 15568 30008
rect 15620 30036 15626 30048
rect 15841 30039 15899 30045
rect 15841 30036 15853 30039
rect 15620 30008 15853 30036
rect 15620 29996 15626 30008
rect 15841 30005 15853 30008
rect 15887 30005 15899 30039
rect 16390 30036 16396 30048
rect 16351 30008 16396 30036
rect 15841 29999 15899 30005
rect 16390 29996 16396 30008
rect 16448 29996 16454 30048
rect 16574 29996 16580 30048
rect 16632 30036 16638 30048
rect 16853 30039 16911 30045
rect 16853 30036 16865 30039
rect 16632 30008 16865 30036
rect 16632 29996 16638 30008
rect 16853 30005 16865 30008
rect 16899 30005 16911 30039
rect 17494 30036 17500 30048
rect 17455 30008 17500 30036
rect 16853 29999 16911 30005
rect 17494 29996 17500 30008
rect 17552 29996 17558 30048
rect 17788 30036 17816 30067
rect 18515 30039 18573 30045
rect 18515 30036 18527 30039
rect 17788 30008 18527 30036
rect 18515 30005 18527 30008
rect 18561 30036 18573 30039
rect 19150 30036 19156 30048
rect 18561 30008 19156 30036
rect 18561 30005 18573 30008
rect 18515 29999 18573 30005
rect 19150 29996 19156 30008
rect 19208 29996 19214 30048
rect 19904 30045 19932 30144
rect 20257 30141 20269 30175
rect 20303 30172 20315 30175
rect 20717 30175 20775 30181
rect 20717 30172 20729 30175
rect 20303 30144 20729 30172
rect 20303 30141 20315 30144
rect 20257 30135 20315 30141
rect 20717 30141 20729 30144
rect 20763 30172 20775 30175
rect 20806 30172 20812 30184
rect 20763 30144 20812 30172
rect 20763 30141 20775 30144
rect 20717 30135 20775 30141
rect 20806 30132 20812 30144
rect 20864 30132 20870 30184
rect 23658 30172 23664 30184
rect 23619 30144 23664 30172
rect 23658 30132 23664 30144
rect 23716 30172 23722 30184
rect 24213 30175 24271 30181
rect 24213 30172 24225 30175
rect 23716 30144 24225 30172
rect 23716 30132 23722 30144
rect 24213 30141 24225 30144
rect 24259 30172 24271 30175
rect 24394 30172 24400 30184
rect 24259 30144 24400 30172
rect 24259 30141 24271 30144
rect 24213 30135 24271 30141
rect 24394 30132 24400 30144
rect 24452 30132 24458 30184
rect 24765 30175 24823 30181
rect 24765 30141 24777 30175
rect 24811 30141 24823 30175
rect 24872 30172 24900 30212
rect 33042 30200 33048 30212
rect 33100 30200 33106 30252
rect 25021 30175 25079 30181
rect 25021 30172 25033 30175
rect 24872 30144 25033 30172
rect 24765 30135 24823 30141
rect 25021 30141 25033 30144
rect 25067 30141 25079 30175
rect 26970 30172 26976 30184
rect 26931 30144 26976 30172
rect 25021 30135 25079 30141
rect 20962 30107 21020 30113
rect 20962 30104 20974 30107
rect 20548 30076 20974 30104
rect 20548 30048 20576 30076
rect 20962 30073 20974 30076
rect 21008 30073 21020 30107
rect 20962 30067 21020 30073
rect 23477 30107 23535 30113
rect 23477 30073 23489 30107
rect 23523 30104 23535 30107
rect 24026 30104 24032 30116
rect 23523 30076 24032 30104
rect 23523 30073 23535 30076
rect 23477 30067 23535 30073
rect 24026 30064 24032 30076
rect 24084 30104 24090 30116
rect 24780 30104 24808 30135
rect 26970 30132 26976 30144
rect 27028 30172 27034 30184
rect 27525 30175 27583 30181
rect 27525 30172 27537 30175
rect 27028 30144 27537 30172
rect 27028 30132 27034 30144
rect 27525 30141 27537 30144
rect 27571 30141 27583 30175
rect 27525 30135 27583 30141
rect 35437 30175 35495 30181
rect 35437 30141 35449 30175
rect 35483 30172 35495 30175
rect 35710 30172 35716 30184
rect 35483 30144 35716 30172
rect 35483 30141 35495 30144
rect 35437 30135 35495 30141
rect 35710 30132 35716 30144
rect 35768 30172 35774 30184
rect 35989 30175 36047 30181
rect 35989 30172 36001 30175
rect 35768 30144 36001 30172
rect 35768 30132 35774 30144
rect 35989 30141 36001 30144
rect 36035 30141 36047 30175
rect 35989 30135 36047 30141
rect 32861 30107 32919 30113
rect 32861 30104 32873 30107
rect 24084 30076 24808 30104
rect 32232 30076 32873 30104
rect 24084 30064 24090 30076
rect 32232 30048 32260 30076
rect 32861 30073 32873 30076
rect 32907 30073 32919 30107
rect 32861 30067 32919 30073
rect 19889 30039 19947 30045
rect 19889 30005 19901 30039
rect 19935 30036 19947 30039
rect 20070 30036 20076 30048
rect 19935 30008 20076 30036
rect 19935 30005 19947 30008
rect 19889 29999 19947 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 20530 30036 20536 30048
rect 20491 30008 20536 30036
rect 20530 29996 20536 30008
rect 20588 29996 20594 30048
rect 23842 30036 23848 30048
rect 23803 30008 23848 30036
rect 23842 29996 23848 30008
rect 23900 29996 23906 30048
rect 26142 30036 26148 30048
rect 26103 30008 26148 30036
rect 26142 29996 26148 30008
rect 26200 29996 26206 30048
rect 27154 30036 27160 30048
rect 27115 30008 27160 30036
rect 27154 29996 27160 30008
rect 27212 29996 27218 30048
rect 32214 30036 32220 30048
rect 32175 30008 32220 30036
rect 32214 29996 32220 30008
rect 32272 29996 32278 30048
rect 32401 30039 32459 30045
rect 32401 30005 32413 30039
rect 32447 30036 32459 30039
rect 32490 30036 32496 30048
rect 32447 30008 32496 30036
rect 32447 30005 32459 30008
rect 32401 29999 32459 30005
rect 32490 29996 32496 30008
rect 32548 29996 32554 30048
rect 32766 30036 32772 30048
rect 32727 30008 32772 30036
rect 32766 29996 32772 30008
rect 32824 29996 32830 30048
rect 35345 30039 35403 30045
rect 35345 30005 35357 30039
rect 35391 30036 35403 30039
rect 35618 30036 35624 30048
rect 35391 30008 35624 30036
rect 35391 30005 35403 30008
rect 35345 29999 35403 30005
rect 35618 29996 35624 30008
rect 35676 29996 35682 30048
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 2314 29832 2320 29844
rect 2275 29804 2320 29832
rect 2314 29792 2320 29804
rect 2372 29792 2378 29844
rect 2409 29835 2467 29841
rect 2409 29801 2421 29835
rect 2455 29832 2467 29835
rect 2682 29832 2688 29844
rect 2455 29804 2688 29832
rect 2455 29801 2467 29804
rect 2409 29795 2467 29801
rect 2682 29792 2688 29804
rect 2740 29792 2746 29844
rect 5994 29832 6000 29844
rect 5955 29804 6000 29832
rect 5994 29792 6000 29804
rect 6052 29792 6058 29844
rect 6270 29792 6276 29844
rect 6328 29832 6334 29844
rect 7837 29835 7895 29841
rect 7837 29832 7849 29835
rect 6328 29804 7849 29832
rect 6328 29792 6334 29804
rect 7837 29801 7849 29804
rect 7883 29801 7895 29835
rect 7837 29795 7895 29801
rect 8570 29792 8576 29844
rect 8628 29832 8634 29844
rect 8849 29835 8907 29841
rect 8849 29832 8861 29835
rect 8628 29804 8861 29832
rect 8628 29792 8634 29804
rect 8849 29801 8861 29804
rect 8895 29801 8907 29835
rect 8849 29795 8907 29801
rect 10686 29792 10692 29844
rect 10744 29832 10750 29844
rect 11057 29835 11115 29841
rect 11057 29832 11069 29835
rect 10744 29804 11069 29832
rect 10744 29792 10750 29804
rect 11057 29801 11069 29804
rect 11103 29801 11115 29835
rect 11422 29832 11428 29844
rect 11383 29804 11428 29832
rect 11057 29795 11115 29801
rect 11422 29792 11428 29804
rect 11480 29792 11486 29844
rect 14185 29835 14243 29841
rect 14185 29801 14197 29835
rect 14231 29832 14243 29835
rect 14274 29832 14280 29844
rect 14231 29804 14280 29832
rect 14231 29801 14243 29804
rect 14185 29795 14243 29801
rect 14274 29792 14280 29804
rect 14332 29792 14338 29844
rect 15654 29792 15660 29844
rect 15712 29832 15718 29844
rect 16123 29835 16181 29841
rect 16123 29832 16135 29835
rect 15712 29804 16135 29832
rect 15712 29792 15718 29804
rect 16123 29801 16135 29804
rect 16169 29801 16181 29835
rect 17494 29832 17500 29844
rect 17407 29804 17500 29832
rect 16123 29795 16181 29801
rect 17494 29792 17500 29804
rect 17552 29832 17558 29844
rect 18509 29835 18567 29841
rect 18509 29832 18521 29835
rect 17552 29804 18521 29832
rect 17552 29792 17558 29804
rect 18509 29801 18521 29804
rect 18555 29832 18567 29835
rect 18782 29832 18788 29844
rect 18555 29804 18788 29832
rect 18555 29801 18567 29804
rect 18509 29795 18567 29801
rect 18782 29792 18788 29804
rect 18840 29792 18846 29844
rect 20530 29792 20536 29844
rect 20588 29832 20594 29844
rect 22281 29835 22339 29841
rect 22281 29832 22293 29835
rect 20588 29804 22293 29832
rect 20588 29792 20594 29804
rect 22281 29801 22293 29804
rect 22327 29801 22339 29835
rect 22281 29795 22339 29801
rect 23842 29792 23848 29844
rect 23900 29832 23906 29844
rect 24578 29832 24584 29844
rect 23900 29804 24584 29832
rect 23900 29792 23906 29804
rect 24578 29792 24584 29804
rect 24636 29832 24642 29844
rect 24949 29835 25007 29841
rect 24949 29832 24961 29835
rect 24636 29804 24961 29832
rect 24636 29792 24642 29804
rect 24949 29801 24961 29804
rect 24995 29801 25007 29835
rect 24949 29795 25007 29801
rect 25041 29835 25099 29841
rect 25041 29801 25053 29835
rect 25087 29832 25099 29835
rect 27154 29832 27160 29844
rect 25087 29804 27160 29832
rect 25087 29801 25099 29804
rect 25041 29795 25099 29801
rect 2332 29764 2360 29792
rect 2332 29736 3004 29764
rect 2774 29656 2780 29708
rect 2832 29696 2838 29708
rect 2832 29668 2877 29696
rect 2832 29656 2838 29668
rect 2498 29588 2504 29640
rect 2556 29628 2562 29640
rect 2976 29637 3004 29736
rect 3050 29724 3056 29776
rect 3108 29764 3114 29776
rect 4494 29767 4552 29773
rect 4494 29764 4506 29767
rect 3108 29736 4506 29764
rect 3108 29724 3114 29736
rect 4494 29733 4506 29736
rect 4540 29764 4552 29767
rect 4614 29764 4620 29776
rect 4540 29736 4620 29764
rect 4540 29733 4552 29736
rect 4494 29727 4552 29733
rect 4614 29724 4620 29736
rect 4672 29724 4678 29776
rect 9858 29724 9864 29776
rect 9916 29773 9922 29776
rect 9916 29767 9980 29773
rect 9916 29733 9934 29767
rect 9968 29733 9980 29767
rect 9916 29727 9980 29733
rect 9916 29724 9922 29727
rect 12894 29724 12900 29776
rect 12952 29764 12958 29776
rect 13050 29767 13108 29773
rect 13050 29764 13062 29767
rect 12952 29736 13062 29764
rect 12952 29724 12958 29736
rect 13050 29733 13062 29736
rect 13096 29733 13108 29767
rect 18138 29764 18144 29776
rect 18099 29736 18144 29764
rect 13050 29727 13108 29733
rect 18138 29724 18144 29736
rect 18196 29724 18202 29776
rect 24118 29764 24124 29776
rect 24079 29736 24124 29764
rect 24118 29724 24124 29736
rect 24176 29724 24182 29776
rect 24394 29764 24400 29776
rect 24355 29736 24400 29764
rect 24394 29724 24400 29736
rect 24452 29724 24458 29776
rect 24486 29724 24492 29776
rect 24544 29764 24550 29776
rect 25056 29764 25084 29795
rect 27154 29792 27160 29804
rect 27212 29792 27218 29844
rect 35894 29832 35900 29844
rect 35855 29804 35900 29832
rect 35894 29792 35900 29804
rect 35952 29792 35958 29844
rect 24544 29736 25084 29764
rect 24544 29724 24550 29736
rect 3878 29696 3884 29708
rect 3791 29668 3884 29696
rect 3878 29656 3884 29668
rect 3936 29696 3942 29708
rect 4249 29699 4307 29705
rect 4249 29696 4261 29699
rect 3936 29668 4261 29696
rect 3936 29656 3942 29668
rect 4249 29665 4261 29668
rect 4295 29696 4307 29699
rect 5350 29696 5356 29708
rect 4295 29668 5356 29696
rect 4295 29665 4307 29668
rect 4249 29659 4307 29665
rect 5350 29656 5356 29668
rect 5408 29656 5414 29708
rect 6546 29696 6552 29708
rect 5644 29668 6552 29696
rect 2869 29631 2927 29637
rect 2869 29628 2881 29631
rect 2556 29600 2881 29628
rect 2556 29588 2562 29600
rect 2869 29597 2881 29600
rect 2915 29597 2927 29631
rect 2869 29591 2927 29597
rect 2961 29631 3019 29637
rect 2961 29597 2973 29631
rect 3007 29597 3019 29631
rect 2961 29591 3019 29597
rect 5644 29572 5672 29668
rect 6546 29656 6552 29668
rect 6604 29696 6610 29708
rect 6713 29699 6771 29705
rect 6713 29696 6725 29699
rect 6604 29668 6725 29696
rect 6604 29656 6610 29668
rect 6713 29665 6725 29668
rect 6759 29665 6771 29699
rect 6713 29659 6771 29665
rect 8573 29699 8631 29705
rect 8573 29665 8585 29699
rect 8619 29696 8631 29699
rect 8662 29696 8668 29708
rect 8619 29668 8668 29696
rect 8619 29665 8631 29668
rect 8573 29659 8631 29665
rect 8662 29656 8668 29668
rect 8720 29656 8726 29708
rect 9677 29699 9735 29705
rect 9677 29665 9689 29699
rect 9723 29696 9735 29699
rect 9766 29696 9772 29708
rect 9723 29668 9772 29696
rect 9723 29665 9735 29668
rect 9677 29659 9735 29665
rect 6365 29631 6423 29637
rect 6365 29597 6377 29631
rect 6411 29628 6423 29631
rect 6454 29628 6460 29640
rect 6411 29600 6460 29628
rect 6411 29597 6423 29600
rect 6365 29591 6423 29597
rect 6454 29588 6460 29600
rect 6512 29588 6518 29640
rect 7742 29588 7748 29640
rect 7800 29628 7806 29640
rect 8205 29631 8263 29637
rect 8205 29628 8217 29631
rect 7800 29600 8217 29628
rect 7800 29588 7806 29600
rect 8205 29597 8217 29600
rect 8251 29628 8263 29631
rect 8478 29628 8484 29640
rect 8251 29600 8484 29628
rect 8251 29597 8263 29600
rect 8205 29591 8263 29597
rect 8478 29588 8484 29600
rect 8536 29628 8542 29640
rect 9692 29628 9720 29659
rect 9766 29656 9772 29668
rect 9824 29656 9830 29708
rect 14182 29656 14188 29708
rect 14240 29696 14246 29708
rect 14829 29699 14887 29705
rect 14829 29696 14841 29699
rect 14240 29668 14841 29696
rect 14240 29656 14246 29668
rect 14829 29665 14841 29668
rect 14875 29696 14887 29699
rect 15010 29696 15016 29708
rect 14875 29668 15016 29696
rect 14875 29665 14887 29668
rect 14829 29659 14887 29665
rect 15010 29656 15016 29668
rect 15068 29656 15074 29708
rect 15378 29656 15384 29708
rect 15436 29696 15442 29708
rect 16393 29699 16451 29705
rect 16393 29696 16405 29699
rect 15436 29668 16405 29696
rect 15436 29656 15442 29668
rect 16393 29665 16405 29668
rect 16439 29696 16451 29699
rect 16758 29696 16764 29708
rect 16439 29668 16764 29696
rect 16439 29665 16451 29668
rect 16393 29659 16451 29665
rect 16758 29656 16764 29668
rect 16816 29656 16822 29708
rect 19610 29696 19616 29708
rect 19571 29668 19616 29696
rect 19610 29656 19616 29668
rect 19668 29656 19674 29708
rect 20806 29656 20812 29708
rect 20864 29696 20870 29708
rect 21174 29705 21180 29708
rect 20901 29699 20959 29705
rect 20901 29696 20913 29699
rect 20864 29668 20913 29696
rect 20864 29656 20870 29668
rect 20901 29665 20913 29668
rect 20947 29665 20959 29699
rect 21168 29696 21180 29705
rect 21135 29668 21180 29696
rect 20901 29659 20959 29665
rect 21168 29659 21180 29668
rect 21174 29656 21180 29659
rect 21232 29656 21238 29708
rect 32493 29699 32551 29705
rect 32493 29665 32505 29699
rect 32539 29696 32551 29699
rect 32766 29696 32772 29708
rect 32539 29668 32772 29696
rect 32539 29665 32551 29668
rect 32493 29659 32551 29665
rect 32766 29656 32772 29668
rect 32824 29696 32830 29708
rect 33594 29696 33600 29708
rect 32824 29668 33600 29696
rect 32824 29656 32830 29668
rect 33594 29656 33600 29668
rect 33652 29696 33658 29708
rect 33761 29699 33819 29705
rect 33761 29696 33773 29699
rect 33652 29668 33773 29696
rect 33652 29656 33658 29668
rect 33761 29665 33773 29668
rect 33807 29665 33819 29699
rect 33761 29659 33819 29665
rect 34514 29656 34520 29708
rect 34572 29696 34578 29708
rect 35526 29696 35532 29708
rect 34572 29668 35532 29696
rect 34572 29656 34578 29668
rect 35526 29656 35532 29668
rect 35584 29656 35590 29708
rect 35713 29699 35771 29705
rect 35713 29665 35725 29699
rect 35759 29696 35771 29699
rect 35802 29696 35808 29708
rect 35759 29668 35808 29696
rect 35759 29665 35771 29668
rect 35713 29659 35771 29665
rect 35802 29656 35808 29668
rect 35860 29656 35866 29708
rect 8536 29600 9720 29628
rect 8536 29588 8542 29600
rect 11054 29588 11060 29640
rect 11112 29628 11118 29640
rect 12161 29631 12219 29637
rect 12161 29628 12173 29631
rect 11112 29600 12173 29628
rect 11112 29588 11118 29600
rect 12161 29597 12173 29600
rect 12207 29628 12219 29631
rect 12805 29631 12863 29637
rect 12805 29628 12817 29631
rect 12207 29600 12817 29628
rect 12207 29597 12219 29600
rect 12161 29591 12219 29597
rect 12805 29597 12817 29600
rect 12851 29597 12863 29631
rect 12805 29591 12863 29597
rect 15470 29588 15476 29640
rect 15528 29628 15534 29640
rect 15565 29631 15623 29637
rect 15565 29628 15577 29631
rect 15528 29600 15577 29628
rect 15528 29588 15534 29600
rect 15565 29597 15577 29600
rect 15611 29628 15623 29631
rect 15657 29631 15715 29637
rect 15657 29628 15669 29631
rect 15611 29600 15669 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 15657 29597 15669 29600
rect 15703 29628 15715 29631
rect 15838 29628 15844 29640
rect 15703 29600 15844 29628
rect 15703 29597 15715 29600
rect 15657 29591 15715 29597
rect 15838 29588 15844 29600
rect 15896 29588 15902 29640
rect 16163 29631 16221 29637
rect 16163 29597 16175 29631
rect 16209 29628 16221 29631
rect 16298 29628 16304 29640
rect 16209 29600 16304 29628
rect 16209 29597 16221 29600
rect 16163 29591 16221 29597
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 19705 29631 19763 29637
rect 19705 29628 19717 29631
rect 19392 29600 19717 29628
rect 19392 29588 19398 29600
rect 19705 29597 19717 29600
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 19797 29631 19855 29637
rect 19797 29597 19809 29631
rect 19843 29628 19855 29631
rect 20530 29628 20536 29640
rect 19843 29600 20536 29628
rect 19843 29597 19855 29600
rect 19797 29591 19855 29597
rect 5626 29560 5632 29572
rect 5539 29532 5632 29560
rect 5626 29520 5632 29532
rect 5684 29520 5690 29572
rect 19058 29520 19064 29572
rect 19116 29560 19122 29572
rect 19812 29560 19840 29591
rect 20530 29588 20536 29600
rect 20588 29588 20594 29640
rect 25130 29588 25136 29640
rect 25188 29628 25194 29640
rect 25593 29631 25651 29637
rect 25593 29628 25605 29631
rect 25188 29600 25605 29628
rect 25188 29588 25194 29600
rect 25593 29597 25605 29600
rect 25639 29628 25651 29631
rect 26142 29628 26148 29640
rect 25639 29600 26148 29628
rect 25639 29597 25651 29600
rect 25593 29591 25651 29597
rect 26142 29588 26148 29600
rect 26200 29588 26206 29640
rect 26513 29631 26571 29637
rect 26513 29597 26525 29631
rect 26559 29628 26571 29631
rect 26786 29628 26792 29640
rect 26559 29600 26792 29628
rect 26559 29597 26571 29600
rect 26513 29591 26571 29597
rect 26786 29588 26792 29600
rect 26844 29588 26850 29640
rect 33502 29628 33508 29640
rect 33463 29600 33508 29628
rect 33502 29588 33508 29600
rect 33560 29588 33566 29640
rect 19116 29532 19840 29560
rect 19116 29520 19122 29532
rect 12529 29495 12587 29501
rect 12529 29461 12541 29495
rect 12575 29492 12587 29495
rect 12710 29492 12716 29504
rect 12575 29464 12716 29492
rect 12575 29461 12587 29464
rect 12529 29455 12587 29461
rect 12710 29452 12716 29464
rect 12768 29452 12774 29504
rect 13998 29452 14004 29504
rect 14056 29492 14062 29504
rect 14461 29495 14519 29501
rect 14461 29492 14473 29495
rect 14056 29464 14473 29492
rect 14056 29452 14062 29464
rect 14461 29461 14473 29464
rect 14507 29492 14519 29495
rect 14550 29492 14556 29504
rect 14507 29464 14556 29492
rect 14507 29461 14519 29464
rect 14461 29455 14519 29461
rect 14550 29452 14556 29464
rect 14608 29452 14614 29504
rect 19153 29495 19211 29501
rect 19153 29461 19165 29495
rect 19199 29492 19211 29495
rect 19242 29492 19248 29504
rect 19199 29464 19248 29492
rect 19199 29461 19211 29464
rect 19153 29455 19211 29461
rect 19242 29452 19248 29464
rect 19300 29452 19306 29504
rect 24581 29495 24639 29501
rect 24581 29461 24593 29495
rect 24627 29492 24639 29495
rect 24762 29492 24768 29504
rect 24627 29464 24768 29492
rect 24627 29461 24639 29464
rect 24581 29455 24639 29461
rect 24762 29452 24768 29464
rect 24820 29452 24826 29504
rect 26142 29452 26148 29504
rect 26200 29492 26206 29504
rect 27062 29492 27068 29504
rect 26200 29464 27068 29492
rect 26200 29452 26206 29464
rect 27062 29452 27068 29464
rect 27120 29452 27126 29504
rect 34698 29452 34704 29504
rect 34756 29492 34762 29504
rect 34885 29495 34943 29501
rect 34885 29492 34897 29495
rect 34756 29464 34897 29492
rect 34756 29452 34762 29464
rect 34885 29461 34897 29464
rect 34931 29461 34943 29495
rect 34885 29455 34943 29461
rect 35253 29495 35311 29501
rect 35253 29461 35265 29495
rect 35299 29492 35311 29495
rect 35894 29492 35900 29504
rect 35299 29464 35900 29492
rect 35299 29461 35311 29464
rect 35253 29455 35311 29461
rect 35894 29452 35900 29464
rect 35952 29452 35958 29504
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 2498 29288 2504 29300
rect 2459 29260 2504 29288
rect 2498 29248 2504 29260
rect 2556 29248 2562 29300
rect 4062 29288 4068 29300
rect 4023 29260 4068 29288
rect 4062 29248 4068 29260
rect 4120 29248 4126 29300
rect 4433 29291 4491 29297
rect 4433 29257 4445 29291
rect 4479 29288 4491 29291
rect 4614 29288 4620 29300
rect 4479 29260 4620 29288
rect 4479 29257 4491 29260
rect 4433 29251 4491 29257
rect 4614 29248 4620 29260
rect 4672 29248 4678 29300
rect 5074 29248 5080 29300
rect 5132 29288 5138 29300
rect 5169 29291 5227 29297
rect 5169 29288 5181 29291
rect 5132 29260 5181 29288
rect 5132 29248 5138 29260
rect 5169 29257 5181 29260
rect 5215 29257 5227 29291
rect 6546 29288 6552 29300
rect 6507 29260 6552 29288
rect 5169 29251 5227 29257
rect 6546 29248 6552 29260
rect 6604 29248 6610 29300
rect 9950 29288 9956 29300
rect 9911 29260 9956 29288
rect 9950 29248 9956 29260
rect 10008 29248 10014 29300
rect 11330 29288 11336 29300
rect 11291 29260 11336 29288
rect 11330 29248 11336 29260
rect 11388 29248 11394 29300
rect 11422 29248 11428 29300
rect 11480 29288 11486 29300
rect 11793 29291 11851 29297
rect 11793 29288 11805 29291
rect 11480 29260 11805 29288
rect 11480 29248 11486 29260
rect 11793 29257 11805 29260
rect 11839 29257 11851 29291
rect 11793 29251 11851 29257
rect 9769 29223 9827 29229
rect 9769 29189 9781 29223
rect 9815 29220 9827 29223
rect 9858 29220 9864 29232
rect 9815 29192 9864 29220
rect 9815 29189 9827 29192
rect 9769 29183 9827 29189
rect 9858 29180 9864 29192
rect 9916 29180 9922 29232
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29152 5135 29155
rect 5626 29152 5632 29164
rect 5123 29124 5632 29152
rect 5123 29121 5135 29124
rect 5077 29115 5135 29121
rect 5626 29112 5632 29124
rect 5684 29112 5690 29164
rect 5721 29155 5779 29161
rect 5721 29121 5733 29155
rect 5767 29152 5779 29155
rect 5994 29152 6000 29164
rect 5767 29124 6000 29152
rect 5767 29121 5779 29124
rect 5721 29115 5779 29121
rect 5994 29112 6000 29124
rect 6052 29112 6058 29164
rect 6454 29112 6460 29164
rect 6512 29152 6518 29164
rect 7101 29155 7159 29161
rect 7101 29152 7113 29155
rect 6512 29124 7113 29152
rect 6512 29112 6518 29124
rect 7101 29121 7113 29124
rect 7147 29152 7159 29155
rect 7742 29152 7748 29164
rect 7147 29124 7748 29152
rect 7147 29121 7159 29124
rect 7101 29115 7159 29121
rect 7742 29112 7748 29124
rect 7800 29112 7806 29164
rect 10594 29152 10600 29164
rect 10507 29124 10600 29152
rect 10594 29112 10600 29124
rect 10652 29152 10658 29164
rect 11348 29152 11376 29248
rect 10652 29124 11376 29152
rect 11808 29152 11836 29251
rect 12894 29248 12900 29300
rect 12952 29288 12958 29300
rect 13449 29291 13507 29297
rect 13449 29288 13461 29291
rect 12952 29260 13461 29288
rect 12952 29248 12958 29260
rect 13449 29257 13461 29260
rect 13495 29257 13507 29291
rect 13449 29251 13507 29257
rect 15565 29291 15623 29297
rect 15565 29257 15577 29291
rect 15611 29288 15623 29291
rect 15654 29288 15660 29300
rect 15611 29260 15660 29288
rect 15611 29257 15623 29260
rect 15565 29251 15623 29257
rect 15654 29248 15660 29260
rect 15712 29248 15718 29300
rect 16574 29248 16580 29300
rect 16632 29288 16638 29300
rect 17037 29291 17095 29297
rect 17037 29288 17049 29291
rect 16632 29260 17049 29288
rect 16632 29248 16638 29260
rect 17037 29257 17049 29260
rect 17083 29257 17095 29291
rect 17310 29288 17316 29300
rect 17271 29260 17316 29288
rect 17037 29251 17095 29257
rect 17310 29248 17316 29260
rect 17368 29248 17374 29300
rect 17770 29288 17776 29300
rect 17731 29260 17776 29288
rect 17770 29248 17776 29260
rect 17828 29248 17834 29300
rect 18414 29288 18420 29300
rect 18375 29260 18420 29288
rect 18414 29248 18420 29260
rect 18472 29248 18478 29300
rect 18877 29291 18935 29297
rect 18877 29257 18889 29291
rect 18923 29288 18935 29291
rect 19610 29288 19616 29300
rect 18923 29260 19616 29288
rect 18923 29257 18935 29260
rect 18877 29251 18935 29257
rect 19610 29248 19616 29260
rect 19668 29248 19674 29300
rect 20806 29248 20812 29300
rect 20864 29288 20870 29300
rect 21818 29288 21824 29300
rect 20864 29260 21824 29288
rect 20864 29248 20870 29260
rect 21818 29248 21824 29260
rect 21876 29248 21882 29300
rect 24578 29288 24584 29300
rect 24539 29260 24584 29288
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 26142 29288 26148 29300
rect 26103 29260 26148 29288
rect 26142 29248 26148 29260
rect 26200 29248 26206 29300
rect 26418 29288 26424 29300
rect 26379 29260 26424 29288
rect 26418 29248 26424 29260
rect 26476 29248 26482 29300
rect 26786 29288 26792 29300
rect 26747 29260 26792 29288
rect 26786 29248 26792 29260
rect 26844 29248 26850 29300
rect 12434 29180 12440 29232
rect 12492 29220 12498 29232
rect 14001 29223 14059 29229
rect 12492 29192 12537 29220
rect 12492 29180 12498 29192
rect 14001 29189 14013 29223
rect 14047 29220 14059 29223
rect 15194 29220 15200 29232
rect 14047 29192 15200 29220
rect 14047 29189 14059 29192
rect 14001 29183 14059 29189
rect 15194 29180 15200 29192
rect 15252 29180 15258 29232
rect 19150 29220 19156 29232
rect 19111 29192 19156 29220
rect 19150 29180 19156 29192
rect 19208 29180 19214 29232
rect 21177 29223 21235 29229
rect 21177 29189 21189 29223
rect 21223 29220 21235 29223
rect 21542 29220 21548 29232
rect 21223 29192 21548 29220
rect 21223 29189 21235 29192
rect 21177 29183 21235 29189
rect 21542 29180 21548 29192
rect 21600 29180 21606 29232
rect 23845 29223 23903 29229
rect 23845 29189 23857 29223
rect 23891 29220 23903 29223
rect 24210 29220 24216 29232
rect 23891 29192 24216 29220
rect 23891 29189 23903 29192
rect 23845 29183 23903 29189
rect 24210 29180 24216 29192
rect 24268 29180 24274 29232
rect 24305 29223 24363 29229
rect 24305 29189 24317 29223
rect 24351 29220 24363 29223
rect 24486 29220 24492 29232
rect 24351 29192 24492 29220
rect 24351 29189 24363 29192
rect 24305 29183 24363 29189
rect 24486 29180 24492 29192
rect 24544 29180 24550 29232
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 11808 29124 13093 29152
rect 10652 29112 10658 29124
rect 13081 29121 13093 29124
rect 13127 29152 13139 29155
rect 13722 29152 13728 29164
rect 13127 29124 13728 29152
rect 13127 29121 13139 29124
rect 13081 29115 13139 29121
rect 13722 29112 13728 29124
rect 13780 29112 13786 29164
rect 14274 29112 14280 29164
rect 14332 29152 14338 29164
rect 14553 29155 14611 29161
rect 14553 29152 14565 29155
rect 14332 29124 14565 29152
rect 14332 29112 14338 29124
rect 14553 29121 14565 29124
rect 14599 29121 14611 29155
rect 14553 29115 14611 29121
rect 15010 29112 15016 29164
rect 15068 29152 15074 29164
rect 15657 29155 15715 29161
rect 15657 29152 15669 29155
rect 15068 29124 15669 29152
rect 15068 29112 15074 29124
rect 15657 29121 15669 29124
rect 15703 29121 15715 29155
rect 15657 29115 15715 29121
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 19800 29155 19858 29161
rect 19800 29152 19812 29155
rect 19300 29124 19812 29152
rect 19300 29112 19306 29124
rect 19800 29121 19812 29124
rect 19846 29121 19858 29155
rect 20070 29152 20076 29164
rect 20031 29124 20076 29152
rect 19800 29115 19858 29121
rect 20070 29112 20076 29124
rect 20128 29112 20134 29164
rect 2038 29044 2044 29096
rect 2096 29084 2102 29096
rect 2685 29087 2743 29093
rect 2685 29084 2697 29087
rect 2096 29056 2697 29084
rect 2096 29044 2102 29056
rect 2685 29053 2697 29056
rect 2731 29053 2743 29087
rect 2685 29047 2743 29053
rect 5537 29087 5595 29093
rect 5537 29053 5549 29087
rect 5583 29084 5595 29087
rect 5810 29084 5816 29096
rect 5583 29056 5816 29084
rect 5583 29053 5595 29056
rect 5537 29047 5595 29053
rect 5810 29044 5816 29056
rect 5868 29084 5874 29096
rect 6270 29084 6276 29096
rect 5868 29056 6276 29084
rect 5868 29044 5874 29056
rect 6270 29044 6276 29056
rect 6328 29044 6334 29096
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 10321 29087 10379 29093
rect 10321 29084 10333 29087
rect 9732 29056 10333 29084
rect 9732 29044 9738 29056
rect 10321 29053 10333 29056
rect 10367 29084 10379 29087
rect 10965 29087 11023 29093
rect 10965 29084 10977 29087
rect 10367 29056 10977 29084
rect 10367 29053 10379 29056
rect 10321 29047 10379 29053
rect 10965 29053 10977 29056
rect 11011 29053 11023 29087
rect 10965 29047 11023 29053
rect 12710 29044 12716 29096
rect 12768 29084 12774 29096
rect 12805 29087 12863 29093
rect 12805 29084 12817 29087
rect 12768 29056 12817 29084
rect 12768 29044 12774 29056
rect 12805 29053 12817 29056
rect 12851 29053 12863 29087
rect 12805 29047 12863 29053
rect 15197 29087 15255 29093
rect 15197 29053 15209 29087
rect 15243 29084 15255 29087
rect 15378 29084 15384 29096
rect 15243 29056 15384 29084
rect 15243 29053 15255 29056
rect 15197 29047 15255 29053
rect 15378 29044 15384 29056
rect 15436 29044 15442 29096
rect 15924 29087 15982 29093
rect 15924 29053 15936 29087
rect 15970 29084 15982 29087
rect 17310 29084 17316 29096
rect 15970 29056 17316 29084
rect 15970 29053 15982 29056
rect 15924 29047 15982 29053
rect 17310 29044 17316 29056
rect 17368 29044 17374 29096
rect 18874 29044 18880 29096
rect 18932 29084 18938 29096
rect 19337 29087 19395 29093
rect 19337 29084 19349 29087
rect 18932 29056 19349 29084
rect 18932 29044 18938 29056
rect 19337 29053 19349 29056
rect 19383 29084 19395 29087
rect 20346 29084 20352 29096
rect 19383 29056 20352 29084
rect 19383 29053 19395 29056
rect 19337 29047 19395 29053
rect 20346 29044 20352 29056
rect 20404 29044 20410 29096
rect 20714 29044 20720 29096
rect 20772 29084 20778 29096
rect 21174 29084 21180 29096
rect 20772 29056 21180 29084
rect 20772 29044 20778 29056
rect 21174 29044 21180 29056
rect 21232 29084 21238 29096
rect 21453 29087 21511 29093
rect 21453 29084 21465 29087
rect 21232 29056 21465 29084
rect 21232 29044 21238 29056
rect 21453 29053 21465 29056
rect 21499 29084 21511 29087
rect 21910 29084 21916 29096
rect 21499 29056 21916 29084
rect 21499 29053 21511 29056
rect 21453 29047 21511 29053
rect 21910 29044 21916 29056
rect 21968 29044 21974 29096
rect 23477 29087 23535 29093
rect 23477 29053 23489 29087
rect 23523 29084 23535 29087
rect 23661 29087 23719 29093
rect 23661 29084 23673 29087
rect 23523 29056 23673 29084
rect 23523 29053 23535 29056
rect 23477 29047 23535 29053
rect 23661 29053 23673 29056
rect 23707 29084 23719 29087
rect 23934 29084 23940 29096
rect 23707 29056 23940 29084
rect 23707 29053 23719 29056
rect 23661 29047 23719 29053
rect 23934 29044 23940 29056
rect 23992 29044 23998 29096
rect 24026 29044 24032 29096
rect 24084 29084 24090 29096
rect 24765 29087 24823 29093
rect 24765 29084 24777 29087
rect 24084 29056 24777 29084
rect 24084 29044 24090 29056
rect 24765 29053 24777 29056
rect 24811 29084 24823 29087
rect 26804 29084 26832 29248
rect 26878 29180 26884 29232
rect 26936 29220 26942 29232
rect 26973 29223 27031 29229
rect 26973 29220 26985 29223
rect 26936 29192 26985 29220
rect 26936 29180 26942 29192
rect 26973 29189 26985 29192
rect 27019 29189 27031 29223
rect 26973 29183 27031 29189
rect 34790 29180 34796 29232
rect 34848 29220 34854 29232
rect 34885 29223 34943 29229
rect 34885 29220 34897 29223
rect 34848 29192 34897 29220
rect 34848 29180 34854 29192
rect 34885 29189 34897 29192
rect 34931 29189 34943 29223
rect 34885 29183 34943 29189
rect 34974 29180 34980 29232
rect 35032 29220 35038 29232
rect 35710 29220 35716 29232
rect 35032 29192 35716 29220
rect 35032 29180 35038 29192
rect 35710 29180 35716 29192
rect 35768 29180 35774 29232
rect 27062 29112 27068 29164
rect 27120 29152 27126 29164
rect 27525 29155 27583 29161
rect 27525 29152 27537 29155
rect 27120 29124 27537 29152
rect 27120 29112 27126 29124
rect 27525 29121 27537 29124
rect 27571 29121 27583 29155
rect 27525 29115 27583 29121
rect 35529 29155 35587 29161
rect 35529 29121 35541 29155
rect 35575 29152 35587 29155
rect 35894 29152 35900 29164
rect 35575 29124 35900 29152
rect 35575 29121 35587 29124
rect 35529 29115 35587 29121
rect 35894 29112 35900 29124
rect 35952 29112 35958 29164
rect 27341 29087 27399 29093
rect 27341 29084 27353 29087
rect 24811 29056 25268 29084
rect 26804 29056 27353 29084
rect 24811 29053 24823 29056
rect 24765 29047 24823 29053
rect 1765 29019 1823 29025
rect 1765 28985 1777 29019
rect 1811 29016 1823 29019
rect 2133 29019 2191 29025
rect 2133 29016 2145 29019
rect 1811 28988 2145 29016
rect 1811 28985 1823 28988
rect 1765 28979 1823 28985
rect 2133 28985 2145 28988
rect 2179 29016 2191 29019
rect 2774 29016 2780 29028
rect 2179 28988 2780 29016
rect 2179 28985 2191 28988
rect 2133 28979 2191 28985
rect 2774 28976 2780 28988
rect 2832 29016 2838 29028
rect 2930 29019 2988 29025
rect 2930 29016 2942 29019
rect 2832 28988 2942 29016
rect 2832 28976 2838 28988
rect 2930 28985 2942 28988
rect 2976 28985 2988 29019
rect 2930 28979 2988 28985
rect 7653 29019 7711 29025
rect 7653 28985 7665 29019
rect 7699 29016 7711 29019
rect 7990 29019 8048 29025
rect 7990 29016 8002 29019
rect 7699 28988 8002 29016
rect 7699 28985 7711 28988
rect 7653 28979 7711 28985
rect 7990 28985 8002 28988
rect 8036 29016 8048 29019
rect 8294 29016 8300 29028
rect 8036 28988 8300 29016
rect 8036 28985 8048 28988
rect 7990 28979 8048 28985
rect 8294 28976 8300 28988
rect 8352 28976 8358 29028
rect 12161 29019 12219 29025
rect 12161 29016 12173 29019
rect 10980 28988 12173 29016
rect 10980 28960 11008 28988
rect 12161 28985 12173 28988
rect 12207 29016 12219 29019
rect 12897 29019 12955 29025
rect 12897 29016 12909 29019
rect 12207 28988 12909 29016
rect 12207 28985 12219 28988
rect 12161 28979 12219 28985
rect 12897 28985 12909 28988
rect 12943 28985 12955 29019
rect 13814 29016 13820 29028
rect 13775 28988 13820 29016
rect 12897 28979 12955 28985
rect 13814 28976 13820 28988
rect 13872 29016 13878 29028
rect 14369 29019 14427 29025
rect 14369 29016 14381 29019
rect 13872 28988 14381 29016
rect 13872 28976 13878 28988
rect 14369 28985 14381 28988
rect 14415 28985 14427 29019
rect 14369 28979 14427 28985
rect 19150 28976 19156 29028
rect 19208 29016 19214 29028
rect 19208 28988 19380 29016
rect 19208 28976 19214 28988
rect 9122 28948 9128 28960
rect 9083 28920 9128 28948
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 10410 28908 10416 28960
rect 10468 28948 10474 28960
rect 10468 28920 10513 28948
rect 10468 28908 10474 28920
rect 10962 28908 10968 28960
rect 11020 28908 11026 28960
rect 14458 28908 14464 28960
rect 14516 28948 14522 28960
rect 19352 28948 19380 28988
rect 21266 28976 21272 29028
rect 21324 29016 21330 29028
rect 22005 29019 22063 29025
rect 22005 29016 22017 29019
rect 21324 28988 22017 29016
rect 21324 28976 21330 28988
rect 22005 28985 22017 28988
rect 22051 28985 22063 29019
rect 25010 29019 25068 29025
rect 25010 29016 25022 29019
rect 22005 28979 22063 28985
rect 24780 28988 25022 29016
rect 24780 28960 24808 28988
rect 25010 28985 25022 28988
rect 25056 29016 25068 29019
rect 25130 29016 25136 29028
rect 25056 28988 25136 29016
rect 25056 28985 25068 28988
rect 25010 28979 25068 28985
rect 25130 28976 25136 28988
rect 25188 28976 25194 29028
rect 19803 28951 19861 28957
rect 19803 28948 19815 28951
rect 14516 28920 14561 28948
rect 19352 28920 19815 28948
rect 14516 28908 14522 28920
rect 19803 28917 19815 28920
rect 19849 28948 19861 28951
rect 20530 28948 20536 28960
rect 19849 28920 20536 28948
rect 19849 28917 19861 28920
rect 19803 28911 19861 28917
rect 20530 28908 20536 28920
rect 20588 28908 20594 28960
rect 24762 28908 24768 28960
rect 24820 28908 24826 28960
rect 25240 28948 25268 29056
rect 27341 29053 27353 29056
rect 27387 29053 27399 29087
rect 31478 29084 31484 29096
rect 31439 29056 31484 29084
rect 27341 29047 27399 29053
rect 31478 29044 31484 29056
rect 31536 29044 31542 29096
rect 34333 29087 34391 29093
rect 34333 29053 34345 29087
rect 34379 29084 34391 29087
rect 35253 29087 35311 29093
rect 35253 29084 35265 29087
rect 34379 29056 35265 29084
rect 34379 29053 34391 29056
rect 34333 29047 34391 29053
rect 35253 29053 35265 29056
rect 35299 29084 35311 29087
rect 35710 29084 35716 29096
rect 35299 29056 35716 29084
rect 35299 29053 35311 29056
rect 35253 29047 35311 29053
rect 35710 29044 35716 29056
rect 35768 29044 35774 29096
rect 26418 28976 26424 29028
rect 26476 29016 26482 29028
rect 27433 29019 27491 29025
rect 27433 29016 27445 29019
rect 26476 28988 27445 29016
rect 26476 28976 26482 28988
rect 27433 28985 27445 28988
rect 27479 28985 27491 29019
rect 31726 29019 31784 29025
rect 31726 29016 31738 29019
rect 27433 28979 27491 28985
rect 31312 28988 31738 29016
rect 25498 28948 25504 28960
rect 25240 28920 25504 28948
rect 25498 28908 25504 28920
rect 25556 28908 25562 28960
rect 31202 28908 31208 28960
rect 31260 28948 31266 28960
rect 31312 28957 31340 28988
rect 31726 28985 31738 28988
rect 31772 28985 31784 29019
rect 31726 28979 31784 28985
rect 33502 28976 33508 29028
rect 33560 29016 33566 29028
rect 35345 29019 35403 29025
rect 35345 29016 35357 29019
rect 33560 28988 34008 29016
rect 33560 28976 33566 28988
rect 31297 28951 31355 28957
rect 31297 28948 31309 28951
rect 31260 28920 31309 28948
rect 31260 28908 31266 28920
rect 31297 28917 31309 28920
rect 31343 28917 31355 28951
rect 31297 28911 31355 28917
rect 32674 28908 32680 28960
rect 32732 28948 32738 28960
rect 32861 28951 32919 28957
rect 32861 28948 32873 28951
rect 32732 28920 32873 28948
rect 32732 28908 32738 28920
rect 32861 28917 32873 28920
rect 32907 28917 32919 28951
rect 33594 28948 33600 28960
rect 33555 28920 33600 28948
rect 32861 28911 32919 28917
rect 33594 28908 33600 28920
rect 33652 28908 33658 28960
rect 33980 28957 34008 28988
rect 34716 28988 35357 29016
rect 34716 28960 34744 28988
rect 35345 28985 35357 28988
rect 35391 28985 35403 29019
rect 35345 28979 35403 28985
rect 35802 28976 35808 29028
rect 35860 29016 35866 29028
rect 35897 29019 35955 29025
rect 35897 29016 35909 29019
rect 35860 28988 35909 29016
rect 35860 28976 35866 28988
rect 35897 28985 35909 28988
rect 35943 28985 35955 29019
rect 35897 28979 35955 28985
rect 33965 28951 34023 28957
rect 33965 28917 33977 28951
rect 34011 28948 34023 28951
rect 34238 28948 34244 28960
rect 34011 28920 34244 28948
rect 34011 28917 34023 28920
rect 33965 28911 34023 28917
rect 34238 28908 34244 28920
rect 34296 28908 34302 28960
rect 34698 28948 34704 28960
rect 34659 28920 34704 28948
rect 34698 28908 34704 28920
rect 34756 28908 34762 28960
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 2774 28704 2780 28756
rect 2832 28744 2838 28756
rect 3145 28747 3203 28753
rect 3145 28744 3157 28747
rect 2832 28716 3157 28744
rect 2832 28704 2838 28716
rect 3145 28713 3157 28716
rect 3191 28713 3203 28747
rect 3145 28707 3203 28713
rect 3329 28747 3387 28753
rect 3329 28713 3341 28747
rect 3375 28744 3387 28747
rect 3513 28747 3571 28753
rect 3513 28744 3525 28747
rect 3375 28716 3525 28744
rect 3375 28713 3387 28716
rect 3329 28707 3387 28713
rect 3513 28713 3525 28716
rect 3559 28744 3571 28747
rect 3878 28744 3884 28756
rect 3559 28716 3884 28744
rect 3559 28713 3571 28716
rect 3513 28707 3571 28713
rect 3878 28704 3884 28716
rect 3936 28704 3942 28756
rect 4614 28704 4620 28756
rect 4672 28744 4678 28756
rect 5445 28747 5503 28753
rect 5445 28744 5457 28747
rect 4672 28716 5457 28744
rect 4672 28704 4678 28716
rect 5445 28713 5457 28716
rect 5491 28713 5503 28747
rect 5810 28744 5816 28756
rect 5771 28716 5816 28744
rect 5445 28707 5503 28713
rect 5810 28704 5816 28716
rect 5868 28704 5874 28756
rect 8294 28704 8300 28756
rect 8352 28744 8358 28756
rect 8481 28747 8539 28753
rect 8481 28744 8493 28747
rect 8352 28716 8493 28744
rect 8352 28704 8358 28716
rect 8481 28713 8493 28716
rect 8527 28713 8539 28747
rect 8481 28707 8539 28713
rect 9861 28747 9919 28753
rect 9861 28713 9873 28747
rect 9907 28744 9919 28747
rect 10226 28744 10232 28756
rect 9907 28716 10232 28744
rect 9907 28713 9919 28716
rect 9861 28707 9919 28713
rect 10226 28704 10232 28716
rect 10284 28704 10290 28756
rect 10594 28744 10600 28756
rect 10555 28716 10600 28744
rect 10594 28704 10600 28716
rect 10652 28704 10658 28756
rect 13357 28747 13415 28753
rect 13357 28713 13369 28747
rect 13403 28744 13415 28747
rect 14093 28747 14151 28753
rect 14093 28744 14105 28747
rect 13403 28716 14105 28744
rect 13403 28713 13415 28716
rect 13357 28707 13415 28713
rect 14093 28713 14105 28716
rect 14139 28744 14151 28747
rect 14458 28744 14464 28756
rect 14139 28716 14464 28744
rect 14139 28713 14151 28716
rect 14093 28707 14151 28713
rect 14458 28704 14464 28716
rect 14516 28704 14522 28756
rect 15286 28704 15292 28756
rect 15344 28744 15350 28756
rect 15657 28747 15715 28753
rect 15657 28744 15669 28747
rect 15344 28716 15669 28744
rect 15344 28704 15350 28716
rect 15657 28713 15669 28716
rect 15703 28713 15715 28747
rect 15657 28707 15715 28713
rect 18785 28747 18843 28753
rect 18785 28713 18797 28747
rect 18831 28744 18843 28747
rect 19242 28744 19248 28756
rect 18831 28716 19248 28744
rect 18831 28713 18843 28716
rect 18785 28707 18843 28713
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 19613 28747 19671 28753
rect 19613 28713 19625 28747
rect 19659 28744 19671 28747
rect 20070 28744 20076 28756
rect 19659 28716 20076 28744
rect 19659 28713 19671 28716
rect 19613 28707 19671 28713
rect 1854 28636 1860 28688
rect 1912 28676 1918 28688
rect 2032 28679 2090 28685
rect 2032 28676 2044 28679
rect 1912 28648 2044 28676
rect 1912 28636 1918 28648
rect 2032 28645 2044 28648
rect 2078 28676 2090 28679
rect 2498 28676 2504 28688
rect 2078 28648 2504 28676
rect 2078 28645 2090 28648
rect 2032 28639 2090 28645
rect 2498 28636 2504 28648
rect 2556 28636 2562 28688
rect 3896 28608 3924 28704
rect 4154 28636 4160 28688
rect 4212 28676 4218 28688
rect 4310 28679 4368 28685
rect 4310 28676 4322 28679
rect 4212 28648 4322 28676
rect 4212 28636 4218 28648
rect 4310 28645 4322 28648
rect 4356 28645 4368 28679
rect 4310 28639 4368 28645
rect 11232 28679 11290 28685
rect 11232 28645 11244 28679
rect 11278 28676 11290 28679
rect 12342 28676 12348 28688
rect 11278 28648 12348 28676
rect 11278 28645 11290 28648
rect 11232 28639 11290 28645
rect 12342 28636 12348 28648
rect 12400 28636 12406 28688
rect 14274 28636 14280 28688
rect 14332 28676 14338 28688
rect 14369 28679 14427 28685
rect 14369 28676 14381 28679
rect 14332 28648 14381 28676
rect 14332 28636 14338 28648
rect 14369 28645 14381 28648
rect 14415 28645 14427 28679
rect 14369 28639 14427 28645
rect 15194 28636 15200 28688
rect 15252 28676 15258 28688
rect 15749 28679 15807 28685
rect 15749 28676 15761 28679
rect 15252 28648 15761 28676
rect 15252 28636 15258 28648
rect 15749 28645 15761 28648
rect 15795 28676 15807 28679
rect 15838 28676 15844 28688
rect 15795 28648 15844 28676
rect 15795 28645 15807 28648
rect 15749 28639 15807 28645
rect 15838 28636 15844 28648
rect 15896 28636 15902 28688
rect 19058 28676 19064 28688
rect 19019 28648 19064 28676
rect 19058 28636 19064 28648
rect 19116 28636 19122 28688
rect 19518 28636 19524 28688
rect 19576 28676 19582 28688
rect 19628 28676 19656 28707
rect 20070 28704 20076 28716
rect 20128 28704 20134 28756
rect 20717 28747 20775 28753
rect 20717 28713 20729 28747
rect 20763 28744 20775 28747
rect 20806 28744 20812 28756
rect 20763 28716 20812 28744
rect 20763 28713 20775 28716
rect 20717 28707 20775 28713
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 22094 28704 22100 28756
rect 22152 28744 22158 28756
rect 22281 28747 22339 28753
rect 22281 28744 22293 28747
rect 22152 28716 22293 28744
rect 22152 28704 22158 28716
rect 22281 28713 22293 28716
rect 22327 28713 22339 28747
rect 23658 28744 23664 28756
rect 23619 28716 23664 28744
rect 22281 28707 22339 28713
rect 23658 28704 23664 28716
rect 23716 28704 23722 28756
rect 24121 28747 24179 28753
rect 24121 28713 24133 28747
rect 24167 28744 24179 28747
rect 24762 28744 24768 28756
rect 24167 28716 24768 28744
rect 24167 28713 24179 28716
rect 24121 28707 24179 28713
rect 24762 28704 24768 28716
rect 24820 28704 24826 28756
rect 31202 28744 31208 28756
rect 31163 28716 31208 28744
rect 31202 28704 31208 28716
rect 31260 28704 31266 28756
rect 33594 28704 33600 28756
rect 33652 28744 33658 28756
rect 33781 28747 33839 28753
rect 33781 28744 33793 28747
rect 33652 28716 33793 28744
rect 33652 28704 33658 28716
rect 33781 28713 33793 28716
rect 33827 28713 33839 28747
rect 33781 28707 33839 28713
rect 35710 28704 35716 28756
rect 35768 28744 35774 28756
rect 35989 28747 36047 28753
rect 35989 28744 36001 28747
rect 35768 28716 36001 28744
rect 35768 28704 35774 28716
rect 35989 28713 36001 28716
rect 36035 28713 36047 28747
rect 35989 28707 36047 28713
rect 19576 28648 19656 28676
rect 19576 28636 19582 28648
rect 4065 28611 4123 28617
rect 4065 28608 4077 28611
rect 3896 28580 4077 28608
rect 4065 28577 4077 28580
rect 4111 28577 4123 28611
rect 4065 28571 4123 28577
rect 7282 28568 7288 28620
rect 7340 28608 7346 28620
rect 8386 28608 8392 28620
rect 7340 28580 8392 28608
rect 7340 28568 7346 28580
rect 8386 28568 8392 28580
rect 8444 28608 8450 28620
rect 9122 28608 9128 28620
rect 8444 28580 9128 28608
rect 8444 28568 8450 28580
rect 9122 28568 9128 28580
rect 9180 28568 9186 28620
rect 9677 28611 9735 28617
rect 9677 28577 9689 28611
rect 9723 28608 9735 28611
rect 10226 28608 10232 28620
rect 9723 28580 10232 28608
rect 9723 28577 9735 28580
rect 9677 28571 9735 28577
rect 10226 28568 10232 28580
rect 10284 28568 10290 28620
rect 12618 28568 12624 28620
rect 12676 28608 12682 28620
rect 13173 28611 13231 28617
rect 13173 28608 13185 28611
rect 12676 28580 13185 28608
rect 12676 28568 12682 28580
rect 13173 28577 13185 28580
rect 13219 28608 13231 28611
rect 13446 28608 13452 28620
rect 13219 28580 13452 28608
rect 13219 28577 13231 28580
rect 13173 28571 13231 28577
rect 13446 28568 13452 28580
rect 13504 28568 13510 28620
rect 20824 28608 20852 28704
rect 21174 28617 21180 28620
rect 20901 28611 20959 28617
rect 20901 28608 20913 28611
rect 20824 28580 20913 28608
rect 20901 28577 20913 28580
rect 20947 28577 20959 28611
rect 21168 28608 21180 28617
rect 21135 28580 21180 28608
rect 20901 28571 20959 28577
rect 21168 28571 21180 28580
rect 21174 28568 21180 28571
rect 21232 28568 21238 28620
rect 23676 28608 23704 28704
rect 24480 28679 24538 28685
rect 24480 28645 24492 28679
rect 24526 28676 24538 28679
rect 26142 28676 26148 28688
rect 24526 28648 26148 28676
rect 24526 28645 24538 28648
rect 24480 28639 24538 28645
rect 26142 28636 26148 28648
rect 26200 28636 26206 28688
rect 34146 28636 34152 28688
rect 34204 28676 34210 28688
rect 34974 28676 34980 28688
rect 34204 28648 34980 28676
rect 34204 28636 34210 28648
rect 34974 28636 34980 28648
rect 35032 28636 35038 28688
rect 24213 28611 24271 28617
rect 24213 28608 24225 28611
rect 23676 28580 24225 28608
rect 24213 28577 24225 28580
rect 24259 28577 24271 28611
rect 24213 28571 24271 28577
rect 25590 28568 25596 28620
rect 25648 28608 25654 28620
rect 26769 28611 26827 28617
rect 26769 28608 26781 28611
rect 25648 28580 26781 28608
rect 25648 28568 25654 28580
rect 26769 28577 26781 28580
rect 26815 28608 26827 28611
rect 27246 28608 27252 28620
rect 26815 28580 27252 28608
rect 26815 28577 26827 28580
rect 26769 28571 26827 28577
rect 27246 28568 27252 28580
rect 27304 28568 27310 28620
rect 29914 28568 29920 28620
rect 29972 28608 29978 28620
rect 30081 28611 30139 28617
rect 30081 28608 30093 28611
rect 29972 28580 30093 28608
rect 29972 28568 29978 28580
rect 30081 28577 30093 28580
rect 30127 28577 30139 28611
rect 30081 28571 30139 28577
rect 32214 28568 32220 28620
rect 32272 28608 32278 28620
rect 32674 28617 32680 28620
rect 32657 28611 32680 28617
rect 32657 28608 32669 28611
rect 32272 28580 32669 28608
rect 32272 28568 32278 28580
rect 32657 28577 32669 28580
rect 32732 28608 32738 28620
rect 32732 28580 32805 28608
rect 32657 28571 32680 28577
rect 32674 28568 32680 28571
rect 32732 28568 32738 28580
rect 34698 28568 34704 28620
rect 34756 28608 34762 28620
rect 34865 28611 34923 28617
rect 34865 28608 34877 28611
rect 34756 28580 34877 28608
rect 34756 28568 34762 28580
rect 34865 28577 34877 28580
rect 34911 28577 34923 28611
rect 34865 28571 34923 28577
rect 1765 28543 1823 28549
rect 1765 28509 1777 28543
rect 1811 28509 1823 28543
rect 1765 28503 1823 28509
rect 7469 28543 7527 28549
rect 7469 28509 7481 28543
rect 7515 28540 7527 28543
rect 8662 28540 8668 28552
rect 7515 28512 8668 28540
rect 7515 28509 7527 28512
rect 7469 28503 7527 28509
rect 1780 28404 1808 28503
rect 8662 28500 8668 28512
rect 8720 28500 8726 28552
rect 9490 28540 9496 28552
rect 9403 28512 9496 28540
rect 9490 28500 9496 28512
rect 9548 28540 9554 28552
rect 9766 28540 9772 28552
rect 9548 28512 9772 28540
rect 9548 28500 9554 28512
rect 9766 28500 9772 28512
rect 9824 28540 9830 28552
rect 10965 28543 11023 28549
rect 10965 28540 10977 28543
rect 9824 28512 10977 28540
rect 9824 28500 9830 28512
rect 10965 28509 10977 28512
rect 11011 28509 11023 28543
rect 10965 28503 11023 28509
rect 14642 28500 14648 28552
rect 14700 28540 14706 28552
rect 15562 28540 15568 28552
rect 14700 28512 15568 28540
rect 14700 28500 14706 28512
rect 15562 28500 15568 28512
rect 15620 28540 15626 28552
rect 15841 28543 15899 28549
rect 15841 28540 15853 28543
rect 15620 28512 15853 28540
rect 15620 28500 15626 28512
rect 15841 28509 15853 28512
rect 15887 28509 15899 28543
rect 16850 28540 16856 28552
rect 16811 28512 16856 28540
rect 15841 28503 15899 28509
rect 16850 28500 16856 28512
rect 16908 28500 16914 28552
rect 19702 28540 19708 28552
rect 19663 28512 19708 28540
rect 19702 28500 19708 28512
rect 19760 28500 19766 28552
rect 19794 28500 19800 28552
rect 19852 28540 19858 28552
rect 20714 28540 20720 28552
rect 19852 28512 20720 28540
rect 19852 28500 19858 28512
rect 20714 28500 20720 28512
rect 20772 28500 20778 28552
rect 23201 28543 23259 28549
rect 23201 28509 23213 28543
rect 23247 28540 23259 28543
rect 23842 28540 23848 28552
rect 23247 28512 23848 28540
rect 23247 28509 23259 28512
rect 23201 28503 23259 28509
rect 23842 28500 23848 28512
rect 23900 28500 23906 28552
rect 26510 28540 26516 28552
rect 26423 28512 26516 28540
rect 26510 28500 26516 28512
rect 26568 28500 26574 28552
rect 29733 28543 29791 28549
rect 29733 28509 29745 28543
rect 29779 28540 29791 28543
rect 29822 28540 29828 28552
rect 29779 28512 29828 28540
rect 29779 28509 29791 28512
rect 29733 28503 29791 28509
rect 29822 28500 29828 28512
rect 29880 28500 29886 28552
rect 32401 28543 32459 28549
rect 32401 28509 32413 28543
rect 32447 28509 32459 28543
rect 34609 28543 34667 28549
rect 34609 28540 34621 28543
rect 32401 28503 32459 28509
rect 34440 28512 34621 28540
rect 8021 28475 8079 28481
rect 8021 28441 8033 28475
rect 8067 28472 8079 28475
rect 10229 28475 10287 28481
rect 10229 28472 10241 28475
rect 8067 28444 10241 28472
rect 8067 28441 8079 28444
rect 8021 28435 8079 28441
rect 10229 28441 10241 28444
rect 10275 28472 10287 28475
rect 10410 28472 10416 28484
rect 10275 28444 10416 28472
rect 10275 28441 10287 28444
rect 10229 28435 10287 28441
rect 10410 28432 10416 28444
rect 10468 28432 10474 28484
rect 15289 28475 15347 28481
rect 15289 28441 15301 28475
rect 15335 28472 15347 28475
rect 16482 28472 16488 28484
rect 15335 28444 16488 28472
rect 15335 28441 15347 28444
rect 15289 28435 15347 28441
rect 16482 28432 16488 28444
rect 16540 28432 16546 28484
rect 25498 28432 25504 28484
rect 25556 28472 25562 28484
rect 25869 28475 25927 28481
rect 25869 28472 25881 28475
rect 25556 28444 25881 28472
rect 25556 28432 25562 28444
rect 25869 28441 25881 28444
rect 25915 28472 25927 28475
rect 26528 28472 26556 28500
rect 25915 28444 26556 28472
rect 25915 28441 25927 28444
rect 25869 28435 25927 28441
rect 2038 28404 2044 28416
rect 1780 28376 2044 28404
rect 2038 28364 2044 28376
rect 2096 28404 2102 28416
rect 3329 28407 3387 28413
rect 3329 28404 3341 28407
rect 2096 28376 3341 28404
rect 2096 28364 2102 28376
rect 3329 28373 3341 28376
rect 3375 28373 3387 28407
rect 7834 28404 7840 28416
rect 7795 28376 7840 28404
rect 3329 28367 3387 28373
rect 7834 28364 7840 28376
rect 7892 28364 7898 28416
rect 12345 28407 12403 28413
rect 12345 28373 12357 28407
rect 12391 28404 12403 28407
rect 12621 28407 12679 28413
rect 12621 28404 12633 28407
rect 12391 28376 12633 28404
rect 12391 28373 12403 28376
rect 12345 28367 12403 28373
rect 12621 28373 12633 28376
rect 12667 28404 12679 28407
rect 12802 28404 12808 28416
rect 12667 28376 12808 28404
rect 12667 28373 12679 28376
rect 12621 28367 12679 28373
rect 12802 28364 12808 28376
rect 12860 28364 12866 28416
rect 12986 28404 12992 28416
rect 12947 28376 12992 28404
rect 12986 28364 12992 28376
rect 13044 28364 13050 28416
rect 15010 28364 15016 28416
rect 15068 28404 15074 28416
rect 15105 28407 15163 28413
rect 15105 28404 15117 28407
rect 15068 28376 15117 28404
rect 15068 28364 15074 28376
rect 15105 28373 15117 28376
rect 15151 28404 15163 28407
rect 15378 28404 15384 28416
rect 15151 28376 15384 28404
rect 15151 28373 15163 28376
rect 15105 28367 15163 28373
rect 15378 28364 15384 28376
rect 15436 28364 15442 28416
rect 16298 28404 16304 28416
rect 16259 28376 16304 28404
rect 16298 28364 16304 28376
rect 16356 28364 16362 28416
rect 20346 28404 20352 28416
rect 20259 28376 20352 28404
rect 20346 28364 20352 28376
rect 20404 28404 20410 28416
rect 20530 28404 20536 28416
rect 20404 28376 20536 28404
rect 20404 28364 20410 28376
rect 20530 28364 20536 28376
rect 20588 28364 20594 28416
rect 25590 28404 25596 28416
rect 25551 28376 25596 28404
rect 25590 28364 25596 28376
rect 25648 28364 25654 28416
rect 27890 28404 27896 28416
rect 27851 28376 27896 28404
rect 27890 28364 27896 28376
rect 27948 28364 27954 28416
rect 31478 28364 31484 28416
rect 31536 28404 31542 28416
rect 31573 28407 31631 28413
rect 31573 28404 31585 28407
rect 31536 28376 31585 28404
rect 31536 28364 31542 28376
rect 31573 28373 31585 28376
rect 31619 28404 31631 28407
rect 32416 28404 32444 28503
rect 34238 28404 34244 28416
rect 31619 28376 34244 28404
rect 31619 28373 31631 28376
rect 31573 28367 31631 28373
rect 34238 28364 34244 28376
rect 34296 28404 34302 28416
rect 34440 28413 34468 28512
rect 34609 28509 34621 28512
rect 34655 28509 34667 28543
rect 34609 28503 34667 28509
rect 34425 28407 34483 28413
rect 34425 28404 34437 28407
rect 34296 28376 34437 28404
rect 34296 28364 34302 28376
rect 34425 28373 34437 28376
rect 34471 28373 34483 28407
rect 34425 28367 34483 28373
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 1854 28200 1860 28212
rect 1815 28172 1860 28200
rect 1854 28160 1860 28172
rect 1912 28160 1918 28212
rect 4062 28160 4068 28212
rect 4120 28200 4126 28212
rect 4157 28203 4215 28209
rect 4157 28200 4169 28203
rect 4120 28172 4169 28200
rect 4120 28160 4126 28172
rect 4157 28169 4169 28172
rect 4203 28169 4215 28203
rect 4157 28163 4215 28169
rect 4525 28203 4583 28209
rect 4525 28169 4537 28203
rect 4571 28200 4583 28203
rect 5350 28200 5356 28212
rect 4571 28172 5356 28200
rect 4571 28169 4583 28172
rect 4525 28163 4583 28169
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 7282 28200 7288 28212
rect 7243 28172 7288 28200
rect 7282 28160 7288 28172
rect 7340 28160 7346 28212
rect 8294 28160 8300 28212
rect 8352 28200 8358 28212
rect 8757 28203 8815 28209
rect 8757 28200 8769 28203
rect 8352 28172 8769 28200
rect 8352 28160 8358 28172
rect 8757 28169 8769 28172
rect 8803 28169 8815 28203
rect 8757 28163 8815 28169
rect 9861 28203 9919 28209
rect 9861 28169 9873 28203
rect 9907 28200 9919 28203
rect 10962 28200 10968 28212
rect 9907 28172 10968 28200
rect 9907 28169 9919 28172
rect 9861 28163 9919 28169
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 11885 28203 11943 28209
rect 11885 28169 11897 28203
rect 11931 28200 11943 28203
rect 12253 28203 12311 28209
rect 12253 28200 12265 28203
rect 11931 28172 12265 28200
rect 11931 28169 11943 28172
rect 11885 28163 11943 28169
rect 12253 28169 12265 28172
rect 12299 28200 12311 28203
rect 12342 28200 12348 28212
rect 12299 28172 12348 28200
rect 12299 28169 12311 28172
rect 12253 28163 12311 28169
rect 12342 28160 12348 28172
rect 12400 28200 12406 28212
rect 13446 28200 13452 28212
rect 12400 28172 12940 28200
rect 13407 28172 13452 28200
rect 12400 28160 12406 28172
rect 9585 28135 9643 28141
rect 9585 28101 9597 28135
rect 9631 28132 9643 28135
rect 10781 28135 10839 28141
rect 10781 28132 10793 28135
rect 9631 28104 10793 28132
rect 9631 28101 9643 28104
rect 9585 28095 9643 28101
rect 8389 28067 8447 28073
rect 8389 28033 8401 28067
rect 8435 28064 8447 28067
rect 8662 28064 8668 28076
rect 8435 28036 8668 28064
rect 8435 28033 8447 28036
rect 8389 28027 8447 28033
rect 8662 28024 8668 28036
rect 8720 28064 8726 28076
rect 9214 28064 9220 28076
rect 8720 28036 9220 28064
rect 8720 28024 8726 28036
rect 9214 28024 9220 28036
rect 9272 28024 9278 28076
rect 7558 27956 7564 28008
rect 7616 27996 7622 28008
rect 9692 28005 9720 28104
rect 10781 28101 10793 28104
rect 10827 28101 10839 28135
rect 12437 28135 12495 28141
rect 12437 28132 12449 28135
rect 10781 28095 10839 28101
rect 11256 28104 12449 28132
rect 11256 28073 11284 28104
rect 12437 28101 12449 28104
rect 12483 28101 12495 28135
rect 12437 28095 12495 28101
rect 10689 28067 10747 28073
rect 10689 28033 10701 28067
rect 10735 28064 10747 28067
rect 11241 28067 11299 28073
rect 11241 28064 11253 28067
rect 10735 28036 11253 28064
rect 10735 28033 10747 28036
rect 10689 28027 10747 28033
rect 11241 28033 11253 28036
rect 11287 28033 11299 28067
rect 11241 28027 11299 28033
rect 11330 28024 11336 28076
rect 11388 28064 11394 28076
rect 12912 28073 12940 28172
rect 13446 28160 13452 28172
rect 13504 28160 13510 28212
rect 14642 28200 14648 28212
rect 14603 28172 14648 28200
rect 14642 28160 14648 28172
rect 14700 28160 14706 28212
rect 15286 28200 15292 28212
rect 15247 28172 15292 28200
rect 15286 28160 15292 28172
rect 15344 28160 15350 28212
rect 15473 28203 15531 28209
rect 15473 28169 15485 28203
rect 15519 28200 15531 28203
rect 16298 28200 16304 28212
rect 15519 28172 16304 28200
rect 15519 28169 15531 28172
rect 15473 28163 15531 28169
rect 16298 28160 16304 28172
rect 16356 28160 16362 28212
rect 16390 28160 16396 28212
rect 16448 28200 16454 28212
rect 16485 28203 16543 28209
rect 16485 28200 16497 28203
rect 16448 28172 16497 28200
rect 16448 28160 16454 28172
rect 16485 28169 16497 28172
rect 16531 28169 16543 28203
rect 16485 28163 16543 28169
rect 19337 28203 19395 28209
rect 19337 28169 19349 28203
rect 19383 28200 19395 28203
rect 19518 28200 19524 28212
rect 19383 28172 19524 28200
rect 19383 28169 19395 28172
rect 19337 28163 19395 28169
rect 19518 28160 19524 28172
rect 19576 28160 19582 28212
rect 19702 28160 19708 28212
rect 19760 28200 19766 28212
rect 19978 28200 19984 28212
rect 19760 28172 19984 28200
rect 19760 28160 19766 28172
rect 19978 28160 19984 28172
rect 20036 28200 20042 28212
rect 20073 28203 20131 28209
rect 20073 28200 20085 28203
rect 20036 28172 20085 28200
rect 20036 28160 20042 28172
rect 20073 28169 20085 28172
rect 20119 28169 20131 28203
rect 23842 28200 23848 28212
rect 23803 28172 23848 28200
rect 20073 28163 20131 28169
rect 23842 28160 23848 28172
rect 23900 28160 23906 28212
rect 27246 28200 27252 28212
rect 27207 28172 27252 28200
rect 27246 28160 27252 28172
rect 27304 28160 27310 28212
rect 29641 28203 29699 28209
rect 29641 28169 29653 28203
rect 29687 28200 29699 28203
rect 29914 28200 29920 28212
rect 29687 28172 29920 28200
rect 29687 28169 29699 28172
rect 29641 28163 29699 28169
rect 29914 28160 29920 28172
rect 29972 28200 29978 28212
rect 31481 28203 31539 28209
rect 31481 28200 31493 28203
rect 29972 28172 31493 28200
rect 29972 28160 29978 28172
rect 31481 28169 31493 28172
rect 31527 28169 31539 28203
rect 32214 28200 32220 28212
rect 32175 28172 32220 28200
rect 31481 28163 31539 28169
rect 16408 28132 16436 28160
rect 15948 28104 16436 28132
rect 18969 28135 19027 28141
rect 12897 28067 12955 28073
rect 11388 28036 11433 28064
rect 11388 28024 11394 28036
rect 12897 28033 12909 28067
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 12986 28024 12992 28076
rect 13044 28064 13050 28076
rect 15948 28073 15976 28104
rect 18969 28101 18981 28135
rect 19015 28132 19027 28135
rect 19794 28132 19800 28144
rect 19015 28104 19800 28132
rect 19015 28101 19027 28104
rect 18969 28095 19027 28101
rect 19794 28092 19800 28104
rect 19852 28092 19858 28144
rect 23750 28092 23756 28144
rect 23808 28132 23814 28144
rect 24029 28135 24087 28141
rect 24029 28132 24041 28135
rect 23808 28104 24041 28132
rect 23808 28092 23814 28104
rect 24029 28101 24041 28104
rect 24075 28101 24087 28135
rect 24029 28095 24087 28101
rect 15933 28067 15991 28073
rect 13044 28036 13089 28064
rect 13044 28024 13050 28036
rect 15933 28033 15945 28067
rect 15979 28033 15991 28067
rect 15933 28027 15991 28033
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16301 28067 16359 28073
rect 16301 28064 16313 28067
rect 16163 28036 16313 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16301 28033 16313 28036
rect 16347 28064 16359 28067
rect 16482 28064 16488 28076
rect 16347 28036 16488 28064
rect 16347 28033 16359 28036
rect 16301 28027 16359 28033
rect 16482 28024 16488 28036
rect 16540 28024 16546 28076
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 19613 28067 19671 28073
rect 19613 28064 19625 28067
rect 19484 28036 19625 28064
rect 19484 28024 19490 28036
rect 19613 28033 19625 28036
rect 19659 28033 19671 28067
rect 19613 28027 19671 28033
rect 23477 28067 23535 28073
rect 23477 28033 23489 28067
rect 23523 28064 23535 28067
rect 24673 28067 24731 28073
rect 24673 28064 24685 28067
rect 23523 28036 24685 28064
rect 23523 28033 23535 28036
rect 23477 28027 23535 28033
rect 24673 28033 24685 28036
rect 24719 28064 24731 28067
rect 25501 28067 25559 28073
rect 25501 28064 25513 28067
rect 24719 28036 25513 28064
rect 24719 28033 24731 28036
rect 24673 28027 24731 28033
rect 25501 28033 25513 28036
rect 25547 28064 25559 28067
rect 31496 28064 31524 28163
rect 32214 28160 32220 28172
rect 32272 28160 32278 28212
rect 34698 28200 34704 28212
rect 34659 28172 34704 28200
rect 34698 28160 34704 28172
rect 34756 28160 34762 28212
rect 31941 28067 31999 28073
rect 31941 28064 31953 28067
rect 25547 28036 25728 28064
rect 31496 28036 31953 28064
rect 25547 28033 25559 28036
rect 25501 28027 25559 28033
rect 8205 27999 8263 28005
rect 8205 27996 8217 27999
rect 7616 27968 8217 27996
rect 7616 27956 7622 27968
rect 8205 27965 8217 27968
rect 8251 27965 8263 27999
rect 8205 27959 8263 27965
rect 9677 27999 9735 28005
rect 9677 27965 9689 27999
rect 9723 27965 9735 27999
rect 12802 27996 12808 28008
rect 12763 27968 12808 27996
rect 9677 27959 9735 27965
rect 12802 27956 12808 27968
rect 12860 27956 12866 28008
rect 15562 27956 15568 28008
rect 15620 27996 15626 28008
rect 15841 27999 15899 28005
rect 15841 27996 15853 27999
rect 15620 27968 15853 27996
rect 15620 27956 15626 27968
rect 15841 27965 15853 27968
rect 15887 27996 15899 27999
rect 16850 27996 16856 28008
rect 15887 27968 16856 27996
rect 15887 27965 15899 27968
rect 15841 27959 15899 27965
rect 16850 27956 16856 27968
rect 16908 27956 16914 28008
rect 20717 27999 20775 28005
rect 20717 27965 20729 27999
rect 20763 27996 20775 27999
rect 20806 27996 20812 28008
rect 20763 27968 20812 27996
rect 20763 27965 20775 27968
rect 20717 27959 20775 27965
rect 20806 27956 20812 27968
rect 20864 27956 20870 28008
rect 23842 27956 23848 28008
rect 23900 27996 23906 28008
rect 24397 27999 24455 28005
rect 24397 27996 24409 27999
rect 23900 27968 24409 27996
rect 23900 27956 23906 27968
rect 24397 27965 24409 27968
rect 24443 27965 24455 27999
rect 24397 27959 24455 27965
rect 25406 27956 25412 28008
rect 25464 27996 25470 28008
rect 25593 27999 25651 28005
rect 25593 27996 25605 27999
rect 25464 27968 25605 27996
rect 25464 27956 25470 27968
rect 25593 27965 25605 27968
rect 25639 27965 25651 27999
rect 25700 27996 25728 28036
rect 31941 28033 31953 28036
rect 31987 28033 31999 28067
rect 31941 28027 31999 28033
rect 32766 28024 32772 28076
rect 32824 28064 32830 28076
rect 32953 28067 33011 28073
rect 32953 28064 32965 28067
rect 32824 28036 32965 28064
rect 32824 28024 32830 28036
rect 32953 28033 32965 28036
rect 32999 28064 33011 28067
rect 33042 28064 33048 28076
rect 32999 28036 33048 28064
rect 32999 28033 33011 28036
rect 32953 28027 33011 28033
rect 33042 28024 33048 28036
rect 33100 28064 33106 28076
rect 33778 28064 33784 28076
rect 33100 28036 33784 28064
rect 33100 28024 33106 28036
rect 33778 28024 33784 28036
rect 33836 28024 33842 28076
rect 25866 28005 25872 28008
rect 25860 27996 25872 28005
rect 25700 27968 25872 27996
rect 25593 27959 25651 27965
rect 25860 27959 25872 27968
rect 25866 27956 25872 27959
rect 25924 27956 25930 28008
rect 29089 27999 29147 28005
rect 29089 27965 29101 27999
rect 29135 27996 29147 27999
rect 29822 27996 29828 28008
rect 29135 27968 29828 27996
rect 29135 27965 29147 27968
rect 29089 27959 29147 27965
rect 29822 27956 29828 27968
rect 29880 27996 29886 28008
rect 30101 27999 30159 28005
rect 30101 27996 30113 27999
rect 29880 27968 30113 27996
rect 29880 27956 29886 27968
rect 30101 27965 30113 27968
rect 30147 27996 30159 27999
rect 30147 27968 31156 27996
rect 30147 27965 30159 27968
rect 30101 27959 30159 27965
rect 7282 27888 7288 27940
rect 7340 27928 7346 27940
rect 7834 27928 7840 27940
rect 7340 27900 7840 27928
rect 7340 27888 7346 27900
rect 7834 27888 7840 27900
rect 7892 27928 7898 27940
rect 8113 27931 8171 27937
rect 8113 27928 8125 27931
rect 7892 27900 8125 27928
rect 7892 27888 7898 27900
rect 8113 27897 8125 27900
rect 8159 27897 8171 27931
rect 8113 27891 8171 27897
rect 15013 27931 15071 27937
rect 15013 27897 15025 27931
rect 15059 27928 15071 27931
rect 15286 27928 15292 27940
rect 15059 27900 15292 27928
rect 15059 27897 15071 27900
rect 15013 27891 15071 27897
rect 15286 27888 15292 27900
rect 15344 27928 15350 27940
rect 16301 27931 16359 27937
rect 16301 27928 16313 27931
rect 15344 27900 16313 27928
rect 15344 27888 15350 27900
rect 16301 27897 16313 27900
rect 16347 27897 16359 27931
rect 16301 27891 16359 27897
rect 20984 27931 21042 27937
rect 20984 27897 20996 27931
rect 21030 27928 21042 27931
rect 21818 27928 21824 27940
rect 21030 27900 21824 27928
rect 21030 27897 21042 27900
rect 20984 27891 21042 27897
rect 21818 27888 21824 27900
rect 21876 27928 21882 27940
rect 22373 27931 22431 27937
rect 22373 27928 22385 27931
rect 21876 27900 22385 27928
rect 21876 27888 21882 27900
rect 22373 27897 22385 27900
rect 22419 27897 22431 27931
rect 22373 27891 22431 27897
rect 25133 27931 25191 27937
rect 25133 27897 25145 27931
rect 25179 27928 25191 27931
rect 26142 27928 26148 27940
rect 25179 27900 26148 27928
rect 25179 27897 25191 27900
rect 25133 27891 25191 27897
rect 26142 27888 26148 27900
rect 26200 27888 26206 27940
rect 30009 27931 30067 27937
rect 30009 27897 30021 27931
rect 30055 27928 30067 27931
rect 30346 27931 30404 27937
rect 30346 27928 30358 27931
rect 30055 27900 30358 27928
rect 30055 27897 30067 27900
rect 30009 27891 30067 27897
rect 30346 27897 30358 27900
rect 30392 27928 30404 27931
rect 31018 27928 31024 27940
rect 30392 27900 31024 27928
rect 30392 27897 30404 27900
rect 30346 27891 30404 27897
rect 31018 27888 31024 27900
rect 31076 27888 31082 27940
rect 31128 27928 31156 27968
rect 31202 27956 31208 28008
rect 31260 27996 31266 28008
rect 34977 27999 35035 28005
rect 34977 27996 34989 27999
rect 31260 27968 32904 27996
rect 31260 27956 31266 27968
rect 31478 27928 31484 27940
rect 31128 27900 31484 27928
rect 31478 27888 31484 27900
rect 31536 27888 31542 27940
rect 31849 27931 31907 27937
rect 31849 27897 31861 27931
rect 31895 27928 31907 27931
rect 31941 27931 31999 27937
rect 31941 27928 31953 27931
rect 31895 27900 31953 27928
rect 31895 27897 31907 27900
rect 31849 27891 31907 27897
rect 31941 27897 31953 27900
rect 31987 27928 31999 27931
rect 32769 27931 32827 27937
rect 32769 27928 32781 27931
rect 31987 27900 32781 27928
rect 31987 27897 31999 27900
rect 31941 27891 31999 27897
rect 32769 27897 32781 27900
rect 32815 27897 32827 27931
rect 32769 27891 32827 27897
rect 2038 27820 2044 27872
rect 2096 27860 2102 27872
rect 2133 27863 2191 27869
rect 2133 27860 2145 27863
rect 2096 27832 2145 27860
rect 2096 27820 2102 27832
rect 2133 27829 2145 27832
rect 2179 27829 2191 27863
rect 7558 27860 7564 27872
rect 7519 27832 7564 27860
rect 2133 27823 2191 27829
rect 7558 27820 7564 27832
rect 7616 27820 7622 27872
rect 7742 27860 7748 27872
rect 7703 27832 7748 27860
rect 7742 27820 7748 27832
rect 7800 27820 7806 27872
rect 9214 27860 9220 27872
rect 9175 27832 9220 27860
rect 9214 27820 9220 27832
rect 9272 27820 9278 27872
rect 10226 27860 10232 27872
rect 10187 27832 10232 27860
rect 10226 27820 10232 27832
rect 10284 27820 10290 27872
rect 11146 27860 11152 27872
rect 11107 27832 11152 27860
rect 11146 27820 11152 27832
rect 11204 27820 11210 27872
rect 20625 27863 20683 27869
rect 20625 27829 20637 27863
rect 20671 27860 20683 27863
rect 21174 27860 21180 27872
rect 20671 27832 21180 27860
rect 20671 27829 20683 27832
rect 20625 27823 20683 27829
rect 21174 27820 21180 27832
rect 21232 27860 21238 27872
rect 22094 27860 22100 27872
rect 21232 27832 22100 27860
rect 21232 27820 21238 27832
rect 22094 27820 22100 27832
rect 22152 27860 22158 27872
rect 22152 27832 22245 27860
rect 22152 27820 22158 27832
rect 24486 27820 24492 27872
rect 24544 27860 24550 27872
rect 26973 27863 27031 27869
rect 24544 27832 24589 27860
rect 24544 27820 24550 27832
rect 26973 27829 26985 27863
rect 27019 27860 27031 27863
rect 27062 27860 27068 27872
rect 27019 27832 27068 27860
rect 27019 27829 27031 27832
rect 26973 27823 27031 27829
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 32306 27860 32312 27872
rect 32267 27832 32312 27860
rect 32306 27820 32312 27832
rect 32364 27820 32370 27872
rect 32677 27863 32735 27869
rect 32677 27829 32689 27863
rect 32723 27860 32735 27863
rect 32876 27860 32904 27968
rect 34716 27968 34989 27996
rect 33962 27888 33968 27940
rect 34020 27928 34026 27940
rect 34606 27928 34612 27940
rect 34020 27900 34612 27928
rect 34020 27888 34026 27900
rect 34606 27888 34612 27900
rect 34664 27888 34670 27940
rect 34716 27872 34744 27968
rect 34977 27965 34989 27968
rect 35023 27965 35035 27999
rect 34977 27959 35035 27965
rect 34992 27928 35020 27959
rect 35066 27956 35072 28008
rect 35124 27996 35130 28008
rect 35244 27999 35302 28005
rect 35244 27996 35256 27999
rect 35124 27968 35256 27996
rect 35124 27956 35130 27968
rect 35244 27965 35256 27968
rect 35290 27996 35302 27999
rect 35710 27996 35716 28008
rect 35290 27968 35716 27996
rect 35290 27965 35302 27968
rect 35244 27959 35302 27965
rect 35710 27956 35716 27968
rect 35768 27956 35774 28008
rect 36633 27931 36691 27937
rect 36633 27928 36645 27931
rect 34992 27900 36645 27928
rect 36633 27897 36645 27900
rect 36679 27928 36691 27931
rect 37458 27928 37464 27940
rect 36679 27900 37464 27928
rect 36679 27897 36691 27900
rect 36633 27891 36691 27897
rect 37458 27888 37464 27900
rect 37516 27888 37522 27940
rect 33321 27863 33379 27869
rect 33321 27860 33333 27863
rect 32723 27832 33333 27860
rect 32723 27829 32735 27832
rect 32677 27823 32735 27829
rect 33321 27829 33333 27832
rect 33367 27829 33379 27863
rect 33778 27860 33784 27872
rect 33739 27832 33784 27860
rect 33321 27823 33379 27829
rect 33778 27820 33784 27832
rect 33836 27820 33842 27872
rect 34149 27863 34207 27869
rect 34149 27829 34161 27863
rect 34195 27860 34207 27863
rect 34238 27860 34244 27872
rect 34195 27832 34244 27860
rect 34195 27829 34207 27832
rect 34149 27823 34207 27829
rect 34238 27820 34244 27832
rect 34296 27860 34302 27872
rect 34698 27860 34704 27872
rect 34296 27832 34704 27860
rect 34296 27820 34302 27832
rect 34698 27820 34704 27832
rect 34756 27820 34762 27872
rect 36354 27860 36360 27872
rect 36315 27832 36360 27860
rect 36354 27820 36360 27832
rect 36412 27820 36418 27872
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 2498 27616 2504 27668
rect 2556 27656 2562 27668
rect 2777 27659 2835 27665
rect 2777 27656 2789 27659
rect 2556 27628 2789 27656
rect 2556 27616 2562 27628
rect 2777 27625 2789 27628
rect 2823 27625 2835 27659
rect 2777 27619 2835 27625
rect 8294 27616 8300 27668
rect 8352 27656 8358 27668
rect 8573 27659 8631 27665
rect 8573 27656 8585 27659
rect 8352 27628 8585 27656
rect 8352 27616 8358 27628
rect 8573 27625 8585 27628
rect 8619 27625 8631 27659
rect 9490 27656 9496 27668
rect 9451 27628 9496 27656
rect 8573 27619 8631 27625
rect 9490 27616 9496 27628
rect 9548 27616 9554 27668
rect 11146 27656 11152 27668
rect 10980 27628 11152 27656
rect 2038 27588 2044 27600
rect 1412 27560 2044 27588
rect 1412 27529 1440 27560
rect 2038 27548 2044 27560
rect 2096 27548 2102 27600
rect 9508 27588 9536 27616
rect 7208 27560 9536 27588
rect 10873 27591 10931 27597
rect 1670 27529 1676 27532
rect 1397 27523 1455 27529
rect 1397 27489 1409 27523
rect 1443 27489 1455 27523
rect 1664 27520 1676 27529
rect 1631 27492 1676 27520
rect 1397 27483 1455 27489
rect 1664 27483 1676 27492
rect 1670 27480 1676 27483
rect 1728 27480 1734 27532
rect 6638 27480 6644 27532
rect 6696 27520 6702 27532
rect 7208 27529 7236 27560
rect 10873 27557 10885 27591
rect 10919 27588 10931 27591
rect 10980 27588 11008 27628
rect 11146 27616 11152 27628
rect 11204 27656 11210 27668
rect 12250 27656 12256 27668
rect 11204 27628 12256 27656
rect 11204 27616 11210 27628
rect 12250 27616 12256 27628
rect 12308 27616 12314 27668
rect 12342 27616 12348 27668
rect 12400 27656 12406 27668
rect 12802 27656 12808 27668
rect 12400 27628 12808 27656
rect 12400 27616 12406 27628
rect 12802 27616 12808 27628
rect 12860 27616 12866 27668
rect 15562 27656 15568 27668
rect 15523 27628 15568 27656
rect 15562 27616 15568 27628
rect 15620 27616 15626 27668
rect 15838 27656 15844 27668
rect 15799 27628 15844 27656
rect 15838 27616 15844 27628
rect 15896 27616 15902 27668
rect 20806 27616 20812 27668
rect 20864 27656 20870 27668
rect 21913 27659 21971 27665
rect 21913 27656 21925 27659
rect 20864 27628 21925 27656
rect 20864 27616 20870 27628
rect 21913 27625 21925 27628
rect 21959 27625 21971 27659
rect 21913 27619 21971 27625
rect 23753 27659 23811 27665
rect 23753 27625 23765 27659
rect 23799 27656 23811 27659
rect 24486 27656 24492 27668
rect 23799 27628 24492 27656
rect 23799 27625 23811 27628
rect 23753 27619 23811 27625
rect 24486 27616 24492 27628
rect 24544 27656 24550 27668
rect 24857 27659 24915 27665
rect 24857 27656 24869 27659
rect 24544 27628 24869 27656
rect 24544 27616 24550 27628
rect 24857 27625 24869 27628
rect 24903 27625 24915 27659
rect 31018 27656 31024 27668
rect 30979 27628 31024 27656
rect 24857 27619 24915 27625
rect 31018 27616 31024 27628
rect 31076 27616 31082 27668
rect 32306 27616 32312 27668
rect 32364 27656 32370 27668
rect 32585 27659 32643 27665
rect 32585 27656 32597 27659
rect 32364 27628 32597 27656
rect 32364 27616 32370 27628
rect 32585 27625 32597 27628
rect 32631 27625 32643 27659
rect 35066 27656 35072 27668
rect 35027 27628 35072 27656
rect 32585 27619 32643 27625
rect 35066 27616 35072 27628
rect 35124 27616 35130 27668
rect 21266 27588 21272 27600
rect 10919 27560 11008 27588
rect 21227 27560 21272 27588
rect 10919 27557 10931 27560
rect 10873 27551 10931 27557
rect 21266 27548 21272 27560
rect 21324 27548 21330 27600
rect 24121 27591 24179 27597
rect 24121 27557 24133 27591
rect 24167 27588 24179 27591
rect 25225 27591 25283 27597
rect 25225 27588 25237 27591
rect 24167 27560 25237 27588
rect 24167 27557 24179 27560
rect 24121 27551 24179 27557
rect 25225 27557 25237 27560
rect 25271 27588 25283 27591
rect 25406 27588 25412 27600
rect 25271 27560 25412 27588
rect 25271 27557 25283 27560
rect 25225 27551 25283 27557
rect 25406 27548 25412 27560
rect 25464 27588 25470 27600
rect 26878 27588 26884 27600
rect 25464 27560 26884 27588
rect 25464 27548 25470 27560
rect 26878 27548 26884 27560
rect 26936 27548 26942 27600
rect 29822 27588 29828 27600
rect 29656 27560 29828 27588
rect 7193 27523 7251 27529
rect 7193 27520 7205 27523
rect 6696 27492 7205 27520
rect 6696 27480 6702 27492
rect 7193 27489 7205 27492
rect 7239 27489 7251 27523
rect 7193 27483 7251 27489
rect 7282 27480 7288 27532
rect 7340 27520 7346 27532
rect 7449 27523 7507 27529
rect 7449 27520 7461 27523
rect 7340 27492 7461 27520
rect 7340 27480 7346 27492
rect 7449 27489 7461 27492
rect 7495 27489 7507 27523
rect 9950 27520 9956 27532
rect 9911 27492 9956 27520
rect 7449 27483 7507 27489
rect 9950 27480 9956 27492
rect 10008 27480 10014 27532
rect 11054 27520 11060 27532
rect 11015 27492 11060 27520
rect 11054 27480 11060 27492
rect 11112 27480 11118 27532
rect 11324 27523 11382 27529
rect 11324 27489 11336 27523
rect 11370 27520 11382 27523
rect 11790 27520 11796 27532
rect 11370 27492 11796 27520
rect 11370 27489 11382 27492
rect 11324 27483 11382 27489
rect 11790 27480 11796 27492
rect 11848 27520 11854 27532
rect 12342 27520 12348 27532
rect 11848 27492 12348 27520
rect 11848 27480 11854 27492
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 12434 27480 12440 27532
rect 12492 27520 12498 27532
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 12492 27492 13277 27520
rect 12492 27480 12498 27492
rect 13265 27489 13277 27492
rect 13311 27520 13323 27523
rect 13446 27520 13452 27532
rect 13311 27492 13452 27520
rect 13311 27489 13323 27492
rect 13265 27483 13323 27489
rect 13446 27480 13452 27492
rect 13504 27480 13510 27532
rect 16482 27520 16488 27532
rect 16443 27492 16488 27520
rect 16482 27480 16488 27492
rect 16540 27480 16546 27532
rect 19334 27480 19340 27532
rect 19392 27520 19398 27532
rect 19613 27523 19671 27529
rect 19613 27520 19625 27523
rect 19392 27492 19625 27520
rect 19392 27480 19398 27492
rect 19613 27489 19625 27492
rect 19659 27489 19671 27523
rect 22830 27520 22836 27532
rect 22791 27492 22836 27520
rect 19613 27483 19671 27489
rect 22830 27480 22836 27492
rect 22888 27480 22894 27532
rect 29454 27480 29460 27532
rect 29512 27520 29518 27532
rect 29656 27529 29684 27560
rect 29822 27548 29828 27560
rect 29880 27548 29886 27600
rect 31941 27591 31999 27597
rect 31941 27557 31953 27591
rect 31987 27588 31999 27591
rect 32490 27588 32496 27600
rect 31987 27560 32496 27588
rect 31987 27557 31999 27560
rect 31941 27551 31999 27557
rect 32490 27548 32496 27560
rect 32548 27548 32554 27600
rect 32766 27548 32772 27600
rect 32824 27548 32830 27600
rect 34606 27548 34612 27600
rect 34664 27588 34670 27600
rect 35342 27588 35348 27600
rect 34664 27560 35348 27588
rect 34664 27548 34670 27560
rect 35342 27548 35348 27560
rect 35400 27548 35406 27600
rect 35894 27548 35900 27600
rect 35952 27588 35958 27600
rect 36998 27588 37004 27600
rect 35952 27560 37004 27588
rect 35952 27548 35958 27560
rect 36998 27548 37004 27560
rect 37056 27548 37062 27600
rect 29549 27523 29607 27529
rect 29549 27520 29561 27523
rect 29512 27492 29561 27520
rect 29512 27480 29518 27492
rect 29549 27489 29561 27492
rect 29595 27520 29607 27523
rect 29641 27523 29699 27529
rect 29641 27520 29653 27523
rect 29595 27492 29653 27520
rect 29595 27489 29607 27492
rect 29549 27483 29607 27489
rect 29641 27489 29653 27492
rect 29687 27489 29699 27523
rect 29641 27483 29699 27489
rect 29908 27523 29966 27529
rect 29908 27489 29920 27523
rect 29954 27520 29966 27523
rect 30834 27520 30840 27532
rect 29954 27492 30840 27520
rect 29954 27489 29966 27492
rect 29908 27483 29966 27489
rect 30834 27480 30840 27492
rect 30892 27480 30898 27532
rect 31573 27523 31631 27529
rect 31573 27489 31585 27523
rect 31619 27520 31631 27523
rect 32784 27520 32812 27548
rect 31619 27492 32812 27520
rect 34057 27523 34115 27529
rect 31619 27489 31631 27492
rect 31573 27483 31631 27489
rect 34057 27489 34069 27523
rect 34103 27520 34115 27523
rect 34422 27520 34428 27532
rect 34103 27492 34428 27520
rect 34103 27489 34115 27492
rect 34057 27483 34115 27489
rect 34422 27480 34428 27492
rect 34480 27480 34486 27532
rect 35428 27523 35486 27529
rect 35428 27489 35440 27523
rect 35474 27520 35486 27523
rect 36354 27520 36360 27532
rect 35474 27492 36360 27520
rect 35474 27489 35486 27492
rect 35428 27483 35486 27489
rect 36354 27480 36360 27492
rect 36412 27480 36418 27532
rect 19058 27412 19064 27464
rect 19116 27452 19122 27464
rect 19705 27455 19763 27461
rect 19705 27452 19717 27455
rect 19116 27424 19717 27452
rect 19116 27412 19122 27424
rect 19705 27421 19717 27424
rect 19751 27421 19763 27455
rect 19886 27452 19892 27464
rect 19847 27424 19892 27452
rect 19705 27415 19763 27421
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 20717 27455 20775 27461
rect 20717 27421 20729 27455
rect 20763 27452 20775 27455
rect 21361 27455 21419 27461
rect 21361 27452 21373 27455
rect 20763 27424 21373 27452
rect 20763 27421 20775 27424
rect 20717 27415 20775 27421
rect 21361 27421 21373 27424
rect 21407 27421 21419 27455
rect 21361 27415 21419 27421
rect 21545 27455 21603 27461
rect 21545 27421 21557 27455
rect 21591 27452 21603 27455
rect 22094 27452 22100 27464
rect 21591 27424 22100 27452
rect 21591 27421 21603 27424
rect 21545 27415 21603 27421
rect 10134 27384 10140 27396
rect 10095 27356 10140 27384
rect 10134 27344 10140 27356
rect 10192 27344 10198 27396
rect 13449 27387 13507 27393
rect 13449 27353 13461 27387
rect 13495 27384 13507 27387
rect 13722 27384 13728 27396
rect 13495 27356 13728 27384
rect 13495 27353 13507 27356
rect 13449 27347 13507 27353
rect 13722 27344 13728 27356
rect 13780 27344 13786 27396
rect 18966 27344 18972 27396
rect 19024 27384 19030 27396
rect 19245 27387 19303 27393
rect 19245 27384 19257 27387
rect 19024 27356 19257 27384
rect 19024 27344 19030 27356
rect 19245 27353 19257 27356
rect 19291 27353 19303 27387
rect 19245 27347 19303 27353
rect 20901 27387 20959 27393
rect 20901 27353 20913 27387
rect 20947 27384 20959 27387
rect 21082 27384 21088 27396
rect 20947 27356 21088 27384
rect 20947 27353 20959 27356
rect 20901 27347 20959 27353
rect 21082 27344 21088 27356
rect 21140 27344 21146 27396
rect 21376 27384 21404 27415
rect 22094 27412 22100 27424
rect 22152 27412 22158 27464
rect 22646 27412 22652 27464
rect 22704 27452 22710 27464
rect 22925 27455 22983 27461
rect 22925 27452 22937 27455
rect 22704 27424 22937 27452
rect 22704 27412 22710 27424
rect 22925 27421 22937 27424
rect 22971 27421 22983 27455
rect 23106 27452 23112 27464
rect 23067 27424 23112 27452
rect 22925 27415 22983 27421
rect 23106 27412 23112 27424
rect 23164 27412 23170 27464
rect 25314 27452 25320 27464
rect 25275 27424 25320 27452
rect 25314 27412 25320 27424
rect 25372 27412 25378 27464
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27452 25467 27455
rect 25590 27452 25596 27464
rect 25455 27424 25596 27452
rect 25455 27421 25467 27424
rect 25409 27415 25467 27421
rect 22465 27387 22523 27393
rect 22465 27384 22477 27387
rect 21376 27356 22477 27384
rect 22465 27353 22477 27356
rect 22511 27353 22523 27387
rect 22465 27347 22523 27353
rect 24765 27387 24823 27393
rect 24765 27353 24777 27387
rect 24811 27384 24823 27387
rect 25424 27384 25452 27415
rect 25590 27412 25596 27424
rect 25648 27412 25654 27464
rect 26510 27452 26516 27464
rect 26471 27424 26516 27452
rect 26510 27412 26516 27424
rect 26568 27412 26574 27464
rect 32769 27455 32827 27461
rect 32769 27421 32781 27455
rect 32815 27452 32827 27455
rect 33502 27452 33508 27464
rect 32815 27424 33508 27452
rect 32815 27421 32827 27424
rect 32769 27415 32827 27421
rect 33502 27412 33508 27424
rect 33560 27412 33566 27464
rect 34698 27412 34704 27464
rect 34756 27452 34762 27464
rect 35161 27455 35219 27461
rect 35161 27452 35173 27455
rect 34756 27424 35173 27452
rect 34756 27412 34762 27424
rect 35161 27421 35173 27424
rect 35207 27421 35219 27455
rect 35161 27415 35219 27421
rect 24811 27356 25452 27384
rect 33520 27384 33548 27412
rect 34609 27387 34667 27393
rect 34609 27384 34621 27387
rect 33520 27356 34621 27384
rect 24811 27353 24823 27356
rect 24765 27347 24823 27353
rect 34609 27353 34621 27356
rect 34655 27353 34667 27387
rect 34609 27347 34667 27353
rect 12342 27276 12348 27328
rect 12400 27316 12406 27328
rect 12437 27319 12495 27325
rect 12437 27316 12449 27319
rect 12400 27288 12449 27316
rect 12400 27276 12406 27288
rect 12437 27285 12449 27288
rect 12483 27285 12495 27319
rect 12437 27279 12495 27285
rect 12805 27319 12863 27325
rect 12805 27285 12817 27319
rect 12851 27316 12863 27319
rect 12894 27316 12900 27328
rect 12851 27288 12900 27316
rect 12851 27285 12863 27288
rect 12805 27279 12863 27285
rect 12894 27276 12900 27288
rect 12952 27276 12958 27328
rect 15378 27276 15384 27328
rect 15436 27316 15442 27328
rect 16209 27319 16267 27325
rect 16209 27316 16221 27319
rect 15436 27288 16221 27316
rect 15436 27276 15442 27288
rect 16209 27285 16221 27288
rect 16255 27285 16267 27319
rect 16666 27316 16672 27328
rect 16627 27288 16672 27316
rect 16209 27279 16267 27285
rect 16666 27276 16672 27288
rect 16724 27276 16730 27328
rect 20349 27319 20407 27325
rect 20349 27285 20361 27319
rect 20395 27316 20407 27319
rect 20990 27316 20996 27328
rect 20395 27288 20996 27316
rect 20395 27285 20407 27288
rect 20349 27279 20407 27285
rect 20990 27276 20996 27288
rect 21048 27276 21054 27328
rect 25590 27276 25596 27328
rect 25648 27316 25654 27328
rect 25869 27319 25927 27325
rect 25869 27316 25881 27319
rect 25648 27288 25881 27316
rect 25648 27276 25654 27288
rect 25869 27285 25881 27288
rect 25915 27316 25927 27319
rect 26973 27319 27031 27325
rect 26973 27316 26985 27319
rect 25915 27288 26985 27316
rect 25915 27285 25927 27288
rect 25869 27279 25927 27285
rect 26973 27285 26985 27288
rect 27019 27316 27031 27319
rect 27798 27316 27804 27328
rect 27019 27288 27804 27316
rect 27019 27285 27031 27288
rect 26973 27279 27031 27285
rect 27798 27276 27804 27288
rect 27856 27276 27862 27328
rect 32122 27316 32128 27328
rect 32083 27288 32128 27316
rect 32122 27276 32128 27288
rect 32180 27276 32186 27328
rect 33226 27316 33232 27328
rect 33187 27288 33232 27316
rect 33226 27276 33232 27288
rect 33284 27276 33290 27328
rect 34238 27316 34244 27328
rect 34199 27288 34244 27316
rect 34238 27276 34244 27288
rect 34296 27276 34302 27328
rect 36541 27319 36599 27325
rect 36541 27285 36553 27319
rect 36587 27316 36599 27319
rect 36814 27316 36820 27328
rect 36587 27288 36820 27316
rect 36587 27285 36599 27288
rect 36541 27279 36599 27285
rect 36814 27276 36820 27288
rect 36872 27276 36878 27328
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 2038 27112 2044 27124
rect 1999 27084 2044 27112
rect 2038 27072 2044 27084
rect 2096 27072 2102 27124
rect 6638 27112 6644 27124
rect 6599 27084 6644 27112
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 7742 27112 7748 27124
rect 7703 27084 7748 27112
rect 7742 27072 7748 27084
rect 7800 27072 7806 27124
rect 8202 27112 8208 27124
rect 8163 27084 8208 27112
rect 8202 27072 8208 27084
rect 8260 27072 8266 27124
rect 9950 27112 9956 27124
rect 9911 27084 9956 27112
rect 9950 27072 9956 27084
rect 10008 27112 10014 27124
rect 10689 27115 10747 27121
rect 10689 27112 10701 27115
rect 10008 27084 10701 27112
rect 10008 27072 10014 27084
rect 10689 27081 10701 27084
rect 10735 27081 10747 27115
rect 11790 27112 11796 27124
rect 11751 27084 11796 27112
rect 10689 27075 10747 27081
rect 11790 27072 11796 27084
rect 11848 27072 11854 27124
rect 12250 27072 12256 27124
rect 12308 27112 12314 27124
rect 12437 27115 12495 27121
rect 12437 27112 12449 27115
rect 12308 27084 12449 27112
rect 12308 27072 12314 27084
rect 12437 27081 12449 27084
rect 12483 27081 12495 27115
rect 13446 27112 13452 27124
rect 13407 27084 13452 27112
rect 12437 27075 12495 27081
rect 13446 27072 13452 27084
rect 13504 27072 13510 27124
rect 15286 27112 15292 27124
rect 15247 27084 15292 27112
rect 15286 27072 15292 27084
rect 15344 27072 15350 27124
rect 16482 27072 16488 27124
rect 16540 27112 16546 27124
rect 17129 27115 17187 27121
rect 17129 27112 17141 27115
rect 16540 27084 17141 27112
rect 16540 27072 16546 27084
rect 17129 27081 17141 27084
rect 17175 27112 17187 27115
rect 18506 27112 18512 27124
rect 17175 27084 18512 27112
rect 17175 27081 17187 27084
rect 17129 27075 17187 27081
rect 18506 27072 18512 27084
rect 18564 27072 18570 27124
rect 18969 27115 19027 27121
rect 18969 27081 18981 27115
rect 19015 27112 19027 27115
rect 19058 27112 19064 27124
rect 19015 27084 19064 27112
rect 19015 27081 19027 27084
rect 18969 27075 19027 27081
rect 19058 27072 19064 27084
rect 19116 27072 19122 27124
rect 19334 27112 19340 27124
rect 19295 27084 19340 27112
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 20349 27115 20407 27121
rect 20349 27081 20361 27115
rect 20395 27112 20407 27115
rect 21174 27112 21180 27124
rect 20395 27084 21180 27112
rect 20395 27081 20407 27084
rect 20349 27075 20407 27081
rect 21174 27072 21180 27084
rect 21232 27072 21238 27124
rect 21818 27112 21824 27124
rect 21779 27084 21824 27112
rect 21818 27072 21824 27084
rect 21876 27112 21882 27124
rect 23106 27112 23112 27124
rect 21876 27084 23112 27112
rect 21876 27072 21882 27084
rect 23106 27072 23112 27084
rect 23164 27112 23170 27124
rect 23201 27115 23259 27121
rect 23201 27112 23213 27115
rect 23164 27084 23213 27112
rect 23164 27072 23170 27084
rect 23201 27081 23213 27084
rect 23247 27081 23259 27115
rect 25406 27112 25412 27124
rect 25367 27084 25412 27112
rect 23201 27075 23259 27081
rect 25406 27072 25412 27084
rect 25464 27072 25470 27124
rect 27798 27112 27804 27124
rect 27759 27084 27804 27112
rect 27798 27072 27804 27084
rect 27856 27072 27862 27124
rect 30834 27112 30840 27124
rect 30795 27084 30840 27112
rect 30834 27072 30840 27084
rect 30892 27112 30898 27124
rect 31113 27115 31171 27121
rect 31113 27112 31125 27115
rect 30892 27084 31125 27112
rect 30892 27072 30898 27084
rect 31113 27081 31125 27084
rect 31159 27112 31171 27115
rect 31481 27115 31539 27121
rect 31481 27112 31493 27115
rect 31159 27084 31493 27112
rect 31159 27081 31171 27084
rect 31113 27075 31171 27081
rect 31481 27081 31493 27084
rect 31527 27081 31539 27115
rect 31662 27112 31668 27124
rect 31623 27084 31668 27112
rect 31481 27075 31539 27081
rect 12894 27004 12900 27056
rect 12952 27044 12958 27056
rect 12952 27016 13032 27044
rect 12952 27004 12958 27016
rect 8846 26976 8852 26988
rect 8807 26948 8852 26976
rect 8846 26936 8852 26948
rect 8904 26936 8910 26988
rect 11330 26976 11336 26988
rect 11291 26948 11336 26976
rect 11330 26936 11336 26948
rect 11388 26936 11394 26988
rect 12342 26936 12348 26988
rect 12400 26936 12406 26988
rect 13004 26985 13032 27016
rect 12989 26979 13047 26985
rect 12989 26945 13001 26979
rect 13035 26945 13047 26979
rect 15304 26976 15332 27072
rect 19352 26976 19380 27072
rect 22094 27004 22100 27056
rect 22152 27044 22158 27056
rect 22152 27016 22197 27044
rect 22152 27004 22158 27016
rect 19429 26979 19487 26985
rect 19429 26976 19441 26979
rect 15304 26948 15516 26976
rect 19352 26948 19441 26976
rect 12989 26939 13047 26945
rect 7742 26868 7748 26920
rect 7800 26908 7806 26920
rect 8573 26911 8631 26917
rect 8573 26908 8585 26911
rect 7800 26880 8585 26908
rect 7800 26868 7806 26880
rect 8573 26877 8585 26880
rect 8619 26877 8631 26911
rect 8573 26871 8631 26877
rect 9677 26911 9735 26917
rect 9677 26877 9689 26911
rect 9723 26908 9735 26911
rect 10962 26908 10968 26920
rect 9723 26880 10968 26908
rect 9723 26877 9735 26880
rect 9677 26871 9735 26877
rect 10962 26868 10968 26880
rect 11020 26868 11026 26920
rect 11790 26868 11796 26920
rect 11848 26908 11854 26920
rect 12360 26908 12388 26936
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 11848 26880 12909 26908
rect 11848 26868 11854 26880
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 12897 26871 12955 26877
rect 14369 26911 14427 26917
rect 14369 26877 14381 26911
rect 14415 26908 14427 26911
rect 14415 26880 14780 26908
rect 14415 26877 14427 26880
rect 14369 26871 14427 26877
rect 1670 26840 1676 26852
rect 1583 26812 1676 26840
rect 1670 26800 1676 26812
rect 1728 26840 1734 26852
rect 2682 26840 2688 26852
rect 1728 26812 2688 26840
rect 1728 26800 1734 26812
rect 2682 26800 2688 26812
rect 2740 26800 2746 26852
rect 8665 26843 8723 26849
rect 8665 26840 8677 26843
rect 8036 26812 8677 26840
rect 7282 26772 7288 26784
rect 7243 26744 7288 26772
rect 7282 26732 7288 26744
rect 7340 26732 7346 26784
rect 7834 26732 7840 26784
rect 7892 26772 7898 26784
rect 8036 26781 8064 26812
rect 8665 26809 8677 26812
rect 8711 26809 8723 26843
rect 8665 26803 8723 26809
rect 10597 26843 10655 26849
rect 10597 26809 10609 26843
rect 10643 26840 10655 26843
rect 11149 26843 11207 26849
rect 11149 26840 11161 26843
rect 10643 26812 11161 26840
rect 10643 26809 10655 26812
rect 10597 26803 10655 26809
rect 11149 26809 11161 26812
rect 11195 26840 11207 26843
rect 12342 26840 12348 26852
rect 11195 26812 12348 26840
rect 11195 26809 11207 26812
rect 11149 26803 11207 26809
rect 12342 26800 12348 26812
rect 12400 26800 12406 26852
rect 14752 26784 14780 26880
rect 15286 26868 15292 26920
rect 15344 26908 15350 26920
rect 15381 26911 15439 26917
rect 15381 26908 15393 26911
rect 15344 26880 15393 26908
rect 15344 26868 15350 26880
rect 15381 26877 15393 26880
rect 15427 26877 15439 26911
rect 15488 26908 15516 26948
rect 19429 26945 19441 26948
rect 19475 26945 19487 26979
rect 24578 26976 24584 26988
rect 24539 26948 24584 26976
rect 19429 26939 19487 26945
rect 24578 26936 24584 26948
rect 24636 26936 24642 26988
rect 28721 26979 28779 26985
rect 28721 26945 28733 26979
rect 28767 26976 28779 26979
rect 31496 26976 31524 27075
rect 31662 27072 31668 27084
rect 31720 27072 31726 27124
rect 32306 27072 32312 27124
rect 32364 27112 32370 27124
rect 32677 27115 32735 27121
rect 32677 27112 32689 27115
rect 32364 27084 32689 27112
rect 32364 27072 32370 27084
rect 32677 27081 32689 27084
rect 32723 27081 32735 27115
rect 32677 27075 32735 27081
rect 34333 27115 34391 27121
rect 34333 27081 34345 27115
rect 34379 27112 34391 27115
rect 34422 27112 34428 27124
rect 34379 27084 34428 27112
rect 34379 27081 34391 27084
rect 34333 27075 34391 27081
rect 34422 27072 34428 27084
rect 34480 27072 34486 27124
rect 34701 27115 34759 27121
rect 34701 27081 34713 27115
rect 34747 27112 34759 27115
rect 34790 27112 34796 27124
rect 34747 27084 34796 27112
rect 34747 27081 34759 27084
rect 34701 27075 34759 27081
rect 34790 27072 34796 27084
rect 34848 27112 34854 27124
rect 35989 27115 36047 27121
rect 34848 27084 35388 27112
rect 34848 27072 34854 27084
rect 32125 26979 32183 26985
rect 32125 26976 32137 26979
rect 28767 26948 29408 26976
rect 31496 26948 32137 26976
rect 28767 26945 28779 26948
rect 28721 26939 28779 26945
rect 15637 26911 15695 26917
rect 15637 26908 15649 26911
rect 15488 26880 15649 26908
rect 15381 26871 15439 26877
rect 15637 26877 15649 26880
rect 15683 26877 15695 26911
rect 15637 26871 15695 26877
rect 20441 26911 20499 26917
rect 20441 26877 20453 26911
rect 20487 26908 20499 26911
rect 20990 26908 20996 26920
rect 20487 26880 20996 26908
rect 20487 26877 20499 26880
rect 20441 26871 20499 26877
rect 20990 26868 20996 26880
rect 21048 26868 21054 26920
rect 24489 26911 24547 26917
rect 24489 26877 24501 26911
rect 24535 26908 24547 26911
rect 25406 26908 25412 26920
rect 24535 26880 25412 26908
rect 24535 26877 24547 26880
rect 24489 26871 24547 26877
rect 25406 26868 25412 26880
rect 25464 26868 25470 26920
rect 25590 26908 25596 26920
rect 25551 26880 25596 26908
rect 25590 26868 25596 26880
rect 25648 26868 25654 26920
rect 27706 26868 27712 26920
rect 27764 26908 27770 26920
rect 27985 26911 28043 26917
rect 27985 26908 27997 26911
rect 27764 26880 27997 26908
rect 27764 26868 27770 26880
rect 27985 26877 27997 26880
rect 28031 26908 28043 26911
rect 28261 26911 28319 26917
rect 28261 26908 28273 26911
rect 28031 26880 28273 26908
rect 28031 26877 28043 26880
rect 27985 26871 28043 26877
rect 28261 26877 28273 26880
rect 28307 26877 28319 26911
rect 29380 26908 29408 26948
rect 32125 26945 32137 26948
rect 32171 26945 32183 26979
rect 32125 26939 32183 26945
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26976 32367 26979
rect 32766 26976 32772 26988
rect 32355 26948 32772 26976
rect 32355 26945 32367 26948
rect 32309 26939 32367 26945
rect 32766 26936 32772 26948
rect 32824 26936 32830 26988
rect 33502 26936 33508 26988
rect 33560 26976 33566 26988
rect 35360 26985 35388 27084
rect 35989 27081 36001 27115
rect 36035 27112 36047 27115
rect 36354 27112 36360 27124
rect 36035 27084 36360 27112
rect 36035 27081 36047 27084
rect 35989 27075 36047 27081
rect 36354 27072 36360 27084
rect 36412 27072 36418 27124
rect 37458 27112 37464 27124
rect 37419 27084 37464 27112
rect 37458 27072 37464 27084
rect 37516 27072 37522 27124
rect 33781 26979 33839 26985
rect 33781 26976 33793 26979
rect 33560 26948 33793 26976
rect 33560 26936 33566 26948
rect 33781 26945 33793 26948
rect 33827 26945 33839 26979
rect 33781 26939 33839 26945
rect 35345 26979 35403 26985
rect 35345 26945 35357 26979
rect 35391 26945 35403 26979
rect 35345 26939 35403 26945
rect 35437 26979 35495 26985
rect 35437 26945 35449 26979
rect 35483 26976 35495 26979
rect 36630 26976 36636 26988
rect 35483 26948 36636 26976
rect 35483 26945 35495 26948
rect 35437 26939 35495 26945
rect 29457 26911 29515 26917
rect 29457 26908 29469 26911
rect 29380 26880 29469 26908
rect 28261 26871 28319 26877
rect 29457 26877 29469 26880
rect 29503 26908 29515 26911
rect 29546 26908 29552 26920
rect 29503 26880 29552 26908
rect 29503 26877 29515 26880
rect 29457 26871 29515 26877
rect 29546 26868 29552 26880
rect 29604 26868 29610 26920
rect 33226 26868 33232 26920
rect 33284 26908 33290 26920
rect 33597 26911 33655 26917
rect 33597 26908 33609 26911
rect 33284 26880 33609 26908
rect 33284 26868 33290 26880
rect 33597 26877 33609 26880
rect 33643 26877 33655 26911
rect 33597 26871 33655 26877
rect 19886 26800 19892 26852
rect 19944 26840 19950 26852
rect 20714 26849 20720 26852
rect 19981 26843 20039 26849
rect 19981 26840 19993 26843
rect 19944 26812 19993 26840
rect 19944 26800 19950 26812
rect 19981 26809 19993 26812
rect 20027 26840 20039 26843
rect 20708 26840 20720 26849
rect 20027 26812 20720 26840
rect 20027 26809 20039 26812
rect 19981 26803 20039 26809
rect 20708 26803 20720 26812
rect 20714 26800 20720 26803
rect 20772 26800 20778 26852
rect 22094 26800 22100 26852
rect 22152 26840 22158 26852
rect 22830 26840 22836 26852
rect 22152 26812 22836 26840
rect 22152 26800 22158 26812
rect 22830 26800 22836 26812
rect 22888 26800 22894 26852
rect 23937 26843 23995 26849
rect 23937 26809 23949 26843
rect 23983 26840 23995 26843
rect 25133 26843 25191 26849
rect 23983 26812 24440 26840
rect 23983 26809 23995 26812
rect 23937 26803 23995 26809
rect 8021 26775 8079 26781
rect 8021 26772 8033 26775
rect 7892 26744 8033 26772
rect 7892 26732 7898 26744
rect 8021 26741 8033 26744
rect 8067 26741 8079 26775
rect 11054 26772 11060 26784
rect 11015 26744 11060 26772
rect 8021 26735 8079 26741
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 11790 26732 11796 26784
rect 11848 26772 11854 26784
rect 12161 26775 12219 26781
rect 12161 26772 12173 26775
rect 11848 26744 12173 26772
rect 11848 26732 11854 26744
rect 12161 26741 12173 26744
rect 12207 26741 12219 26775
rect 12161 26735 12219 26741
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 12805 26775 12863 26781
rect 12805 26772 12817 26775
rect 12584 26744 12817 26772
rect 12584 26732 12590 26744
rect 12805 26741 12817 26744
rect 12851 26741 12863 26775
rect 12805 26735 12863 26741
rect 13998 26732 14004 26784
rect 14056 26772 14062 26784
rect 14185 26775 14243 26781
rect 14185 26772 14197 26775
rect 14056 26744 14197 26772
rect 14056 26732 14062 26744
rect 14185 26741 14197 26744
rect 14231 26741 14243 26775
rect 14734 26772 14740 26784
rect 14695 26744 14740 26772
rect 14185 26735 14243 26741
rect 14734 26732 14740 26744
rect 14792 26732 14798 26784
rect 15930 26732 15936 26784
rect 15988 26772 15994 26784
rect 16761 26775 16819 26781
rect 16761 26772 16773 26775
rect 15988 26744 16773 26772
rect 15988 26732 15994 26744
rect 16761 26741 16773 26744
rect 16807 26741 16819 26775
rect 16761 26735 16819 26741
rect 22557 26775 22615 26781
rect 22557 26741 22569 26775
rect 22603 26772 22615 26775
rect 22646 26772 22652 26784
rect 22603 26744 22652 26772
rect 22603 26741 22615 26744
rect 22557 26735 22615 26741
rect 22646 26732 22652 26744
rect 22704 26772 22710 26784
rect 23952 26772 23980 26803
rect 24412 26784 24440 26812
rect 25133 26809 25145 26843
rect 25179 26840 25191 26843
rect 25314 26840 25320 26852
rect 25179 26812 25320 26840
rect 25179 26809 25191 26812
rect 25133 26803 25191 26809
rect 25314 26800 25320 26812
rect 25372 26840 25378 26852
rect 25866 26849 25872 26852
rect 25372 26812 25820 26840
rect 25372 26800 25378 26812
rect 22704 26744 23980 26772
rect 22704 26732 22710 26744
rect 24026 26732 24032 26784
rect 24084 26772 24090 26784
rect 24394 26772 24400 26784
rect 24084 26744 24129 26772
rect 24355 26744 24400 26772
rect 24084 26732 24090 26744
rect 24394 26732 24400 26744
rect 24452 26732 24458 26784
rect 25792 26772 25820 26812
rect 25860 26803 25872 26849
rect 25924 26840 25930 26852
rect 29089 26843 29147 26849
rect 25924 26812 25960 26840
rect 25866 26800 25872 26803
rect 25924 26800 25930 26812
rect 29089 26809 29101 26843
rect 29135 26840 29147 26843
rect 29702 26843 29760 26849
rect 29702 26840 29714 26843
rect 29135 26812 29714 26840
rect 29135 26809 29147 26812
rect 29089 26803 29147 26809
rect 29702 26809 29714 26812
rect 29748 26840 29760 26843
rect 30834 26840 30840 26852
rect 29748 26812 30840 26840
rect 29748 26809 29760 26812
rect 29702 26803 29760 26809
rect 30834 26800 30840 26812
rect 30892 26800 30898 26852
rect 33689 26843 33747 26849
rect 33689 26840 33701 26843
rect 33060 26812 33701 26840
rect 33060 26784 33088 26812
rect 33689 26809 33701 26812
rect 33735 26809 33747 26843
rect 33796 26840 33824 26939
rect 35452 26908 35480 26939
rect 36630 26936 36636 26948
rect 36688 26936 36694 26988
rect 36998 26976 37004 26988
rect 36959 26948 37004 26976
rect 36998 26936 37004 26948
rect 37056 26936 37062 26988
rect 34900 26880 35480 26908
rect 34900 26840 34928 26880
rect 36354 26868 36360 26920
rect 36412 26908 36418 26920
rect 36909 26911 36967 26917
rect 36909 26908 36921 26911
rect 36412 26880 36921 26908
rect 36412 26868 36418 26880
rect 36909 26877 36921 26880
rect 36955 26877 36967 26911
rect 36909 26871 36967 26877
rect 33796 26812 34928 26840
rect 33689 26803 33747 26809
rect 34974 26800 34980 26852
rect 35032 26840 35038 26852
rect 35253 26843 35311 26849
rect 35253 26840 35265 26843
rect 35032 26812 35265 26840
rect 35032 26800 35038 26812
rect 35253 26809 35265 26812
rect 35299 26840 35311 26843
rect 35299 26812 36492 26840
rect 35299 26809 35311 26812
rect 35253 26803 35311 26809
rect 25958 26772 25964 26784
rect 25792 26744 25964 26772
rect 25958 26732 25964 26744
rect 26016 26732 26022 26784
rect 26050 26732 26056 26784
rect 26108 26772 26114 26784
rect 26973 26775 27031 26781
rect 26973 26772 26985 26775
rect 26108 26744 26985 26772
rect 26108 26732 26114 26744
rect 26973 26741 26985 26744
rect 27019 26741 27031 26775
rect 32030 26772 32036 26784
rect 31991 26744 32036 26772
rect 26973 26735 27031 26741
rect 32030 26732 32036 26744
rect 32088 26732 32094 26784
rect 33042 26772 33048 26784
rect 33003 26744 33048 26772
rect 33042 26732 33048 26744
rect 33100 26732 33106 26784
rect 33226 26772 33232 26784
rect 33187 26744 33232 26772
rect 33226 26732 33232 26744
rect 33284 26732 33290 26784
rect 34422 26732 34428 26784
rect 34480 26772 34486 26784
rect 36464 26781 36492 26812
rect 34885 26775 34943 26781
rect 34885 26772 34897 26775
rect 34480 26744 34897 26772
rect 34480 26732 34486 26744
rect 34885 26741 34897 26744
rect 34931 26741 34943 26775
rect 34885 26735 34943 26741
rect 36449 26775 36507 26781
rect 36449 26741 36461 26775
rect 36495 26741 36507 26775
rect 36814 26772 36820 26784
rect 36775 26744 36820 26772
rect 36449 26735 36507 26741
rect 36814 26732 36820 26744
rect 36872 26732 36878 26784
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 7282 26528 7288 26580
rect 7340 26568 7346 26580
rect 8297 26571 8355 26577
rect 8297 26568 8309 26571
rect 7340 26540 8309 26568
rect 7340 26528 7346 26540
rect 8297 26537 8309 26540
rect 8343 26537 8355 26571
rect 8297 26531 8355 26537
rect 8665 26571 8723 26577
rect 8665 26537 8677 26571
rect 8711 26568 8723 26571
rect 8846 26568 8852 26580
rect 8711 26540 8852 26568
rect 8711 26537 8723 26540
rect 8665 26531 8723 26537
rect 8846 26528 8852 26540
rect 8904 26568 8910 26580
rect 10413 26571 10471 26577
rect 10413 26568 10425 26571
rect 8904 26540 10425 26568
rect 8904 26528 8910 26540
rect 10413 26537 10425 26540
rect 10459 26568 10471 26571
rect 11330 26568 11336 26580
rect 10459 26540 11336 26568
rect 10459 26537 10471 26540
rect 10413 26531 10471 26537
rect 11330 26528 11336 26540
rect 11388 26528 11394 26580
rect 15930 26568 15936 26580
rect 15891 26540 15936 26568
rect 15930 26528 15936 26540
rect 15988 26528 15994 26580
rect 19058 26528 19064 26580
rect 19116 26568 19122 26580
rect 19245 26571 19303 26577
rect 19245 26568 19257 26571
rect 19116 26540 19257 26568
rect 19116 26528 19122 26540
rect 19245 26537 19257 26540
rect 19291 26537 19303 26571
rect 19245 26531 19303 26537
rect 19613 26571 19671 26577
rect 19613 26537 19625 26571
rect 19659 26568 19671 26571
rect 19978 26568 19984 26580
rect 19659 26540 19984 26568
rect 19659 26537 19671 26540
rect 19613 26531 19671 26537
rect 6914 26460 6920 26512
rect 6972 26500 6978 26512
rect 7162 26503 7220 26509
rect 7162 26500 7174 26503
rect 6972 26472 7174 26500
rect 6972 26460 6978 26472
rect 7162 26469 7174 26472
rect 7208 26500 7220 26503
rect 7558 26500 7564 26512
rect 7208 26472 7564 26500
rect 7208 26469 7220 26472
rect 7162 26463 7220 26469
rect 7558 26460 7564 26472
rect 7616 26500 7622 26512
rect 8202 26500 8208 26512
rect 7616 26472 8208 26500
rect 7616 26460 7622 26472
rect 8202 26460 8208 26472
rect 8260 26460 8266 26512
rect 10781 26503 10839 26509
rect 10781 26469 10793 26503
rect 10827 26500 10839 26503
rect 11054 26500 11060 26512
rect 10827 26472 11060 26500
rect 10827 26469 10839 26472
rect 10781 26463 10839 26469
rect 11054 26460 11060 26472
rect 11112 26500 11118 26512
rect 12342 26500 12348 26512
rect 11112 26472 12348 26500
rect 11112 26460 11118 26472
rect 12342 26460 12348 26472
rect 12400 26460 12406 26512
rect 19150 26500 19156 26512
rect 19063 26472 19156 26500
rect 19150 26460 19156 26472
rect 19208 26500 19214 26512
rect 19628 26500 19656 26531
rect 19978 26528 19984 26540
rect 20036 26528 20042 26580
rect 20533 26571 20591 26577
rect 20533 26537 20545 26571
rect 20579 26568 20591 26571
rect 20714 26568 20720 26580
rect 20579 26540 20720 26568
rect 20579 26537 20591 26540
rect 20533 26531 20591 26537
rect 20714 26528 20720 26540
rect 20772 26568 20778 26580
rect 22281 26571 22339 26577
rect 22281 26568 22293 26571
rect 20772 26540 22293 26568
rect 20772 26528 20778 26540
rect 22281 26537 22293 26540
rect 22327 26537 22339 26571
rect 22281 26531 22339 26537
rect 23845 26571 23903 26577
rect 23845 26537 23857 26571
rect 23891 26568 23903 26571
rect 23934 26568 23940 26580
rect 23891 26540 23940 26568
rect 23891 26537 23903 26540
rect 23845 26531 23903 26537
rect 23934 26528 23940 26540
rect 23992 26568 23998 26580
rect 24578 26568 24584 26580
rect 23992 26540 24584 26568
rect 23992 26528 23998 26540
rect 24578 26528 24584 26540
rect 24636 26528 24642 26580
rect 24857 26571 24915 26577
rect 24857 26537 24869 26571
rect 24903 26568 24915 26571
rect 24946 26568 24952 26580
rect 24903 26540 24952 26568
rect 24903 26537 24915 26540
rect 24857 26531 24915 26537
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 25225 26571 25283 26577
rect 25225 26537 25237 26571
rect 25271 26568 25283 26571
rect 26510 26568 26516 26580
rect 25271 26540 26516 26568
rect 25271 26537 25283 26540
rect 25225 26531 25283 26537
rect 19208 26472 19656 26500
rect 24765 26503 24823 26509
rect 19208 26460 19214 26472
rect 24765 26469 24777 26503
rect 24811 26500 24823 26503
rect 25240 26500 25268 26531
rect 26510 26528 26516 26540
rect 26568 26528 26574 26580
rect 30834 26568 30840 26580
rect 30795 26540 30840 26568
rect 30834 26528 30840 26540
rect 30892 26528 30898 26580
rect 31018 26528 31024 26580
rect 31076 26568 31082 26580
rect 31665 26571 31723 26577
rect 31665 26568 31677 26571
rect 31076 26540 31677 26568
rect 31076 26528 31082 26540
rect 31665 26537 31677 26540
rect 31711 26568 31723 26571
rect 32030 26568 32036 26580
rect 31711 26540 32036 26568
rect 31711 26537 31723 26540
rect 31665 26531 31723 26537
rect 32030 26528 32036 26540
rect 32088 26528 32094 26580
rect 32125 26571 32183 26577
rect 32125 26537 32137 26571
rect 32171 26568 32183 26571
rect 33042 26568 33048 26580
rect 32171 26540 33048 26568
rect 32171 26537 32183 26540
rect 32125 26531 32183 26537
rect 33042 26528 33048 26540
rect 33100 26528 33106 26580
rect 34974 26568 34980 26580
rect 34935 26540 34980 26568
rect 34974 26528 34980 26540
rect 35032 26528 35038 26580
rect 24811 26472 25268 26500
rect 30852 26500 30880 26528
rect 32493 26503 32551 26509
rect 32493 26500 32505 26503
rect 30852 26472 32505 26500
rect 24811 26469 24823 26472
rect 24765 26463 24823 26469
rect 32493 26469 32505 26472
rect 32539 26500 32551 26503
rect 32674 26500 32680 26512
rect 32539 26472 32680 26500
rect 32539 26469 32551 26472
rect 32493 26463 32551 26469
rect 32674 26460 32680 26472
rect 32732 26460 32738 26512
rect 33778 26460 33784 26512
rect 33836 26500 33842 26512
rect 34149 26503 34207 26509
rect 34149 26500 34161 26503
rect 33836 26472 34161 26500
rect 33836 26460 33842 26472
rect 34149 26469 34161 26472
rect 34195 26469 34207 26503
rect 34149 26463 34207 26469
rect 7006 26392 7012 26444
rect 7064 26392 7070 26444
rect 11324 26435 11382 26441
rect 11324 26401 11336 26435
rect 11370 26432 11382 26435
rect 11790 26432 11796 26444
rect 11370 26404 11796 26432
rect 11370 26401 11382 26404
rect 11324 26395 11382 26401
rect 11790 26392 11796 26404
rect 11848 26392 11854 26444
rect 15838 26432 15844 26444
rect 15799 26404 15844 26432
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 17034 26432 17040 26444
rect 16995 26404 17040 26432
rect 17034 26392 17040 26404
rect 17092 26392 17098 26444
rect 18785 26435 18843 26441
rect 18785 26401 18797 26435
rect 18831 26432 18843 26435
rect 20714 26432 20720 26444
rect 18831 26404 20720 26432
rect 18831 26401 18843 26404
rect 18785 26395 18843 26401
rect 6917 26367 6975 26373
rect 6917 26333 6929 26367
rect 6963 26364 6975 26367
rect 7024 26364 7052 26392
rect 6963 26336 7052 26364
rect 6963 26333 6975 26336
rect 6917 26327 6975 26333
rect 10962 26324 10968 26376
rect 11020 26364 11026 26376
rect 11057 26367 11115 26373
rect 11057 26364 11069 26367
rect 11020 26336 11069 26364
rect 11020 26324 11026 26336
rect 11057 26333 11069 26336
rect 11103 26333 11115 26367
rect 11057 26327 11115 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26364 15163 26367
rect 15746 26364 15752 26376
rect 15151 26336 15752 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 15746 26324 15752 26336
rect 15804 26364 15810 26376
rect 16117 26367 16175 26373
rect 16117 26364 16129 26367
rect 15804 26336 16129 26364
rect 15804 26324 15810 26336
rect 16117 26333 16129 26336
rect 16163 26364 16175 26367
rect 16666 26364 16672 26376
rect 16163 26336 16672 26364
rect 16163 26333 16175 26336
rect 16117 26327 16175 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 19702 26364 19708 26376
rect 19663 26336 19708 26364
rect 19702 26324 19708 26336
rect 19760 26324 19766 26376
rect 19812 26373 19840 26404
rect 20714 26392 20720 26404
rect 20772 26432 20778 26444
rect 21157 26435 21215 26441
rect 21157 26432 21169 26435
rect 20772 26404 21169 26432
rect 20772 26392 20778 26404
rect 21157 26401 21169 26404
rect 21203 26401 21215 26435
rect 21157 26395 21215 26401
rect 24670 26392 24676 26444
rect 24728 26432 24734 26444
rect 24728 26404 25544 26432
rect 24728 26392 24734 26404
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26333 19855 26367
rect 20898 26364 20904 26376
rect 20859 26336 20904 26364
rect 19797 26327 19855 26333
rect 20898 26324 20904 26336
rect 20956 26324 20962 26376
rect 25314 26364 25320 26376
rect 25275 26336 25320 26364
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 25516 26373 25544 26404
rect 25958 26392 25964 26444
rect 26016 26432 26022 26444
rect 27249 26435 27307 26441
rect 27249 26432 27261 26435
rect 26016 26404 27261 26432
rect 26016 26392 26022 26404
rect 27249 26401 27261 26404
rect 27295 26432 27307 26435
rect 27522 26432 27528 26444
rect 27295 26404 27528 26432
rect 27295 26401 27307 26404
rect 27249 26395 27307 26401
rect 27522 26392 27528 26404
rect 27580 26392 27586 26444
rect 28994 26392 29000 26444
rect 29052 26432 29058 26444
rect 29713 26435 29771 26441
rect 29713 26432 29725 26435
rect 29052 26404 29725 26432
rect 29052 26392 29058 26404
rect 29713 26401 29725 26404
rect 29759 26432 29771 26435
rect 30282 26432 30288 26444
rect 29759 26404 30288 26432
rect 29759 26401 29771 26404
rect 29713 26395 29771 26401
rect 30282 26392 30288 26404
rect 30340 26392 30346 26444
rect 33502 26432 33508 26444
rect 31312 26404 33508 26432
rect 31312 26376 31340 26404
rect 33502 26392 33508 26404
rect 33560 26392 33566 26444
rect 33870 26392 33876 26444
rect 33928 26432 33934 26444
rect 34057 26435 34115 26441
rect 34057 26432 34069 26435
rect 33928 26404 34069 26432
rect 33928 26392 33934 26404
rect 34057 26401 34069 26404
rect 34103 26401 34115 26435
rect 34057 26395 34115 26401
rect 34698 26392 34704 26444
rect 34756 26432 34762 26444
rect 35509 26435 35567 26441
rect 35509 26432 35521 26435
rect 34756 26404 35521 26432
rect 34756 26392 34762 26404
rect 35509 26401 35521 26404
rect 35555 26432 35567 26435
rect 36814 26432 36820 26444
rect 35555 26404 36820 26432
rect 35555 26401 35567 26404
rect 35509 26395 35567 26401
rect 36814 26392 36820 26404
rect 36872 26392 36878 26444
rect 25501 26367 25559 26373
rect 25501 26333 25513 26367
rect 25547 26364 25559 26367
rect 26050 26364 26056 26376
rect 25547 26336 26056 26364
rect 25547 26333 25559 26336
rect 25501 26327 25559 26333
rect 26050 26324 26056 26336
rect 26108 26324 26114 26376
rect 26234 26364 26240 26376
rect 26195 26336 26240 26364
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 26326 26324 26332 26376
rect 26384 26364 26390 26376
rect 26513 26367 26571 26373
rect 26513 26364 26525 26367
rect 26384 26336 26525 26364
rect 26384 26324 26390 26336
rect 26513 26333 26525 26336
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 26694 26324 26700 26376
rect 26752 26364 26758 26376
rect 26836 26367 26894 26373
rect 26836 26364 26848 26367
rect 26752 26336 26848 26364
rect 26752 26324 26758 26336
rect 26836 26333 26848 26336
rect 26882 26333 26894 26367
rect 26836 26327 26894 26333
rect 26970 26324 26976 26376
rect 27028 26364 27034 26376
rect 29365 26367 29423 26373
rect 29365 26364 29377 26367
rect 27028 26336 27073 26364
rect 29012 26336 29377 26364
rect 27028 26324 27034 26336
rect 12437 26299 12495 26305
rect 12437 26265 12449 26299
rect 12483 26296 12495 26299
rect 12526 26296 12532 26308
rect 12483 26268 12532 26296
rect 12483 26265 12495 26268
rect 12437 26259 12495 26265
rect 12526 26256 12532 26268
rect 12584 26296 12590 26308
rect 12713 26299 12771 26305
rect 12713 26296 12725 26299
rect 12584 26268 12725 26296
rect 12584 26256 12590 26268
rect 12713 26265 12725 26268
rect 12759 26265 12771 26299
rect 15473 26299 15531 26305
rect 15473 26296 15485 26299
rect 12713 26259 12771 26265
rect 15120 26268 15485 26296
rect 15120 26240 15148 26268
rect 15473 26265 15485 26268
rect 15519 26265 15531 26299
rect 17218 26296 17224 26308
rect 17179 26268 17224 26296
rect 15473 26259 15531 26265
rect 17218 26256 17224 26268
rect 17276 26256 17282 26308
rect 24213 26299 24271 26305
rect 24213 26265 24225 26299
rect 24259 26296 24271 26299
rect 24394 26296 24400 26308
rect 24259 26268 24400 26296
rect 24259 26265 24271 26268
rect 24213 26259 24271 26265
rect 24394 26256 24400 26268
rect 24452 26296 24458 26308
rect 24452 26268 24808 26296
rect 24452 26256 24458 26268
rect 15102 26188 15108 26240
rect 15160 26188 15166 26240
rect 24780 26228 24808 26268
rect 25866 26256 25872 26308
rect 25924 26296 25930 26308
rect 25961 26299 26019 26305
rect 25961 26296 25973 26299
rect 25924 26268 25973 26296
rect 25924 26256 25930 26268
rect 25961 26265 25973 26268
rect 26007 26296 26019 26299
rect 28353 26299 28411 26305
rect 28353 26296 28365 26299
rect 26007 26268 26188 26296
rect 26007 26265 26019 26268
rect 25961 26259 26019 26265
rect 24854 26228 24860 26240
rect 24780 26200 24860 26228
rect 24854 26188 24860 26200
rect 24912 26188 24918 26240
rect 26160 26228 26188 26268
rect 27908 26268 28365 26296
rect 26234 26228 26240 26240
rect 26160 26200 26240 26228
rect 26234 26188 26240 26200
rect 26292 26188 26298 26240
rect 27246 26188 27252 26240
rect 27304 26228 27310 26240
rect 27908 26228 27936 26268
rect 28353 26265 28365 26268
rect 28399 26296 28411 26299
rect 28810 26296 28816 26308
rect 28399 26268 28816 26296
rect 28399 26265 28411 26268
rect 28353 26259 28411 26265
rect 28810 26256 28816 26268
rect 28868 26256 28874 26308
rect 29012 26305 29040 26336
rect 29365 26333 29377 26336
rect 29411 26364 29423 26367
rect 29454 26364 29460 26376
rect 29411 26336 29460 26364
rect 29411 26333 29423 26336
rect 29365 26327 29423 26333
rect 29454 26324 29460 26336
rect 29512 26324 29518 26376
rect 31294 26364 31300 26376
rect 31255 26336 31300 26364
rect 31294 26324 31300 26336
rect 31352 26324 31358 26376
rect 32306 26324 32312 26376
rect 32364 26364 32370 26376
rect 32585 26367 32643 26373
rect 32585 26364 32597 26367
rect 32364 26336 32597 26364
rect 32364 26324 32370 26336
rect 32585 26333 32597 26336
rect 32631 26333 32643 26367
rect 32766 26364 32772 26376
rect 32727 26336 32772 26364
rect 32585 26327 32643 26333
rect 32766 26324 32772 26336
rect 32824 26324 32830 26376
rect 34238 26364 34244 26376
rect 34199 26336 34244 26364
rect 34238 26324 34244 26336
rect 34296 26324 34302 26376
rect 34790 26324 34796 26376
rect 34848 26364 34854 26376
rect 35253 26367 35311 26373
rect 35253 26364 35265 26367
rect 34848 26336 35265 26364
rect 34848 26324 34854 26336
rect 35253 26333 35265 26336
rect 35299 26333 35311 26367
rect 35253 26327 35311 26333
rect 28997 26299 29055 26305
rect 28997 26265 29009 26299
rect 29043 26265 29055 26299
rect 28997 26259 29055 26265
rect 27304 26200 27936 26228
rect 27304 26188 27310 26200
rect 31202 26188 31208 26240
rect 31260 26228 31266 26240
rect 31754 26228 31760 26240
rect 31260 26200 31760 26228
rect 31260 26188 31266 26200
rect 31754 26188 31760 26200
rect 31812 26228 31818 26240
rect 32784 26228 32812 26324
rect 36633 26299 36691 26305
rect 36633 26296 36645 26299
rect 36188 26268 36645 26296
rect 33134 26228 33140 26240
rect 31812 26200 32812 26228
rect 33095 26200 33140 26228
rect 31812 26188 31818 26200
rect 33134 26188 33140 26200
rect 33192 26188 33198 26240
rect 33686 26228 33692 26240
rect 33647 26200 33692 26228
rect 33686 26188 33692 26200
rect 33744 26188 33750 26240
rect 35618 26188 35624 26240
rect 35676 26228 35682 26240
rect 36188 26228 36216 26268
rect 36633 26265 36645 26268
rect 36679 26265 36691 26299
rect 36906 26296 36912 26308
rect 36867 26268 36912 26296
rect 36633 26259 36691 26265
rect 36906 26256 36912 26268
rect 36964 26256 36970 26308
rect 35676 26200 36216 26228
rect 35676 26188 35682 26200
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 6641 26027 6699 26033
rect 6641 25993 6653 26027
rect 6687 26024 6699 26027
rect 6914 26024 6920 26036
rect 6687 25996 6920 26024
rect 6687 25993 6699 25996
rect 6641 25987 6699 25993
rect 6914 25984 6920 25996
rect 6972 25984 6978 26036
rect 8294 26024 8300 26036
rect 8255 25996 8300 26024
rect 8294 25984 8300 25996
rect 8352 25984 8358 26036
rect 11790 26024 11796 26036
rect 11751 25996 11796 26024
rect 11790 25984 11796 25996
rect 11848 25984 11854 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 17034 26024 17040 26036
rect 12492 25996 12537 26024
rect 16995 25996 17040 26024
rect 12492 25984 12498 25996
rect 17034 25984 17040 25996
rect 17092 25984 17098 26036
rect 20717 26027 20775 26033
rect 20717 25993 20729 26027
rect 20763 26024 20775 26027
rect 20806 26024 20812 26036
rect 20763 25996 20812 26024
rect 20763 25993 20775 25996
rect 20717 25987 20775 25993
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 22646 26024 22652 26036
rect 22607 25996 22652 26024
rect 22646 25984 22652 25996
rect 22704 25984 22710 26036
rect 25314 25984 25320 26036
rect 25372 26024 25378 26036
rect 26789 26027 26847 26033
rect 26789 26024 26801 26027
rect 25372 25996 26801 26024
rect 25372 25984 25378 25996
rect 26789 25993 26801 25996
rect 26835 25993 26847 26027
rect 26789 25987 26847 25993
rect 27614 25984 27620 26036
rect 27672 26024 27678 26036
rect 28169 26027 28227 26033
rect 28169 26024 28181 26027
rect 27672 25996 28181 26024
rect 27672 25984 27678 25996
rect 28169 25993 28181 25996
rect 28215 25993 28227 26027
rect 28169 25987 28227 25993
rect 28721 26027 28779 26033
rect 28721 25993 28733 26027
rect 28767 26024 28779 26027
rect 28994 26024 29000 26036
rect 28767 25996 29000 26024
rect 28767 25993 28779 25996
rect 28721 25987 28779 25993
rect 28994 25984 29000 25996
rect 29052 25984 29058 26036
rect 30374 25984 30380 26036
rect 30432 26024 30438 26036
rect 30837 26027 30895 26033
rect 30837 26024 30849 26027
rect 30432 25996 30849 26024
rect 30432 25984 30438 25996
rect 30837 25993 30849 25996
rect 30883 25993 30895 26027
rect 31202 26024 31208 26036
rect 31163 25996 31208 26024
rect 30837 25987 30895 25993
rect 18966 25916 18972 25968
rect 19024 25956 19030 25968
rect 19337 25959 19395 25965
rect 19337 25956 19349 25959
rect 19024 25928 19349 25956
rect 19024 25916 19030 25928
rect 19337 25925 19349 25928
rect 19383 25925 19395 25959
rect 25958 25956 25964 25968
rect 25919 25928 25964 25956
rect 19337 25919 19395 25925
rect 25958 25916 25964 25928
rect 26016 25916 26022 25968
rect 30852 25956 30880 25987
rect 31202 25984 31208 25996
rect 31260 25984 31266 26036
rect 31570 26024 31576 26036
rect 31531 25996 31576 26024
rect 31570 25984 31576 25996
rect 31628 25984 31634 26036
rect 32306 26024 32312 26036
rect 31772 25996 32312 26024
rect 31772 25956 31800 25996
rect 32306 25984 32312 25996
rect 32364 25984 32370 26036
rect 32674 25984 32680 26036
rect 32732 26024 32738 26036
rect 34698 26024 34704 26036
rect 32732 25996 32777 26024
rect 34659 25996 34704 26024
rect 32732 25984 32738 25996
rect 34698 25984 34704 25996
rect 34756 25984 34762 26036
rect 35526 25984 35532 26036
rect 35584 26024 35590 26036
rect 36081 26027 36139 26033
rect 36081 26024 36093 26027
rect 35584 25996 36093 26024
rect 35584 25984 35590 25996
rect 36081 25993 36093 25996
rect 36127 25993 36139 26027
rect 36081 25987 36139 25993
rect 30852 25928 31800 25956
rect 31849 25959 31907 25965
rect 31849 25925 31861 25959
rect 31895 25956 31907 25959
rect 33134 25956 33140 25968
rect 31895 25928 33140 25956
rect 31895 25925 31907 25928
rect 31849 25919 31907 25925
rect 33134 25916 33140 25928
rect 33192 25916 33198 25968
rect 10045 25891 10103 25897
rect 10045 25857 10057 25891
rect 10091 25888 10103 25891
rect 10091 25860 10272 25888
rect 10091 25857 10103 25860
rect 10045 25851 10103 25857
rect 6273 25823 6331 25829
rect 6273 25789 6285 25823
rect 6319 25820 6331 25823
rect 6917 25823 6975 25829
rect 6917 25820 6929 25823
rect 6319 25792 6929 25820
rect 6319 25789 6331 25792
rect 6273 25783 6331 25789
rect 6917 25789 6929 25792
rect 6963 25820 6975 25823
rect 7006 25820 7012 25832
rect 6963 25792 7012 25820
rect 6963 25789 6975 25792
rect 6917 25783 6975 25789
rect 7006 25780 7012 25792
rect 7064 25820 7070 25832
rect 8665 25823 8723 25829
rect 8665 25820 8677 25823
rect 7064 25792 8677 25820
rect 7064 25780 7070 25792
rect 8665 25789 8677 25792
rect 8711 25820 8723 25823
rect 9674 25820 9680 25832
rect 8711 25792 9680 25820
rect 8711 25789 8723 25792
rect 8665 25783 8723 25789
rect 9674 25780 9680 25792
rect 9732 25820 9738 25832
rect 10137 25823 10195 25829
rect 10137 25820 10149 25823
rect 9732 25792 10149 25820
rect 9732 25780 9738 25792
rect 10137 25789 10149 25792
rect 10183 25789 10195 25823
rect 10244 25820 10272 25860
rect 12894 25848 12900 25900
rect 12952 25888 12958 25900
rect 12989 25891 13047 25897
rect 12989 25888 13001 25891
rect 12952 25860 13001 25888
rect 12952 25848 12958 25860
rect 12989 25857 13001 25860
rect 13035 25857 13047 25891
rect 12989 25851 13047 25857
rect 14829 25891 14887 25897
rect 14829 25857 14841 25891
rect 14875 25888 14887 25891
rect 15197 25891 15255 25897
rect 15197 25888 15209 25891
rect 14875 25860 15209 25888
rect 14875 25857 14887 25860
rect 14829 25851 14887 25857
rect 15197 25857 15209 25860
rect 15243 25888 15255 25891
rect 20349 25891 20407 25897
rect 15243 25860 15424 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 10410 25829 10416 25832
rect 10404 25820 10416 25829
rect 10244 25792 10416 25820
rect 10137 25783 10195 25789
rect 10404 25783 10416 25792
rect 7098 25712 7104 25764
rect 7156 25761 7162 25764
rect 7156 25755 7220 25761
rect 7156 25721 7174 25755
rect 7208 25721 7220 25755
rect 10152 25752 10180 25783
rect 10410 25780 10416 25783
rect 10468 25780 10474 25832
rect 14093 25823 14151 25829
rect 14093 25789 14105 25823
rect 14139 25820 14151 25823
rect 14461 25823 14519 25829
rect 14461 25820 14473 25823
rect 14139 25792 14473 25820
rect 14139 25789 14151 25792
rect 14093 25783 14151 25789
rect 14461 25789 14473 25792
rect 14507 25820 14519 25823
rect 15286 25820 15292 25832
rect 14507 25792 15292 25820
rect 14507 25789 14519 25792
rect 14461 25783 14519 25789
rect 15286 25780 15292 25792
rect 15344 25780 15350 25832
rect 15396 25820 15424 25860
rect 20349 25857 20361 25891
rect 20395 25888 20407 25891
rect 21082 25888 21088 25900
rect 20395 25860 21088 25888
rect 20395 25857 20407 25860
rect 20349 25851 20407 25857
rect 21082 25848 21088 25860
rect 21140 25888 21146 25900
rect 21315 25891 21373 25897
rect 21315 25888 21327 25891
rect 21140 25860 21327 25888
rect 21140 25848 21146 25860
rect 21315 25857 21327 25860
rect 21361 25888 21373 25891
rect 22002 25888 22008 25900
rect 21361 25860 22008 25888
rect 21361 25857 21373 25860
rect 21315 25851 21373 25857
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25888 23535 25891
rect 24302 25888 24308 25900
rect 23523 25860 24308 25888
rect 23523 25857 23535 25860
rect 23477 25851 23535 25857
rect 24302 25848 24308 25860
rect 24360 25888 24366 25900
rect 24584 25891 24642 25897
rect 24584 25888 24596 25891
rect 24360 25860 24596 25888
rect 24360 25848 24366 25860
rect 24584 25857 24596 25860
rect 24630 25857 24642 25891
rect 24854 25888 24860 25900
rect 24815 25860 24860 25888
rect 24584 25851 24642 25857
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 26234 25848 26240 25900
rect 26292 25888 26298 25900
rect 27062 25888 27068 25900
rect 26292 25860 27068 25888
rect 26292 25848 26298 25860
rect 27062 25848 27068 25860
rect 27120 25888 27126 25900
rect 27433 25891 27491 25897
rect 27433 25888 27445 25891
rect 27120 25860 27445 25888
rect 27120 25848 27126 25860
rect 27433 25857 27445 25860
rect 27479 25888 27491 25891
rect 27522 25888 27528 25900
rect 27479 25860 27528 25888
rect 27479 25857 27491 25860
rect 27433 25851 27491 25857
rect 27522 25848 27528 25860
rect 27580 25848 27586 25900
rect 29454 25888 29460 25900
rect 29415 25860 29460 25888
rect 29454 25848 29460 25860
rect 29512 25848 29518 25900
rect 33413 25891 33471 25897
rect 33413 25857 33425 25891
rect 33459 25888 33471 25891
rect 34238 25888 34244 25900
rect 33459 25860 34244 25888
rect 33459 25857 33471 25860
rect 33413 25851 33471 25857
rect 34238 25848 34244 25860
rect 34296 25848 34302 25900
rect 15556 25823 15614 25829
rect 15556 25820 15568 25823
rect 15396 25792 15568 25820
rect 15556 25789 15568 25792
rect 15602 25820 15614 25823
rect 15930 25820 15936 25832
rect 15602 25792 15936 25820
rect 15602 25789 15614 25792
rect 15556 25783 15614 25789
rect 15930 25780 15936 25792
rect 15988 25780 15994 25832
rect 18049 25823 18107 25829
rect 18049 25789 18061 25823
rect 18095 25820 18107 25823
rect 18322 25820 18328 25832
rect 18095 25792 18328 25820
rect 18095 25789 18107 25792
rect 18049 25783 18107 25789
rect 18322 25780 18328 25792
rect 18380 25820 18386 25832
rect 18601 25823 18659 25829
rect 18601 25820 18613 25823
rect 18380 25792 18613 25820
rect 18380 25780 18386 25792
rect 18601 25789 18613 25792
rect 18647 25789 18659 25823
rect 18601 25783 18659 25789
rect 19153 25823 19211 25829
rect 19153 25789 19165 25823
rect 19199 25789 19211 25823
rect 19153 25783 19211 25789
rect 10686 25752 10692 25764
rect 10152 25724 10692 25752
rect 7156 25715 7220 25721
rect 7156 25712 7162 25715
rect 10686 25712 10692 25724
rect 10744 25712 10750 25764
rect 12897 25755 12955 25761
rect 12897 25752 12909 25755
rect 12176 25724 12909 25752
rect 11514 25684 11520 25696
rect 11475 25656 11520 25684
rect 11514 25644 11520 25656
rect 11572 25684 11578 25696
rect 12176 25693 12204 25724
rect 12897 25721 12909 25724
rect 12943 25721 12955 25755
rect 12897 25715 12955 25721
rect 12161 25687 12219 25693
rect 12161 25684 12173 25687
rect 11572 25656 12173 25684
rect 11572 25644 11578 25656
rect 12161 25653 12173 25656
rect 12207 25653 12219 25687
rect 12161 25647 12219 25653
rect 12526 25644 12532 25696
rect 12584 25684 12590 25696
rect 12805 25687 12863 25693
rect 12805 25684 12817 25687
rect 12584 25656 12817 25684
rect 12584 25644 12590 25656
rect 12805 25653 12817 25656
rect 12851 25653 12863 25687
rect 12805 25647 12863 25653
rect 15838 25644 15844 25696
rect 15896 25684 15902 25696
rect 16669 25687 16727 25693
rect 16669 25684 16681 25687
rect 15896 25656 16681 25684
rect 15896 25644 15902 25656
rect 16669 25653 16681 25656
rect 16715 25653 16727 25687
rect 16669 25647 16727 25653
rect 18233 25687 18291 25693
rect 18233 25653 18245 25687
rect 18279 25684 18291 25687
rect 18782 25684 18788 25696
rect 18279 25656 18788 25684
rect 18279 25653 18291 25656
rect 18233 25647 18291 25653
rect 18782 25644 18788 25656
rect 18840 25644 18846 25696
rect 19061 25687 19119 25693
rect 19061 25653 19073 25687
rect 19107 25684 19119 25687
rect 19168 25684 19196 25783
rect 20622 25780 20628 25832
rect 20680 25820 20686 25832
rect 20809 25823 20867 25829
rect 20809 25820 20821 25823
rect 20680 25792 20821 25820
rect 20680 25780 20686 25792
rect 20809 25789 20821 25792
rect 20855 25789 20867 25823
rect 21542 25820 21548 25832
rect 20809 25783 20867 25789
rect 20916 25792 21548 25820
rect 19702 25712 19708 25764
rect 19760 25752 19766 25764
rect 19797 25755 19855 25761
rect 19797 25752 19809 25755
rect 19760 25724 19809 25752
rect 19760 25712 19766 25724
rect 19797 25721 19809 25724
rect 19843 25752 19855 25755
rect 20916 25752 20944 25792
rect 21542 25780 21548 25792
rect 21600 25780 21606 25832
rect 23658 25780 23664 25832
rect 23716 25820 23722 25832
rect 24121 25823 24179 25829
rect 24121 25820 24133 25823
rect 23716 25792 24133 25820
rect 23716 25780 23722 25792
rect 24121 25789 24133 25792
rect 24167 25789 24179 25823
rect 27246 25820 27252 25832
rect 27207 25792 27252 25820
rect 24121 25783 24179 25789
rect 27246 25780 27252 25792
rect 27304 25780 27310 25832
rect 31570 25780 31576 25832
rect 31628 25820 31634 25832
rect 31665 25823 31723 25829
rect 31665 25820 31677 25823
rect 31628 25792 31677 25820
rect 31628 25780 31634 25792
rect 31665 25789 31677 25792
rect 31711 25789 31723 25823
rect 33134 25820 33140 25832
rect 33095 25792 33140 25820
rect 31665 25783 31723 25789
rect 33134 25780 33140 25792
rect 33192 25780 33198 25832
rect 35345 25823 35403 25829
rect 35345 25789 35357 25823
rect 35391 25820 35403 25823
rect 35618 25820 35624 25832
rect 35391 25792 35624 25820
rect 35391 25789 35403 25792
rect 35345 25783 35403 25789
rect 35618 25780 35624 25792
rect 35676 25780 35682 25832
rect 35805 25823 35863 25829
rect 35805 25789 35817 25823
rect 35851 25820 35863 25823
rect 36633 25823 36691 25829
rect 36633 25820 36645 25823
rect 35851 25792 36645 25820
rect 35851 25789 35863 25792
rect 35805 25783 35863 25789
rect 36633 25789 36645 25792
rect 36679 25820 36691 25823
rect 37185 25823 37243 25829
rect 37185 25820 37197 25823
rect 36679 25792 37197 25820
rect 36679 25789 36691 25792
rect 36633 25783 36691 25789
rect 37185 25789 37197 25792
rect 37231 25789 37243 25823
rect 37185 25783 37243 25789
rect 19843 25724 20944 25752
rect 19843 25721 19855 25724
rect 19797 25715 19855 25721
rect 26970 25712 26976 25764
rect 27028 25752 27034 25764
rect 27157 25755 27215 25761
rect 27157 25752 27169 25755
rect 27028 25724 27169 25752
rect 27028 25712 27034 25724
rect 27157 25721 27169 25724
rect 27203 25752 27215 25755
rect 27801 25755 27859 25761
rect 27801 25752 27813 25755
rect 27203 25724 27813 25752
rect 27203 25721 27215 25724
rect 27157 25715 27215 25721
rect 27801 25721 27813 25724
rect 27847 25721 27859 25755
rect 27801 25715 27859 25721
rect 29089 25755 29147 25761
rect 29089 25721 29101 25755
rect 29135 25752 29147 25755
rect 29702 25755 29760 25761
rect 29702 25752 29714 25755
rect 29135 25724 29714 25752
rect 29135 25721 29147 25724
rect 29089 25715 29147 25721
rect 29702 25721 29714 25724
rect 29748 25752 29760 25755
rect 30742 25752 30748 25764
rect 29748 25724 30748 25752
rect 29748 25721 29760 25724
rect 29702 25715 29760 25721
rect 30742 25712 30748 25724
rect 30800 25712 30806 25764
rect 35437 25755 35495 25761
rect 35437 25721 35449 25755
rect 35483 25752 35495 25755
rect 35526 25752 35532 25764
rect 35483 25724 35532 25752
rect 35483 25721 35495 25724
rect 35437 25715 35495 25721
rect 35526 25712 35532 25724
rect 35584 25712 35590 25764
rect 19242 25684 19248 25696
rect 19107 25656 19248 25684
rect 19107 25653 19119 25656
rect 19061 25647 19119 25653
rect 19242 25644 19248 25656
rect 19300 25644 19306 25696
rect 20806 25644 20812 25696
rect 20864 25684 20870 25696
rect 21275 25687 21333 25693
rect 21275 25684 21287 25687
rect 20864 25656 21287 25684
rect 20864 25644 20870 25656
rect 21275 25653 21287 25656
rect 21321 25684 21333 25687
rect 24029 25687 24087 25693
rect 24029 25684 24041 25687
rect 21321 25656 24041 25684
rect 21321 25653 21333 25656
rect 21275 25647 21333 25653
rect 24029 25653 24041 25656
rect 24075 25684 24087 25687
rect 24587 25687 24645 25693
rect 24587 25684 24599 25687
rect 24075 25656 24599 25684
rect 24075 25653 24087 25656
rect 24029 25647 24087 25653
rect 24587 25653 24599 25656
rect 24633 25684 24645 25687
rect 26602 25684 26608 25696
rect 24633 25656 26608 25684
rect 24633 25653 24645 25656
rect 24587 25647 24645 25653
rect 26602 25644 26608 25656
rect 26660 25644 26666 25696
rect 32766 25684 32772 25696
rect 32727 25656 32772 25684
rect 32766 25644 32772 25656
rect 32824 25644 32830 25696
rect 32858 25644 32864 25696
rect 32916 25684 32922 25696
rect 33229 25687 33287 25693
rect 33229 25684 33241 25687
rect 32916 25656 33241 25684
rect 32916 25644 32922 25656
rect 33229 25653 33241 25656
rect 33275 25653 33287 25687
rect 33778 25684 33784 25696
rect 33739 25656 33784 25684
rect 33229 25647 33287 25653
rect 33778 25644 33784 25656
rect 33836 25644 33842 25696
rect 33870 25644 33876 25696
rect 33928 25684 33934 25696
rect 34149 25687 34207 25693
rect 34149 25684 34161 25687
rect 33928 25656 34161 25684
rect 33928 25644 33934 25656
rect 34149 25653 34161 25656
rect 34195 25653 34207 25687
rect 34149 25647 34207 25653
rect 34790 25644 34796 25696
rect 34848 25684 34854 25696
rect 36449 25687 36507 25693
rect 36449 25684 36461 25687
rect 34848 25656 36461 25684
rect 34848 25644 34854 25656
rect 36449 25653 36461 25656
rect 36495 25653 36507 25687
rect 36814 25684 36820 25696
rect 36775 25656 36820 25684
rect 36449 25647 36507 25653
rect 36814 25644 36820 25656
rect 36872 25644 36878 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 10597 25483 10655 25489
rect 10597 25449 10609 25483
rect 10643 25480 10655 25483
rect 10686 25480 10692 25492
rect 10643 25452 10692 25480
rect 10643 25449 10655 25452
rect 10597 25443 10655 25449
rect 10686 25440 10692 25452
rect 10744 25480 10750 25492
rect 10962 25480 10968 25492
rect 10744 25452 10968 25480
rect 10744 25440 10750 25452
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 12526 25480 12532 25492
rect 12487 25452 12532 25480
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 19150 25440 19156 25492
rect 19208 25480 19214 25492
rect 19245 25483 19303 25489
rect 19245 25480 19257 25483
rect 19208 25452 19257 25480
rect 19208 25440 19214 25452
rect 19245 25449 19257 25452
rect 19291 25449 19303 25483
rect 20714 25480 20720 25492
rect 20675 25452 20720 25480
rect 19245 25443 19303 25449
rect 20714 25440 20720 25452
rect 20772 25440 20778 25492
rect 21082 25480 21088 25492
rect 21043 25452 21088 25480
rect 21082 25440 21088 25452
rect 21140 25440 21146 25492
rect 21542 25480 21548 25492
rect 21503 25452 21548 25480
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 23658 25480 23664 25492
rect 23619 25452 23664 25480
rect 23658 25440 23664 25452
rect 23716 25440 23722 25492
rect 25314 25440 25320 25492
rect 25372 25480 25378 25492
rect 25869 25483 25927 25489
rect 25869 25480 25881 25483
rect 25372 25452 25881 25480
rect 25372 25440 25378 25452
rect 25869 25449 25881 25452
rect 25915 25449 25927 25483
rect 26234 25480 26240 25492
rect 26195 25452 26240 25480
rect 25869 25443 25927 25449
rect 26234 25440 26240 25452
rect 26292 25440 26298 25492
rect 26881 25483 26939 25489
rect 26881 25449 26893 25483
rect 26927 25480 26939 25483
rect 27246 25480 27252 25492
rect 26927 25452 27252 25480
rect 26927 25449 26939 25452
rect 26881 25443 26939 25449
rect 27246 25440 27252 25452
rect 27304 25440 27310 25492
rect 27522 25480 27528 25492
rect 27483 25452 27528 25480
rect 27522 25440 27528 25452
rect 27580 25440 27586 25492
rect 29273 25483 29331 25489
rect 29273 25449 29285 25483
rect 29319 25480 29331 25483
rect 29454 25480 29460 25492
rect 29319 25452 29460 25480
rect 29319 25449 29331 25452
rect 29273 25443 29331 25449
rect 29454 25440 29460 25452
rect 29512 25440 29518 25492
rect 30742 25480 30748 25492
rect 30703 25452 30748 25480
rect 30742 25440 30748 25452
rect 30800 25440 30806 25492
rect 32493 25483 32551 25489
rect 32493 25449 32505 25483
rect 32539 25480 32551 25483
rect 33778 25480 33784 25492
rect 32539 25452 33784 25480
rect 32539 25449 32551 25452
rect 32493 25443 32551 25449
rect 33778 25440 33784 25452
rect 33836 25440 33842 25492
rect 34238 25440 34244 25492
rect 34296 25480 34302 25492
rect 34425 25483 34483 25489
rect 34425 25480 34437 25483
rect 34296 25452 34437 25480
rect 34296 25440 34302 25452
rect 34425 25449 34437 25452
rect 34471 25449 34483 25483
rect 34425 25443 34483 25449
rect 14001 25415 14059 25421
rect 14001 25381 14013 25415
rect 14047 25412 14059 25415
rect 14090 25412 14096 25424
rect 14047 25384 14096 25412
rect 14047 25381 14059 25384
rect 14001 25375 14059 25381
rect 14090 25372 14096 25384
rect 14148 25372 14154 25424
rect 20349 25415 20407 25421
rect 20349 25381 20361 25415
rect 20395 25412 20407 25415
rect 20622 25412 20628 25424
rect 20395 25384 20628 25412
rect 20395 25381 20407 25384
rect 20349 25375 20407 25381
rect 20622 25372 20628 25384
rect 20680 25372 20686 25424
rect 20990 25372 20996 25424
rect 21048 25412 21054 25424
rect 21821 25415 21879 25421
rect 21821 25412 21833 25415
rect 21048 25384 21833 25412
rect 21048 25372 21054 25384
rect 21821 25381 21833 25384
rect 21867 25381 21879 25415
rect 21821 25375 21879 25381
rect 24121 25415 24179 25421
rect 24121 25381 24133 25415
rect 24167 25412 24179 25415
rect 24210 25412 24216 25424
rect 24167 25384 24216 25412
rect 24167 25381 24179 25384
rect 24121 25375 24179 25381
rect 24210 25372 24216 25384
rect 24268 25412 24274 25424
rect 24480 25415 24538 25421
rect 24480 25412 24492 25415
rect 24268 25384 24492 25412
rect 24268 25372 24274 25384
rect 24480 25381 24492 25384
rect 24526 25412 24538 25415
rect 24670 25412 24676 25424
rect 24526 25384 24676 25412
rect 24526 25381 24538 25384
rect 24480 25375 24538 25381
rect 24670 25372 24676 25384
rect 24728 25372 24734 25424
rect 26970 25372 26976 25424
rect 27028 25412 27034 25424
rect 27157 25415 27215 25421
rect 27157 25412 27169 25415
rect 27028 25384 27169 25412
rect 27028 25372 27034 25384
rect 27157 25381 27169 25384
rect 27203 25381 27215 25415
rect 27157 25375 27215 25381
rect 33321 25415 33379 25421
rect 33321 25381 33333 25415
rect 33367 25412 33379 25415
rect 34256 25412 34284 25440
rect 33367 25384 34284 25412
rect 33367 25381 33379 25384
rect 33321 25375 33379 25381
rect 34698 25372 34704 25424
rect 34756 25412 34762 25424
rect 35244 25415 35302 25421
rect 35244 25412 35256 25415
rect 34756 25384 35256 25412
rect 34756 25372 34762 25384
rect 35244 25381 35256 25384
rect 35290 25412 35302 25415
rect 35618 25412 35624 25424
rect 35290 25384 35624 25412
rect 35290 25381 35302 25384
rect 35244 25375 35302 25381
rect 35618 25372 35624 25384
rect 35676 25372 35682 25424
rect 7006 25304 7012 25356
rect 7064 25344 7070 25356
rect 7101 25347 7159 25353
rect 7101 25344 7113 25347
rect 7064 25316 7113 25344
rect 7064 25304 7070 25316
rect 7101 25313 7113 25316
rect 7147 25313 7159 25347
rect 7101 25307 7159 25313
rect 7190 25304 7196 25356
rect 7248 25344 7254 25356
rect 7357 25347 7415 25353
rect 7357 25344 7369 25347
rect 7248 25316 7369 25344
rect 7248 25304 7254 25316
rect 7357 25313 7369 25316
rect 7403 25313 7415 25347
rect 7357 25307 7415 25313
rect 10042 25304 10048 25356
rect 10100 25344 10106 25356
rect 10945 25347 11003 25353
rect 10945 25344 10957 25347
rect 10100 25316 10957 25344
rect 10100 25304 10106 25316
rect 10945 25313 10957 25316
rect 10991 25344 11003 25347
rect 11514 25344 11520 25356
rect 10991 25316 11520 25344
rect 10991 25313 11003 25316
rect 10945 25307 11003 25313
rect 11514 25304 11520 25316
rect 11572 25304 11578 25356
rect 15102 25344 15108 25356
rect 14108 25316 15108 25344
rect 10686 25276 10692 25288
rect 10647 25248 10692 25276
rect 10686 25236 10692 25248
rect 10744 25236 10750 25288
rect 13722 25236 13728 25288
rect 13780 25276 13786 25288
rect 14108 25285 14136 25316
rect 15102 25304 15108 25316
rect 15160 25304 15166 25356
rect 15545 25347 15603 25353
rect 15545 25344 15557 25347
rect 15212 25316 15557 25344
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 13780 25248 14105 25276
rect 13780 25236 13786 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 14277 25279 14335 25285
rect 14277 25245 14289 25279
rect 14323 25276 14335 25279
rect 14458 25276 14464 25288
rect 14323 25248 14464 25276
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 7009 25143 7067 25149
rect 7009 25109 7021 25143
rect 7055 25140 7067 25143
rect 7098 25140 7104 25152
rect 7055 25112 7104 25140
rect 7055 25109 7067 25112
rect 7009 25103 7067 25109
rect 7098 25100 7104 25112
rect 7156 25140 7162 25152
rect 8202 25140 8208 25152
rect 7156 25112 8208 25140
rect 7156 25100 7162 25112
rect 8202 25100 8208 25112
rect 8260 25140 8266 25152
rect 8481 25143 8539 25149
rect 8481 25140 8493 25143
rect 8260 25112 8493 25140
rect 8260 25100 8266 25112
rect 8481 25109 8493 25112
rect 8527 25109 8539 25143
rect 10134 25140 10140 25152
rect 10095 25112 10140 25140
rect 8481 25103 8539 25109
rect 10134 25100 10140 25112
rect 10192 25100 10198 25152
rect 11054 25100 11060 25152
rect 11112 25140 11118 25152
rect 12069 25143 12127 25149
rect 12069 25140 12081 25143
rect 11112 25112 12081 25140
rect 11112 25100 11118 25112
rect 12069 25109 12081 25112
rect 12115 25140 12127 25143
rect 12526 25140 12532 25152
rect 12115 25112 12532 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 12526 25100 12532 25112
rect 12584 25100 12590 25152
rect 12894 25140 12900 25152
rect 12855 25112 12900 25140
rect 12894 25100 12900 25112
rect 12952 25100 12958 25152
rect 13630 25140 13636 25152
rect 13591 25112 13636 25140
rect 13630 25100 13636 25112
rect 13688 25100 13694 25152
rect 14734 25140 14740 25152
rect 14695 25112 14740 25140
rect 14734 25100 14740 25112
rect 14792 25100 14798 25152
rect 15010 25140 15016 25152
rect 14971 25112 15016 25140
rect 15010 25100 15016 25112
rect 15068 25140 15074 25152
rect 15212 25140 15240 25316
rect 15545 25313 15557 25316
rect 15591 25344 15603 25347
rect 15838 25344 15844 25356
rect 15591 25316 15844 25344
rect 15591 25313 15603 25316
rect 15545 25307 15603 25313
rect 15838 25304 15844 25316
rect 15896 25304 15902 25356
rect 18138 25344 18144 25356
rect 18099 25316 18144 25344
rect 18138 25304 18144 25316
rect 18196 25304 18202 25356
rect 19610 25344 19616 25356
rect 19571 25316 19616 25344
rect 19610 25304 19616 25316
rect 19668 25304 19674 25356
rect 19705 25347 19763 25353
rect 19705 25313 19717 25347
rect 19751 25344 19763 25347
rect 20254 25344 20260 25356
rect 19751 25316 20260 25344
rect 19751 25313 19763 25316
rect 19705 25307 19763 25313
rect 20254 25304 20260 25316
rect 20312 25304 20318 25356
rect 20898 25344 20904 25356
rect 20859 25316 20904 25344
rect 20898 25304 20904 25316
rect 20956 25304 20962 25356
rect 28166 25344 28172 25356
rect 28127 25316 28172 25344
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 28261 25347 28319 25353
rect 28261 25313 28273 25347
rect 28307 25344 28319 25347
rect 28810 25344 28816 25356
rect 28307 25316 28816 25344
rect 28307 25313 28319 25316
rect 28261 25307 28319 25313
rect 28810 25304 28816 25316
rect 28868 25304 28874 25356
rect 28994 25304 29000 25356
rect 29052 25344 29058 25356
rect 29621 25347 29679 25353
rect 29621 25344 29633 25347
rect 29052 25316 29633 25344
rect 29052 25304 29058 25316
rect 29621 25313 29633 25316
rect 29667 25313 29679 25347
rect 29621 25307 29679 25313
rect 31757 25347 31815 25353
rect 31757 25313 31769 25347
rect 31803 25344 31815 25347
rect 31938 25344 31944 25356
rect 31803 25316 31944 25344
rect 31803 25313 31815 25316
rect 31757 25307 31815 25313
rect 31938 25304 31944 25316
rect 31996 25304 32002 25356
rect 32122 25304 32128 25356
rect 32180 25344 32186 25356
rect 32309 25347 32367 25353
rect 32309 25344 32321 25347
rect 32180 25316 32321 25344
rect 32180 25304 32186 25316
rect 32309 25313 32321 25316
rect 32355 25313 32367 25347
rect 32309 25307 32367 25313
rect 33686 25304 33692 25356
rect 33744 25344 33750 25356
rect 33781 25347 33839 25353
rect 33781 25344 33793 25347
rect 33744 25316 33793 25344
rect 33744 25304 33750 25316
rect 33781 25313 33793 25316
rect 33827 25313 33839 25347
rect 33781 25307 33839 25313
rect 15286 25236 15292 25288
rect 15344 25276 15350 25288
rect 15344 25248 15437 25276
rect 15344 25236 15350 25248
rect 16666 25236 16672 25288
rect 16724 25276 16730 25288
rect 16945 25279 17003 25285
rect 16945 25276 16957 25279
rect 16724 25248 16957 25276
rect 16724 25236 16730 25248
rect 16945 25245 16957 25248
rect 16991 25245 17003 25279
rect 16945 25239 17003 25245
rect 19153 25279 19211 25285
rect 19153 25245 19165 25279
rect 19199 25276 19211 25279
rect 19794 25276 19800 25288
rect 19199 25248 19800 25276
rect 19199 25245 19211 25248
rect 19153 25239 19211 25245
rect 19794 25236 19800 25248
rect 19852 25236 19858 25288
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25276 23259 25279
rect 23474 25276 23480 25288
rect 23247 25248 23480 25276
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 23474 25236 23480 25248
rect 23532 25236 23538 25288
rect 23842 25236 23848 25288
rect 23900 25276 23906 25288
rect 24213 25279 24271 25285
rect 24213 25276 24225 25279
rect 23900 25248 24225 25276
rect 23900 25236 23906 25248
rect 24213 25245 24225 25248
rect 24259 25245 24271 25279
rect 28442 25276 28448 25288
rect 28403 25248 28448 25276
rect 24213 25239 24271 25245
rect 28442 25236 28448 25248
rect 28500 25236 28506 25288
rect 29362 25276 29368 25288
rect 29323 25248 29368 25276
rect 29362 25236 29368 25248
rect 29420 25236 29426 25288
rect 32766 25236 32772 25288
rect 32824 25276 32830 25288
rect 33873 25279 33931 25285
rect 33873 25276 33885 25279
rect 32824 25248 33885 25276
rect 32824 25236 32830 25248
rect 33873 25245 33885 25248
rect 33919 25245 33931 25279
rect 34054 25276 34060 25288
rect 34015 25248 34060 25276
rect 33873 25239 33931 25245
rect 34054 25236 34060 25248
rect 34112 25236 34118 25288
rect 34977 25279 35035 25285
rect 34977 25276 34989 25279
rect 34808 25248 34989 25276
rect 15068 25112 15240 25140
rect 15311 25140 15339 25236
rect 31573 25211 31631 25217
rect 31573 25177 31585 25211
rect 31619 25208 31631 25211
rect 34808 25208 34836 25248
rect 34977 25245 34989 25248
rect 35023 25245 35035 25279
rect 34977 25239 35035 25245
rect 31619 25180 34836 25208
rect 31619 25177 31631 25180
rect 31573 25171 31631 25177
rect 34808 25152 34836 25180
rect 15930 25140 15936 25152
rect 15311 25112 15936 25140
rect 15068 25100 15074 25112
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 16669 25143 16727 25149
rect 16669 25140 16681 25143
rect 16632 25112 16681 25140
rect 16632 25100 16638 25112
rect 16669 25109 16681 25112
rect 16715 25109 16727 25143
rect 17402 25140 17408 25152
rect 17363 25112 17408 25140
rect 16669 25103 16727 25109
rect 17402 25100 17408 25112
rect 17460 25100 17466 25152
rect 18325 25143 18383 25149
rect 18325 25109 18337 25143
rect 18371 25140 18383 25143
rect 18598 25140 18604 25152
rect 18371 25112 18604 25140
rect 18371 25109 18383 25112
rect 18325 25103 18383 25109
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 18690 25100 18696 25152
rect 18748 25140 18754 25152
rect 18748 25112 18793 25140
rect 18748 25100 18754 25112
rect 24854 25100 24860 25152
rect 24912 25140 24918 25152
rect 25593 25143 25651 25149
rect 25593 25140 25605 25143
rect 24912 25112 25605 25140
rect 24912 25100 24918 25112
rect 25593 25109 25605 25112
rect 25639 25109 25651 25143
rect 27798 25140 27804 25152
rect 27759 25112 27804 25140
rect 25593 25103 25651 25109
rect 27798 25100 27804 25112
rect 27856 25100 27862 25152
rect 32858 25140 32864 25152
rect 32819 25112 32864 25140
rect 32858 25100 32864 25112
rect 32916 25100 32922 25152
rect 33410 25140 33416 25152
rect 33371 25112 33416 25140
rect 33410 25100 33416 25112
rect 33468 25100 33474 25152
rect 34790 25140 34796 25152
rect 34751 25112 34796 25140
rect 34790 25100 34796 25112
rect 34848 25100 34854 25152
rect 36354 25140 36360 25152
rect 36315 25112 36360 25140
rect 36354 25100 36360 25112
rect 36412 25100 36418 25152
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 6641 24939 6699 24945
rect 6641 24905 6653 24939
rect 6687 24936 6699 24939
rect 7006 24936 7012 24948
rect 6687 24908 7012 24936
rect 6687 24905 6699 24908
rect 6641 24899 6699 24905
rect 7006 24896 7012 24908
rect 7064 24896 7070 24948
rect 9674 24936 9680 24948
rect 9635 24908 9680 24936
rect 9674 24896 9680 24908
rect 9732 24896 9738 24948
rect 10042 24936 10048 24948
rect 10003 24908 10048 24936
rect 10042 24896 10048 24908
rect 10100 24896 10106 24948
rect 12434 24896 12440 24948
rect 12492 24936 12498 24948
rect 14737 24939 14795 24945
rect 12492 24908 12537 24936
rect 12492 24896 12498 24908
rect 14737 24905 14749 24939
rect 14783 24936 14795 24939
rect 15010 24936 15016 24948
rect 14783 24908 15016 24936
rect 14783 24905 14795 24908
rect 14737 24899 14795 24905
rect 15010 24896 15016 24908
rect 15068 24896 15074 24948
rect 18322 24936 18328 24948
rect 18283 24908 18328 24936
rect 18322 24896 18328 24908
rect 18380 24896 18386 24948
rect 19794 24936 19800 24948
rect 19755 24908 19800 24936
rect 19794 24896 19800 24908
rect 19852 24896 19858 24948
rect 20806 24896 20812 24948
rect 20864 24936 20870 24948
rect 21269 24939 21327 24945
rect 21269 24936 21281 24939
rect 20864 24908 21281 24936
rect 20864 24896 20870 24908
rect 21269 24905 21281 24908
rect 21315 24905 21327 24939
rect 21269 24899 21327 24905
rect 23477 24939 23535 24945
rect 23477 24905 23489 24939
rect 23523 24936 23535 24939
rect 23842 24936 23848 24948
rect 23523 24908 23848 24936
rect 23523 24905 23535 24908
rect 23477 24899 23535 24905
rect 23842 24896 23848 24908
rect 23900 24896 23906 24948
rect 24210 24936 24216 24948
rect 24171 24908 24216 24936
rect 24210 24896 24216 24908
rect 24268 24896 24274 24948
rect 27525 24939 27583 24945
rect 27525 24905 27537 24939
rect 27571 24936 27583 24939
rect 28442 24936 28448 24948
rect 27571 24908 28448 24936
rect 27571 24905 27583 24908
rect 27525 24899 27583 24905
rect 28442 24896 28448 24908
rect 28500 24896 28506 24948
rect 28994 24896 29000 24948
rect 29052 24936 29058 24948
rect 30653 24939 30711 24945
rect 30653 24936 30665 24939
rect 29052 24908 30665 24936
rect 29052 24896 29058 24908
rect 30653 24905 30665 24908
rect 30699 24905 30711 24939
rect 30653 24899 30711 24905
rect 12894 24828 12900 24880
rect 12952 24868 12958 24880
rect 12952 24840 13032 24868
rect 12952 24828 12958 24840
rect 11882 24800 11888 24812
rect 11843 24772 11888 24800
rect 11882 24760 11888 24772
rect 11940 24760 11946 24812
rect 13004 24809 13032 24840
rect 15930 24828 15936 24880
rect 15988 24868 15994 24880
rect 17037 24871 17095 24877
rect 17037 24868 17049 24871
rect 15988 24840 17049 24868
rect 15988 24828 15994 24840
rect 17037 24837 17049 24840
rect 17083 24868 17095 24871
rect 17083 24840 18644 24868
rect 17083 24837 17095 24840
rect 17037 24831 17095 24837
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 13722 24800 13728 24812
rect 13683 24772 13728 24800
rect 12989 24763 13047 24769
rect 13722 24760 13728 24772
rect 13780 24760 13786 24812
rect 7374 24732 7380 24744
rect 7335 24704 7380 24732
rect 7374 24692 7380 24704
rect 7432 24692 7438 24744
rect 10134 24732 10140 24744
rect 10095 24704 10140 24732
rect 10134 24692 10140 24704
rect 10192 24692 10198 24744
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 14829 24735 14887 24741
rect 14829 24732 14841 24735
rect 14792 24704 14841 24732
rect 14792 24692 14798 24704
rect 14829 24701 14841 24704
rect 14875 24732 14887 24735
rect 15948 24732 15976 24828
rect 16577 24803 16635 24809
rect 16577 24769 16589 24803
rect 16623 24800 16635 24803
rect 16945 24803 17003 24809
rect 16945 24800 16957 24803
rect 16623 24772 16957 24800
rect 16623 24769 16635 24772
rect 16577 24763 16635 24769
rect 16945 24769 16957 24772
rect 16991 24800 17003 24803
rect 17494 24800 17500 24812
rect 16991 24772 17500 24800
rect 16991 24769 17003 24772
rect 16945 24763 17003 24769
rect 17494 24760 17500 24772
rect 17552 24800 17558 24812
rect 17862 24800 17868 24812
rect 17552 24772 17868 24800
rect 17552 24760 17558 24772
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 18616 24744 18644 24840
rect 18966 24800 18972 24812
rect 18927 24772 18972 24800
rect 18966 24760 18972 24772
rect 19024 24760 19030 24812
rect 19812 24800 19840 24896
rect 20898 24828 20904 24880
rect 20956 24868 20962 24880
rect 21545 24871 21603 24877
rect 21545 24868 21557 24871
rect 20956 24840 21557 24868
rect 20956 24828 20962 24840
rect 21545 24837 21557 24840
rect 21591 24837 21603 24871
rect 21545 24831 21603 24837
rect 19812 24772 20024 24800
rect 19996 24744 20024 24772
rect 20990 24760 20996 24812
rect 21048 24800 21054 24812
rect 21913 24803 21971 24809
rect 21913 24800 21925 24803
rect 21048 24772 21925 24800
rect 21048 24760 21054 24772
rect 21913 24769 21925 24772
rect 21959 24769 21971 24803
rect 23934 24800 23940 24812
rect 23895 24772 23940 24800
rect 21913 24763 21971 24769
rect 23934 24760 23940 24772
rect 23992 24800 23998 24812
rect 28721 24803 28779 24809
rect 23992 24772 24624 24800
rect 23992 24760 23998 24772
rect 14875 24704 15976 24732
rect 17221 24735 17279 24741
rect 14875 24701 14887 24704
rect 14829 24695 14887 24701
rect 17221 24701 17233 24735
rect 17267 24732 17279 24735
rect 17402 24732 17408 24744
rect 17267 24704 17408 24732
rect 17267 24701 17279 24704
rect 17221 24695 17279 24701
rect 17402 24692 17408 24704
rect 17460 24692 17466 24744
rect 18598 24692 18604 24744
rect 18656 24732 18662 24744
rect 19886 24732 19892 24744
rect 18656 24704 19892 24732
rect 18656 24692 18662 24704
rect 19886 24692 19892 24704
rect 19944 24692 19950 24744
rect 19978 24692 19984 24744
rect 20036 24732 20042 24744
rect 20145 24735 20203 24741
rect 20145 24732 20157 24735
rect 20036 24704 20157 24732
rect 20036 24692 20042 24704
rect 20145 24701 20157 24704
rect 20191 24701 20203 24735
rect 20145 24695 20203 24701
rect 24489 24735 24547 24741
rect 24489 24701 24501 24735
rect 24535 24701 24547 24735
rect 24596 24732 24624 24772
rect 28721 24769 28733 24803
rect 28767 24800 28779 24803
rect 28994 24800 29000 24812
rect 28767 24772 29000 24800
rect 28767 24769 28779 24772
rect 28721 24763 28779 24769
rect 28994 24760 29000 24772
rect 29052 24760 29058 24812
rect 30668 24800 30696 24899
rect 32122 24896 32128 24948
rect 32180 24936 32186 24948
rect 32493 24939 32551 24945
rect 32493 24936 32505 24939
rect 32180 24908 32505 24936
rect 32180 24896 32186 24908
rect 32493 24905 32505 24908
rect 32539 24905 32551 24939
rect 32493 24899 32551 24905
rect 32766 24896 32772 24948
rect 32824 24936 32830 24948
rect 33134 24936 33140 24948
rect 32824 24908 33140 24936
rect 32824 24896 32830 24908
rect 33134 24896 33140 24908
rect 33192 24896 33198 24948
rect 33870 24936 33876 24948
rect 33831 24908 33876 24936
rect 33870 24896 33876 24908
rect 33928 24896 33934 24948
rect 34698 24936 34704 24948
rect 34659 24908 34704 24936
rect 34698 24896 34704 24908
rect 34756 24896 34762 24948
rect 36354 24936 36360 24948
rect 36315 24908 36360 24936
rect 36354 24896 36360 24908
rect 36412 24896 36418 24948
rect 36630 24936 36636 24948
rect 36591 24908 36636 24936
rect 36630 24896 36636 24908
rect 36688 24896 36694 24948
rect 31021 24871 31079 24877
rect 31021 24837 31033 24871
rect 31067 24868 31079 24871
rect 31294 24868 31300 24880
rect 31067 24840 31300 24868
rect 31067 24837 31079 24840
rect 31021 24831 31079 24837
rect 31294 24828 31300 24840
rect 31352 24868 31358 24880
rect 31754 24868 31760 24880
rect 31352 24840 31760 24868
rect 31352 24828 31358 24840
rect 31754 24828 31760 24840
rect 31812 24868 31818 24880
rect 31812 24840 32076 24868
rect 31812 24828 31818 24840
rect 32048 24809 32076 24840
rect 31389 24803 31447 24809
rect 31389 24800 31401 24803
rect 30668 24772 31401 24800
rect 31389 24769 31401 24772
rect 31435 24800 31447 24803
rect 31941 24803 31999 24809
rect 31941 24800 31953 24803
rect 31435 24772 31953 24800
rect 31435 24769 31447 24772
rect 31389 24763 31447 24769
rect 31941 24769 31953 24772
rect 31987 24769 31999 24803
rect 31941 24763 31999 24769
rect 32033 24803 32091 24809
rect 32033 24769 32045 24803
rect 32079 24769 32091 24803
rect 32033 24763 32091 24769
rect 32766 24760 32772 24812
rect 32824 24800 32830 24812
rect 34241 24803 34299 24809
rect 34241 24800 34253 24803
rect 32824 24772 34253 24800
rect 32824 24760 32830 24772
rect 34241 24769 34253 24772
rect 34287 24800 34299 24803
rect 35529 24803 35587 24809
rect 34287 24772 35296 24800
rect 34287 24769 34299 24772
rect 34241 24763 34299 24769
rect 24762 24741 24768 24744
rect 24745 24735 24768 24741
rect 24745 24732 24757 24735
rect 24596 24704 24757 24732
rect 24489 24695 24547 24701
rect 24745 24701 24757 24704
rect 24820 24732 24826 24744
rect 29273 24735 29331 24741
rect 24820 24704 24893 24732
rect 24745 24695 24768 24701
rect 7650 24673 7656 24676
rect 7285 24667 7343 24673
rect 7285 24633 7297 24667
rect 7331 24664 7343 24667
rect 7644 24664 7656 24673
rect 7331 24636 7656 24664
rect 7331 24633 7343 24636
rect 7285 24627 7343 24633
rect 7644 24627 7656 24636
rect 7650 24624 7656 24627
rect 7708 24624 7714 24676
rect 10226 24624 10232 24676
rect 10284 24664 10290 24676
rect 15102 24673 15108 24676
rect 10382 24667 10440 24673
rect 10382 24664 10394 24667
rect 10284 24636 10394 24664
rect 10284 24624 10290 24636
rect 10382 24633 10394 24636
rect 10428 24633 10440 24667
rect 12897 24667 12955 24673
rect 12897 24664 12909 24667
rect 10382 24627 10440 24633
rect 12176 24636 12909 24664
rect 12176 24608 12204 24636
rect 12897 24633 12909 24636
rect 12943 24633 12955 24667
rect 15096 24664 15108 24673
rect 15063 24636 15108 24664
rect 12897 24627 12955 24633
rect 15096 24627 15108 24636
rect 15102 24624 15108 24627
rect 15160 24624 15166 24676
rect 18138 24664 18144 24676
rect 17788 24636 18144 24664
rect 17788 24608 17816 24636
rect 18138 24624 18144 24636
rect 18196 24664 18202 24676
rect 18785 24667 18843 24673
rect 18785 24664 18797 24667
rect 18196 24636 18797 24664
rect 18196 24624 18202 24636
rect 18785 24633 18797 24636
rect 18831 24633 18843 24667
rect 18785 24627 18843 24633
rect 19429 24667 19487 24673
rect 19429 24633 19441 24667
rect 19475 24664 19487 24667
rect 19610 24664 19616 24676
rect 19475 24636 19616 24664
rect 19475 24633 19487 24636
rect 19429 24627 19487 24633
rect 19610 24624 19616 24636
rect 19668 24664 19674 24676
rect 22097 24667 22155 24673
rect 22097 24664 22109 24667
rect 19668 24636 22109 24664
rect 19668 24624 19674 24636
rect 22097 24633 22109 24636
rect 22143 24633 22155 24667
rect 24504 24664 24532 24695
rect 24762 24692 24768 24695
rect 24820 24692 24826 24704
rect 29273 24701 29285 24735
rect 29319 24732 29331 24735
rect 29362 24732 29368 24744
rect 29319 24704 29368 24732
rect 29319 24701 29331 24704
rect 29273 24695 29331 24701
rect 29362 24692 29368 24704
rect 29420 24692 29426 24744
rect 33597 24735 33655 24741
rect 33597 24701 33609 24735
rect 33643 24732 33655 24735
rect 33689 24735 33747 24741
rect 33689 24732 33701 24735
rect 33643 24704 33701 24732
rect 33643 24701 33655 24704
rect 33597 24695 33655 24701
rect 33689 24701 33701 24704
rect 33735 24732 33747 24735
rect 34422 24732 34428 24744
rect 33735 24704 34428 24732
rect 33735 24701 33747 24704
rect 33689 24695 33747 24701
rect 34422 24692 34428 24704
rect 34480 24692 34486 24744
rect 35268 24741 35296 24772
rect 35529 24769 35541 24803
rect 35575 24800 35587 24803
rect 35894 24800 35900 24812
rect 35575 24772 35900 24800
rect 35575 24769 35587 24772
rect 35529 24763 35587 24769
rect 35894 24760 35900 24772
rect 35952 24800 35958 24812
rect 36372 24800 36400 24896
rect 37093 24803 37151 24809
rect 37093 24800 37105 24803
rect 35952 24772 36400 24800
rect 36464 24772 37105 24800
rect 35952 24760 35958 24772
rect 36464 24741 36492 24772
rect 37093 24769 37105 24772
rect 37139 24800 37151 24803
rect 37182 24800 37188 24812
rect 37139 24772 37188 24800
rect 37139 24769 37151 24772
rect 37093 24763 37151 24769
rect 37182 24760 37188 24772
rect 37240 24760 37246 24812
rect 35253 24735 35311 24741
rect 35253 24701 35265 24735
rect 35299 24701 35311 24735
rect 35253 24695 35311 24701
rect 36449 24735 36507 24741
rect 36449 24701 36461 24735
rect 36495 24701 36507 24735
rect 36449 24695 36507 24701
rect 24578 24664 24584 24676
rect 24491 24636 24584 24664
rect 22097 24627 22155 24633
rect 24578 24624 24584 24636
rect 24636 24664 24642 24676
rect 26237 24667 26295 24673
rect 26237 24664 26249 24667
rect 24636 24636 26249 24664
rect 24636 24624 24642 24636
rect 26237 24633 26249 24636
rect 26283 24633 26295 24667
rect 26237 24627 26295 24633
rect 27893 24667 27951 24673
rect 27893 24633 27905 24667
rect 27939 24664 27951 24667
rect 28810 24664 28816 24676
rect 27939 24636 28816 24664
rect 27939 24633 27951 24636
rect 27893 24627 27951 24633
rect 28810 24624 28816 24636
rect 28868 24624 28874 24676
rect 29089 24667 29147 24673
rect 29089 24633 29101 24667
rect 29135 24664 29147 24667
rect 29518 24667 29576 24673
rect 29518 24664 29530 24667
rect 29135 24636 29530 24664
rect 29135 24633 29147 24636
rect 29089 24627 29147 24633
rect 29518 24633 29530 24636
rect 29564 24664 29576 24667
rect 30558 24664 30564 24676
rect 29564 24636 30564 24664
rect 29564 24633 29576 24636
rect 29518 24627 29576 24633
rect 30558 24624 30564 24636
rect 30616 24624 30622 24676
rect 33870 24624 33876 24676
rect 33928 24664 33934 24676
rect 35345 24667 35403 24673
rect 35345 24664 35357 24667
rect 33928 24636 35357 24664
rect 33928 24624 33934 24636
rect 35345 24633 35357 24636
rect 35391 24664 35403 24667
rect 35897 24667 35955 24673
rect 35897 24664 35909 24667
rect 35391 24636 35909 24664
rect 35391 24633 35403 24636
rect 35345 24627 35403 24633
rect 35897 24633 35909 24636
rect 35943 24633 35955 24667
rect 35897 24627 35955 24633
rect 8754 24596 8760 24608
rect 8715 24568 8760 24596
rect 8754 24556 8760 24568
rect 8812 24556 8818 24608
rect 11514 24596 11520 24608
rect 11475 24568 11520 24596
rect 11514 24556 11520 24568
rect 11572 24556 11578 24608
rect 12158 24596 12164 24608
rect 12119 24568 12164 24596
rect 12158 24556 12164 24568
rect 12216 24556 12222 24608
rect 12526 24556 12532 24608
rect 12584 24596 12590 24608
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 12584 24568 12817 24596
rect 12584 24556 12590 24568
rect 12805 24565 12817 24568
rect 12851 24565 12863 24599
rect 14090 24596 14096 24608
rect 14051 24568 14096 24596
rect 12805 24559 12863 24565
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 15654 24556 15660 24608
rect 15712 24596 15718 24608
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 15712 24568 16221 24596
rect 15712 24556 15718 24568
rect 16209 24565 16221 24568
rect 16255 24565 16267 24599
rect 17770 24596 17776 24608
rect 17731 24568 17776 24596
rect 16209 24559 16267 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 18690 24596 18696 24608
rect 18651 24568 18696 24596
rect 18690 24556 18696 24568
rect 18748 24556 18754 24608
rect 25866 24596 25872 24608
rect 25827 24568 25872 24596
rect 25866 24556 25872 24568
rect 25924 24556 25930 24608
rect 28166 24556 28172 24608
rect 28224 24596 28230 24608
rect 28261 24599 28319 24605
rect 28261 24596 28273 24599
rect 28224 24568 28273 24596
rect 28224 24556 28230 24568
rect 28261 24565 28273 24568
rect 28307 24596 28319 24599
rect 31481 24599 31539 24605
rect 31481 24596 31493 24599
rect 28307 24568 31493 24596
rect 28307 24565 28319 24568
rect 28261 24559 28319 24565
rect 31481 24565 31493 24568
rect 31527 24565 31539 24599
rect 31846 24596 31852 24608
rect 31807 24568 31852 24596
rect 31481 24559 31539 24565
rect 31846 24556 31852 24568
rect 31904 24556 31910 24608
rect 34790 24556 34796 24608
rect 34848 24596 34854 24608
rect 34885 24599 34943 24605
rect 34885 24596 34897 24599
rect 34848 24568 34897 24596
rect 34848 24556 34854 24568
rect 34885 24565 34897 24568
rect 34931 24565 34943 24599
rect 34885 24559 34943 24565
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 7190 24392 7196 24404
rect 7151 24364 7196 24392
rect 7190 24352 7196 24364
rect 7248 24352 7254 24404
rect 7834 24392 7840 24404
rect 7795 24364 7840 24392
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 10226 24392 10232 24404
rect 10187 24364 10232 24392
rect 10226 24352 10232 24364
rect 10284 24392 10290 24404
rect 11977 24395 12035 24401
rect 11977 24392 11989 24395
rect 10284 24364 11989 24392
rect 10284 24352 10290 24364
rect 11977 24361 11989 24364
rect 12023 24392 12035 24395
rect 12158 24392 12164 24404
rect 12023 24364 12164 24392
rect 12023 24361 12035 24364
rect 11977 24355 12035 24361
rect 12158 24352 12164 24364
rect 12216 24352 12222 24404
rect 14090 24352 14096 24404
rect 14148 24392 14154 24404
rect 15289 24395 15347 24401
rect 15289 24392 15301 24395
rect 14148 24364 15301 24392
rect 14148 24352 14154 24364
rect 15289 24361 15301 24364
rect 15335 24361 15347 24395
rect 15654 24392 15660 24404
rect 15615 24364 15660 24392
rect 15289 24355 15347 24361
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 15749 24395 15807 24401
rect 15749 24361 15761 24395
rect 15795 24392 15807 24395
rect 16482 24392 16488 24404
rect 15795 24364 16488 24392
rect 15795 24361 15807 24364
rect 15749 24355 15807 24361
rect 7208 24324 7236 24352
rect 7926 24324 7932 24336
rect 7208 24296 7932 24324
rect 7926 24284 7932 24296
rect 7984 24324 7990 24336
rect 8297 24327 8355 24333
rect 8297 24324 8309 24327
rect 7984 24296 8309 24324
rect 7984 24284 7990 24296
rect 8297 24293 8309 24296
rect 8343 24324 8355 24327
rect 8754 24324 8760 24336
rect 8343 24296 8760 24324
rect 8343 24293 8355 24296
rect 8297 24287 8355 24293
rect 8754 24284 8760 24296
rect 8812 24284 8818 24336
rect 10962 24284 10968 24336
rect 11020 24284 11026 24336
rect 11514 24284 11520 24336
rect 11572 24324 11578 24336
rect 12526 24324 12532 24336
rect 11572 24296 12532 24324
rect 11572 24284 11578 24296
rect 12526 24284 12532 24296
rect 12584 24284 12590 24336
rect 14921 24327 14979 24333
rect 14921 24293 14933 24327
rect 14967 24324 14979 24327
rect 15102 24324 15108 24336
rect 14967 24296 15108 24324
rect 14967 24293 14979 24296
rect 14921 24287 14979 24293
rect 15102 24284 15108 24296
rect 15160 24324 15166 24336
rect 15764 24324 15792 24355
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 16853 24395 16911 24401
rect 16853 24361 16865 24395
rect 16899 24392 16911 24395
rect 17770 24392 17776 24404
rect 16899 24364 17776 24392
rect 16899 24361 16911 24364
rect 16853 24355 16911 24361
rect 17770 24352 17776 24364
rect 17828 24352 17834 24404
rect 18049 24395 18107 24401
rect 18049 24361 18061 24395
rect 18095 24392 18107 24395
rect 18966 24392 18972 24404
rect 18095 24364 18972 24392
rect 18095 24361 18107 24364
rect 18049 24355 18107 24361
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 19978 24392 19984 24404
rect 19939 24364 19984 24392
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 20254 24392 20260 24404
rect 20215 24364 20260 24392
rect 20254 24352 20260 24364
rect 20312 24392 20318 24404
rect 20901 24395 20959 24401
rect 20901 24392 20913 24395
rect 20312 24364 20913 24392
rect 20312 24352 20318 24364
rect 20901 24361 20913 24364
rect 20947 24361 20959 24395
rect 24302 24392 24308 24404
rect 24263 24364 24308 24392
rect 20901 24355 20959 24361
rect 24302 24352 24308 24364
rect 24360 24352 24366 24404
rect 27249 24395 27307 24401
rect 27249 24361 27261 24395
rect 27295 24392 27307 24395
rect 27522 24392 27528 24404
rect 27295 24364 27528 24392
rect 27295 24361 27307 24364
rect 27249 24355 27307 24361
rect 27522 24352 27528 24364
rect 27580 24352 27586 24404
rect 29181 24395 29239 24401
rect 29181 24361 29193 24395
rect 29227 24392 29239 24395
rect 29362 24392 29368 24404
rect 29227 24364 29368 24392
rect 29227 24361 29239 24364
rect 29181 24355 29239 24361
rect 29362 24352 29368 24364
rect 29420 24352 29426 24404
rect 30558 24352 30564 24404
rect 30616 24392 30622 24404
rect 30653 24395 30711 24401
rect 30653 24392 30665 24395
rect 30616 24364 30665 24392
rect 30616 24352 30622 24364
rect 30653 24361 30665 24364
rect 30699 24361 30711 24395
rect 30653 24355 30711 24361
rect 30742 24352 30748 24404
rect 30800 24392 30806 24404
rect 31481 24395 31539 24401
rect 31481 24392 31493 24395
rect 30800 24364 31493 24392
rect 30800 24352 30806 24364
rect 31481 24361 31493 24364
rect 31527 24392 31539 24395
rect 31846 24392 31852 24404
rect 31527 24364 31852 24392
rect 31527 24361 31539 24364
rect 31481 24355 31539 24361
rect 31846 24352 31852 24364
rect 31904 24352 31910 24404
rect 31938 24352 31944 24404
rect 31996 24392 32002 24404
rect 32309 24395 32367 24401
rect 31996 24364 32041 24392
rect 31996 24352 32002 24364
rect 32309 24361 32321 24395
rect 32355 24392 32367 24395
rect 32858 24392 32864 24404
rect 32355 24364 32864 24392
rect 32355 24361 32367 24364
rect 32309 24355 32367 24361
rect 32858 24352 32864 24364
rect 32916 24352 32922 24404
rect 33042 24352 33048 24404
rect 33100 24392 33106 24404
rect 33505 24395 33563 24401
rect 33505 24392 33517 24395
rect 33100 24364 33517 24392
rect 33100 24352 33106 24364
rect 33505 24361 33517 24364
rect 33551 24392 33563 24395
rect 33686 24392 33692 24404
rect 33551 24364 33692 24392
rect 33551 24361 33563 24364
rect 33505 24355 33563 24361
rect 33686 24352 33692 24364
rect 33744 24352 33750 24404
rect 33873 24395 33931 24401
rect 33873 24361 33885 24395
rect 33919 24392 33931 24395
rect 34054 24392 34060 24404
rect 33919 24364 34060 24392
rect 33919 24361 33931 24364
rect 33873 24355 33931 24361
rect 34054 24352 34060 24364
rect 34112 24352 34118 24404
rect 36633 24395 36691 24401
rect 36633 24361 36645 24395
rect 36679 24392 36691 24395
rect 36906 24392 36912 24404
rect 36679 24364 36912 24392
rect 36679 24361 36691 24364
rect 36633 24355 36691 24361
rect 36906 24352 36912 24364
rect 36964 24352 36970 24404
rect 15160 24296 15792 24324
rect 17788 24324 17816 24352
rect 18325 24327 18383 24333
rect 18325 24324 18337 24327
rect 17788 24296 18337 24324
rect 15160 24284 15166 24296
rect 18325 24293 18337 24296
rect 18371 24293 18383 24327
rect 18325 24287 18383 24293
rect 19886 24284 19892 24336
rect 19944 24324 19950 24336
rect 20625 24327 20683 24333
rect 20625 24324 20637 24327
rect 19944 24296 20637 24324
rect 19944 24284 19950 24296
rect 20625 24293 20637 24296
rect 20671 24293 20683 24327
rect 20625 24287 20683 24293
rect 8202 24256 8208 24268
rect 8163 24228 8208 24256
rect 8202 24216 8208 24228
rect 8260 24216 8266 24268
rect 10686 24216 10692 24268
rect 10744 24256 10750 24268
rect 10853 24259 10911 24265
rect 10853 24256 10865 24259
rect 10744 24228 10865 24256
rect 10744 24216 10750 24228
rect 10853 24225 10865 24228
rect 10899 24256 10911 24259
rect 10980 24256 11008 24284
rect 10899 24228 11008 24256
rect 10899 24225 10911 24228
rect 10853 24219 10911 24225
rect 13262 24216 13268 24268
rect 13320 24256 13326 24268
rect 13630 24256 13636 24268
rect 13320 24228 13636 24256
rect 13320 24216 13326 24228
rect 13630 24216 13636 24228
rect 13688 24256 13694 24268
rect 14093 24259 14151 24265
rect 14093 24256 14105 24259
rect 13688 24228 14105 24256
rect 13688 24216 13694 24228
rect 14093 24225 14105 24228
rect 14139 24225 14151 24259
rect 14093 24219 14151 24225
rect 17221 24259 17279 24265
rect 17221 24225 17233 24259
rect 17267 24256 17279 24259
rect 17770 24256 17776 24268
rect 17267 24228 17776 24256
rect 17267 24225 17279 24228
rect 17221 24219 17279 24225
rect 17770 24216 17776 24228
rect 17828 24216 17834 24268
rect 18874 24265 18880 24268
rect 18868 24256 18880 24265
rect 18835 24228 18880 24256
rect 18868 24219 18880 24228
rect 18874 24216 18880 24219
rect 18932 24216 18938 24268
rect 20640 24256 20668 24287
rect 20714 24284 20720 24336
rect 20772 24324 20778 24336
rect 21269 24327 21327 24333
rect 21269 24324 21281 24327
rect 20772 24296 21281 24324
rect 20772 24284 20778 24296
rect 21269 24293 21281 24296
rect 21315 24293 21327 24327
rect 21269 24287 21327 24293
rect 23474 24284 23480 24336
rect 23532 24324 23538 24336
rect 24673 24327 24731 24333
rect 24673 24324 24685 24327
rect 23532 24296 24685 24324
rect 23532 24284 23538 24296
rect 24673 24293 24685 24296
rect 24719 24293 24731 24327
rect 24673 24287 24731 24293
rect 34508 24327 34566 24333
rect 34508 24293 34520 24327
rect 34554 24324 34566 24327
rect 35894 24324 35900 24336
rect 34554 24296 35900 24324
rect 34554 24293 34566 24296
rect 34508 24287 34566 24293
rect 35894 24284 35900 24296
rect 35952 24284 35958 24336
rect 20990 24256 20996 24268
rect 20640 24228 20996 24256
rect 20990 24216 20996 24228
rect 21048 24216 21054 24268
rect 24026 24216 24032 24268
rect 24084 24256 24090 24268
rect 24765 24259 24823 24265
rect 24765 24256 24777 24259
rect 24084 24228 24777 24256
rect 24084 24216 24090 24228
rect 24765 24225 24777 24228
rect 24811 24225 24823 24259
rect 27430 24256 27436 24268
rect 27391 24228 27436 24256
rect 24765 24219 24823 24225
rect 27430 24216 27436 24228
rect 27488 24216 27494 24268
rect 29546 24265 29552 24268
rect 29540 24219 29552 24265
rect 29604 24256 29610 24268
rect 29604 24228 29640 24256
rect 29546 24216 29552 24219
rect 29604 24216 29610 24228
rect 32030 24216 32036 24268
rect 32088 24256 32094 24268
rect 32125 24259 32183 24265
rect 32125 24256 32137 24259
rect 32088 24228 32137 24256
rect 32088 24216 32094 24228
rect 32125 24225 32137 24228
rect 32171 24225 32183 24259
rect 32125 24219 32183 24225
rect 34241 24259 34299 24265
rect 34241 24225 34253 24259
rect 34287 24256 34299 24259
rect 34882 24256 34888 24268
rect 34287 24228 34888 24256
rect 34287 24225 34299 24228
rect 34241 24219 34299 24225
rect 34882 24216 34888 24228
rect 34940 24256 34946 24268
rect 35526 24256 35532 24268
rect 34940 24228 35532 24256
rect 34940 24216 34946 24228
rect 35526 24216 35532 24228
rect 35584 24216 35590 24268
rect 36446 24256 36452 24268
rect 36407 24228 36452 24256
rect 36446 24216 36452 24228
rect 36504 24216 36510 24268
rect 8478 24188 8484 24200
rect 8439 24160 8484 24188
rect 8478 24148 8484 24160
rect 8536 24148 8542 24200
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10410 24188 10416 24200
rect 10192 24160 10416 24188
rect 10192 24148 10198 24160
rect 10410 24148 10416 24160
rect 10468 24188 10474 24200
rect 10597 24191 10655 24197
rect 10597 24188 10609 24191
rect 10468 24160 10609 24188
rect 10468 24148 10474 24160
rect 10597 24157 10609 24160
rect 10643 24157 10655 24191
rect 10597 24151 10655 24157
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 15746 24188 15752 24200
rect 15252 24160 15752 24188
rect 15252 24148 15258 24160
rect 15746 24148 15752 24160
rect 15804 24188 15810 24200
rect 15841 24191 15899 24197
rect 15841 24188 15853 24191
rect 15804 24160 15853 24188
rect 15804 24148 15810 24160
rect 15841 24157 15853 24160
rect 15887 24157 15899 24191
rect 17310 24188 17316 24200
rect 15841 24151 15899 24157
rect 16040 24160 17316 24188
rect 7374 24080 7380 24132
rect 7432 24120 7438 24132
rect 7561 24123 7619 24129
rect 7561 24120 7573 24123
rect 7432 24092 7573 24120
rect 7432 24080 7438 24092
rect 7561 24089 7573 24092
rect 7607 24120 7619 24123
rect 10152 24120 10180 24148
rect 7607 24092 10180 24120
rect 14277 24123 14335 24129
rect 7607 24089 7619 24092
rect 7561 24083 7619 24089
rect 14277 24089 14289 24123
rect 14323 24120 14335 24123
rect 16040 24120 16068 24160
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 17494 24188 17500 24200
rect 17455 24160 17500 24188
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 18598 24188 18604 24200
rect 18559 24160 18604 24188
rect 18598 24148 18604 24160
rect 18656 24148 18662 24200
rect 21358 24188 21364 24200
rect 21319 24160 21364 24188
rect 21358 24148 21364 24160
rect 21416 24148 21422 24200
rect 21450 24148 21456 24200
rect 21508 24188 21514 24200
rect 21508 24160 21553 24188
rect 21508 24148 21514 24160
rect 24210 24148 24216 24200
rect 24268 24188 24274 24200
rect 24857 24191 24915 24197
rect 24857 24188 24869 24191
rect 24268 24160 24869 24188
rect 24268 24148 24274 24160
rect 24857 24157 24869 24160
rect 24903 24188 24915 24191
rect 25866 24188 25872 24200
rect 24903 24160 25872 24188
rect 24903 24157 24915 24160
rect 24857 24151 24915 24157
rect 25866 24148 25872 24160
rect 25924 24148 25930 24200
rect 28994 24148 29000 24200
rect 29052 24188 29058 24200
rect 29273 24191 29331 24197
rect 29273 24188 29285 24191
rect 29052 24160 29285 24188
rect 29052 24148 29058 24160
rect 29273 24157 29285 24160
rect 29319 24157 29331 24191
rect 29273 24151 29331 24157
rect 14323 24092 16068 24120
rect 16485 24123 16543 24129
rect 14323 24089 14335 24092
rect 14277 24083 14335 24089
rect 16485 24089 16497 24123
rect 16531 24120 16543 24123
rect 16942 24120 16948 24132
rect 16531 24092 16948 24120
rect 16531 24089 16543 24092
rect 16485 24083 16543 24089
rect 16942 24080 16948 24092
rect 17000 24080 17006 24132
rect 13725 24055 13783 24061
rect 13725 24021 13737 24055
rect 13771 24052 13783 24055
rect 14458 24052 14464 24064
rect 13771 24024 14464 24052
rect 13771 24021 13783 24024
rect 13725 24015 13783 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 25130 24012 25136 24064
rect 25188 24052 25194 24064
rect 25317 24055 25375 24061
rect 25317 24052 25329 24055
rect 25188 24024 25329 24052
rect 25188 24012 25194 24024
rect 25317 24021 25329 24024
rect 25363 24021 25375 24055
rect 35618 24052 35624 24064
rect 35579 24024 35624 24052
rect 25317 24015 25375 24021
rect 35618 24012 35624 24024
rect 35676 24012 35682 24064
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 7926 23848 7932 23860
rect 7887 23820 7932 23848
rect 7926 23808 7932 23820
rect 7984 23808 7990 23860
rect 8202 23848 8208 23860
rect 8163 23820 8208 23848
rect 8202 23808 8208 23820
rect 8260 23808 8266 23860
rect 8478 23808 8484 23860
rect 8536 23848 8542 23860
rect 8573 23851 8631 23857
rect 8573 23848 8585 23851
rect 8536 23820 8585 23848
rect 8536 23808 8542 23820
rect 8573 23817 8585 23820
rect 8619 23817 8631 23851
rect 10686 23848 10692 23860
rect 10647 23820 10692 23848
rect 8573 23811 8631 23817
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 10778 23808 10784 23860
rect 10836 23848 10842 23860
rect 11333 23851 11391 23857
rect 11333 23848 11345 23851
rect 10836 23820 11345 23848
rect 10836 23808 10842 23820
rect 11333 23817 11345 23820
rect 11379 23817 11391 23851
rect 13262 23848 13268 23860
rect 13223 23820 13268 23848
rect 11333 23811 11391 23817
rect 13262 23808 13268 23820
rect 13320 23808 13326 23860
rect 15102 23808 15108 23860
rect 15160 23848 15166 23860
rect 15381 23851 15439 23857
rect 15381 23848 15393 23851
rect 15160 23820 15393 23848
rect 15160 23808 15166 23820
rect 15381 23817 15393 23820
rect 15427 23817 15439 23851
rect 15381 23811 15439 23817
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 15749 23851 15807 23857
rect 15749 23848 15761 23851
rect 15712 23820 15761 23848
rect 15712 23808 15718 23820
rect 15749 23817 15761 23820
rect 15795 23817 15807 23851
rect 16390 23848 16396 23860
rect 16351 23820 16396 23848
rect 15749 23811 15807 23817
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 17310 23808 17316 23860
rect 17368 23848 17374 23860
rect 17405 23851 17463 23857
rect 17405 23848 17417 23851
rect 17368 23820 17417 23848
rect 17368 23808 17374 23820
rect 17405 23817 17417 23820
rect 17451 23817 17463 23851
rect 17770 23848 17776 23860
rect 17731 23820 17776 23848
rect 17405 23811 17463 23817
rect 17770 23808 17776 23820
rect 17828 23848 17834 23860
rect 18233 23851 18291 23857
rect 18233 23848 18245 23851
rect 17828 23820 18245 23848
rect 17828 23808 17834 23820
rect 18233 23817 18245 23820
rect 18279 23817 18291 23851
rect 18233 23811 18291 23817
rect 19334 23808 19340 23860
rect 19392 23848 19398 23860
rect 19613 23851 19671 23857
rect 19613 23848 19625 23851
rect 19392 23820 19625 23848
rect 19392 23808 19398 23820
rect 19613 23817 19625 23820
rect 19659 23817 19671 23851
rect 19978 23848 19984 23860
rect 19939 23820 19984 23848
rect 19613 23811 19671 23817
rect 19978 23808 19984 23820
rect 20036 23808 20042 23860
rect 20714 23848 20720 23860
rect 20675 23820 20720 23848
rect 20714 23808 20720 23820
rect 20772 23808 20778 23860
rect 22002 23808 22008 23860
rect 22060 23848 22066 23860
rect 22097 23851 22155 23857
rect 22097 23848 22109 23851
rect 22060 23820 22109 23848
rect 22060 23808 22066 23820
rect 22097 23817 22109 23820
rect 22143 23817 22155 23851
rect 22097 23811 22155 23817
rect 23474 23808 23480 23860
rect 23532 23848 23538 23860
rect 24121 23851 24179 23857
rect 24121 23848 24133 23851
rect 23532 23820 24133 23848
rect 23532 23808 23538 23820
rect 24121 23817 24133 23820
rect 24167 23817 24179 23851
rect 24121 23811 24179 23817
rect 24578 23808 24584 23860
rect 24636 23848 24642 23860
rect 24673 23851 24731 23857
rect 24673 23848 24685 23851
rect 24636 23820 24685 23848
rect 24636 23808 24642 23820
rect 24673 23817 24685 23820
rect 24719 23817 24731 23851
rect 24673 23811 24731 23817
rect 27341 23851 27399 23857
rect 27341 23817 27353 23851
rect 27387 23848 27399 23851
rect 27430 23848 27436 23860
rect 27387 23820 27436 23848
rect 27387 23817 27399 23820
rect 27341 23811 27399 23817
rect 27430 23808 27436 23820
rect 27488 23848 27494 23860
rect 28074 23848 28080 23860
rect 27488 23820 28080 23848
rect 27488 23808 27494 23820
rect 28074 23808 28080 23820
rect 28132 23848 28138 23860
rect 28721 23851 28779 23857
rect 28721 23848 28733 23851
rect 28132 23820 28733 23848
rect 28132 23808 28138 23820
rect 28721 23817 28733 23820
rect 28767 23817 28779 23851
rect 28902 23848 28908 23860
rect 28863 23820 28908 23848
rect 28721 23811 28779 23817
rect 10410 23740 10416 23792
rect 10468 23780 10474 23792
rect 11057 23783 11115 23789
rect 11057 23780 11069 23783
rect 10468 23752 11069 23780
rect 10468 23740 10474 23752
rect 11057 23749 11069 23752
rect 11103 23780 11115 23783
rect 11790 23780 11796 23792
rect 11103 23752 11796 23780
rect 11103 23749 11115 23752
rect 11057 23743 11115 23749
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 15933 23783 15991 23789
rect 15933 23749 15945 23783
rect 15979 23780 15991 23783
rect 15979 23752 17448 23780
rect 15979 23749 15991 23752
rect 15933 23743 15991 23749
rect 17420 23724 17448 23752
rect 18782 23740 18788 23792
rect 18840 23780 18846 23792
rect 20257 23783 20315 23789
rect 20257 23780 20269 23783
rect 18840 23752 20269 23780
rect 18840 23740 18846 23752
rect 20257 23749 20269 23752
rect 20303 23780 20315 23783
rect 21358 23780 21364 23792
rect 20303 23752 21364 23780
rect 20303 23749 20315 23752
rect 20257 23743 20315 23749
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 26421 23783 26479 23789
rect 26421 23749 26433 23783
rect 26467 23780 26479 23783
rect 27522 23780 27528 23792
rect 26467 23752 27528 23780
rect 26467 23749 26479 23752
rect 26421 23743 26479 23749
rect 13633 23715 13691 23721
rect 13633 23681 13645 23715
rect 13679 23712 13691 23715
rect 17037 23715 17095 23721
rect 13679 23684 13860 23712
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 11517 23647 11575 23653
rect 11517 23644 11529 23647
rect 11112 23616 11529 23644
rect 11112 23604 11118 23616
rect 11517 23613 11529 23616
rect 11563 23644 11575 23647
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11563 23616 11805 23644
rect 11563 23613 11575 23616
rect 11517 23607 11575 23613
rect 11793 23613 11805 23616
rect 11839 23644 11851 23647
rect 12342 23644 12348 23656
rect 11839 23616 12348 23644
rect 11839 23613 11851 23616
rect 11793 23607 11851 23613
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12897 23647 12955 23653
rect 12897 23613 12909 23647
rect 12943 23644 12955 23647
rect 13725 23647 13783 23653
rect 13725 23644 13737 23647
rect 12943 23616 13737 23644
rect 12943 23613 12955 23616
rect 12897 23607 12955 23613
rect 13725 23613 13737 23616
rect 13771 23613 13783 23647
rect 13832 23644 13860 23684
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 17037 23675 17095 23681
rect 13992 23647 14050 23653
rect 13992 23644 14004 23647
rect 13832 23616 14004 23644
rect 13725 23607 13783 23613
rect 13992 23613 14004 23616
rect 14038 23644 14050 23647
rect 15654 23644 15660 23656
rect 14038 23616 15660 23644
rect 14038 23613 14050 23616
rect 13992 23607 14050 23613
rect 13740 23576 13768 23607
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 16117 23647 16175 23653
rect 16117 23613 16129 23647
rect 16163 23644 16175 23647
rect 16482 23644 16488 23656
rect 16163 23616 16488 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 16482 23604 16488 23616
rect 16540 23604 16546 23656
rect 17052 23644 17080 23675
rect 17402 23672 17408 23724
rect 17460 23672 17466 23724
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23712 23535 23715
rect 24026 23712 24032 23724
rect 23523 23684 24032 23712
rect 23523 23681 23535 23684
rect 23477 23675 23535 23681
rect 24026 23672 24032 23684
rect 24084 23672 24090 23724
rect 26436 23712 26464 23743
rect 27522 23740 27528 23752
rect 27580 23740 27586 23792
rect 24872 23684 26464 23712
rect 17494 23644 17500 23656
rect 17052 23616 17500 23644
rect 17494 23604 17500 23616
rect 17552 23604 17558 23656
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 18046 23604 18052 23616
rect 18104 23644 18110 23656
rect 18601 23647 18659 23653
rect 18601 23644 18613 23647
rect 18104 23616 18613 23644
rect 18104 23604 18110 23616
rect 18601 23613 18613 23616
rect 18647 23613 18659 23647
rect 18601 23607 18659 23613
rect 19153 23647 19211 23653
rect 19153 23613 19165 23647
rect 19199 23644 19211 23647
rect 19426 23644 19432 23656
rect 19199 23616 19432 23644
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 19426 23604 19432 23616
rect 19484 23604 19490 23656
rect 24872 23653 24900 23684
rect 24857 23647 24915 23653
rect 24857 23613 24869 23647
rect 24903 23613 24915 23647
rect 25130 23644 25136 23656
rect 25091 23616 25136 23644
rect 24857 23607 24915 23613
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 25409 23647 25467 23653
rect 25409 23644 25421 23647
rect 25240 23616 25421 23644
rect 14734 23576 14740 23588
rect 13740 23548 14740 23576
rect 14734 23536 14740 23548
rect 14792 23536 14798 23588
rect 16761 23579 16819 23585
rect 16761 23545 16773 23579
rect 16807 23576 16819 23579
rect 16942 23576 16948 23588
rect 16807 23548 16948 23576
rect 16807 23545 16819 23548
rect 16761 23539 16819 23545
rect 16942 23536 16948 23548
rect 17000 23536 17006 23588
rect 19245 23579 19303 23585
rect 19245 23545 19257 23579
rect 19291 23576 19303 23579
rect 19978 23576 19984 23588
rect 19291 23548 19984 23576
rect 19291 23545 19303 23548
rect 19245 23539 19303 23545
rect 19978 23536 19984 23548
rect 20036 23536 20042 23588
rect 20809 23579 20867 23585
rect 20809 23545 20821 23579
rect 20855 23576 20867 23579
rect 21542 23576 21548 23588
rect 20855 23548 21548 23576
rect 20855 23545 20867 23548
rect 20809 23539 20867 23545
rect 21542 23536 21548 23548
rect 21600 23536 21606 23588
rect 24581 23579 24639 23585
rect 24581 23545 24593 23579
rect 24627 23576 24639 23579
rect 24949 23579 25007 23585
rect 24949 23576 24961 23579
rect 24627 23548 24961 23576
rect 24627 23545 24639 23548
rect 24581 23539 24639 23545
rect 24949 23545 24961 23548
rect 24995 23576 25007 23579
rect 25038 23576 25044 23588
rect 24995 23548 25044 23576
rect 24995 23545 25007 23548
rect 24949 23539 25007 23545
rect 25038 23536 25044 23548
rect 25096 23536 25102 23588
rect 14366 23468 14372 23520
rect 14424 23508 14430 23520
rect 15105 23511 15163 23517
rect 15105 23508 15117 23511
rect 14424 23480 15117 23508
rect 14424 23468 14430 23480
rect 15105 23477 15117 23480
rect 15151 23477 15163 23511
rect 15105 23471 15163 23477
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 16853 23511 16911 23517
rect 16853 23508 16865 23511
rect 16632 23480 16865 23508
rect 16632 23468 16638 23480
rect 16853 23477 16865 23480
rect 16899 23477 16911 23511
rect 16853 23471 16911 23477
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 25240 23508 25268 23616
rect 25409 23613 25421 23616
rect 25455 23644 25467 23647
rect 25961 23647 26019 23653
rect 25961 23644 25973 23647
rect 25455 23616 25973 23644
rect 25455 23613 25467 23616
rect 25409 23607 25467 23613
rect 25961 23613 25973 23616
rect 26007 23613 26019 23647
rect 28736 23644 28764 23811
rect 28902 23808 28908 23820
rect 28960 23808 28966 23860
rect 29546 23848 29552 23860
rect 29507 23820 29552 23848
rect 29546 23808 29552 23820
rect 29604 23848 29610 23860
rect 31294 23848 31300 23860
rect 29604 23820 30420 23848
rect 31255 23820 31300 23848
rect 29604 23808 29610 23820
rect 28810 23740 28816 23792
rect 28868 23780 28874 23792
rect 29917 23783 29975 23789
rect 29917 23780 29929 23783
rect 28868 23752 29929 23780
rect 28868 23740 28874 23752
rect 29917 23749 29929 23752
rect 29963 23749 29975 23783
rect 29917 23743 29975 23749
rect 30392 23780 30420 23820
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 32030 23808 32036 23860
rect 32088 23848 32094 23860
rect 32125 23851 32183 23857
rect 32125 23848 32137 23851
rect 32088 23820 32137 23848
rect 32088 23808 32094 23820
rect 32125 23817 32137 23820
rect 32171 23817 32183 23851
rect 32766 23848 32772 23860
rect 32727 23820 32772 23848
rect 32125 23811 32183 23817
rect 32766 23808 32772 23820
rect 32824 23808 32830 23860
rect 33134 23848 33140 23860
rect 33095 23820 33140 23848
rect 33134 23808 33140 23820
rect 33192 23808 33198 23860
rect 33410 23808 33416 23860
rect 33468 23848 33474 23860
rect 33505 23851 33563 23857
rect 33505 23848 33517 23851
rect 33468 23820 33517 23848
rect 33468 23808 33474 23820
rect 33505 23817 33517 23820
rect 33551 23817 33563 23851
rect 33870 23848 33876 23860
rect 33831 23820 33876 23848
rect 33505 23811 33563 23817
rect 30929 23783 30987 23789
rect 30929 23780 30941 23783
rect 30392 23752 30941 23780
rect 30282 23672 30288 23724
rect 30340 23712 30346 23724
rect 30392 23721 30420 23752
rect 30929 23749 30941 23752
rect 30975 23749 30987 23783
rect 30929 23743 30987 23749
rect 30377 23715 30435 23721
rect 30377 23712 30389 23715
rect 30340 23684 30389 23712
rect 30340 23672 30346 23684
rect 30377 23681 30389 23684
rect 30423 23681 30435 23715
rect 30377 23675 30435 23681
rect 30561 23715 30619 23721
rect 30561 23681 30573 23715
rect 30607 23712 30619 23715
rect 31312 23712 31340 23808
rect 30607 23684 31340 23712
rect 30607 23681 30619 23684
rect 30561 23675 30619 23681
rect 29089 23647 29147 23653
rect 29089 23644 29101 23647
rect 28736 23616 29101 23644
rect 25961 23607 26019 23613
rect 29089 23613 29101 23616
rect 29135 23613 29147 23647
rect 29089 23607 29147 23613
rect 32585 23647 32643 23653
rect 32585 23613 32597 23647
rect 32631 23644 32643 23647
rect 33134 23644 33140 23656
rect 32631 23616 33140 23644
rect 32631 23613 32643 23616
rect 32585 23607 32643 23613
rect 33134 23604 33140 23616
rect 33192 23604 33198 23656
rect 33520 23644 33548 23811
rect 33870 23808 33876 23820
rect 33928 23808 33934 23860
rect 35894 23848 35900 23860
rect 35855 23820 35900 23848
rect 35894 23808 35900 23820
rect 35952 23808 35958 23860
rect 36446 23848 36452 23860
rect 36407 23820 36452 23848
rect 36446 23808 36452 23820
rect 36504 23808 36510 23860
rect 34333 23715 34391 23721
rect 34333 23681 34345 23715
rect 34379 23712 34391 23715
rect 34422 23712 34428 23724
rect 34379 23684 34428 23712
rect 34379 23681 34391 23684
rect 34333 23675 34391 23681
rect 34422 23672 34428 23684
rect 34480 23712 34486 23724
rect 35529 23715 35587 23721
rect 35529 23712 35541 23715
rect 34480 23684 35541 23712
rect 34480 23672 34486 23684
rect 35529 23681 35541 23684
rect 35575 23712 35587 23715
rect 35618 23712 35624 23724
rect 35575 23684 35624 23712
rect 35575 23681 35587 23684
rect 35529 23675 35587 23681
rect 35618 23672 35624 23684
rect 35676 23672 35682 23724
rect 33689 23647 33747 23653
rect 33689 23644 33701 23647
rect 33520 23616 33701 23644
rect 33689 23613 33701 23616
rect 33735 23613 33747 23647
rect 33689 23607 33747 23613
rect 34514 23604 34520 23656
rect 34572 23644 34578 23656
rect 34790 23644 34796 23656
rect 34572 23616 34796 23644
rect 34572 23604 34578 23616
rect 34790 23604 34796 23616
rect 34848 23644 34854 23656
rect 35345 23647 35403 23653
rect 35345 23644 35357 23647
rect 34848 23616 35357 23644
rect 34848 23604 34854 23616
rect 35345 23613 35357 23616
rect 35391 23613 35403 23647
rect 35345 23607 35403 23613
rect 25317 23579 25375 23585
rect 25317 23545 25329 23579
rect 25363 23576 25375 23579
rect 26142 23576 26148 23588
rect 25363 23548 26148 23576
rect 25363 23545 25375 23548
rect 25317 23539 25375 23545
rect 26142 23536 26148 23548
rect 26200 23536 26206 23588
rect 30285 23579 30343 23585
rect 30285 23545 30297 23579
rect 30331 23576 30343 23579
rect 30558 23576 30564 23588
rect 30331 23548 30564 23576
rect 30331 23545 30343 23548
rect 30285 23539 30343 23545
rect 30558 23536 30564 23548
rect 30616 23536 30622 23588
rect 34701 23579 34759 23585
rect 34701 23545 34713 23579
rect 34747 23576 34759 23579
rect 35253 23579 35311 23585
rect 35253 23576 35265 23579
rect 34747 23548 35265 23576
rect 34747 23545 34759 23548
rect 34701 23539 34759 23545
rect 35253 23545 35265 23548
rect 35299 23576 35311 23579
rect 35986 23576 35992 23588
rect 35299 23548 35992 23576
rect 35299 23545 35311 23548
rect 35253 23539 35311 23545
rect 35986 23536 35992 23548
rect 36044 23536 36050 23588
rect 25590 23508 25596 23520
rect 24912 23480 25268 23508
rect 25551 23480 25596 23508
rect 24912 23468 24918 23480
rect 25590 23468 25596 23480
rect 25648 23468 25654 23520
rect 28445 23511 28503 23517
rect 28445 23477 28457 23511
rect 28491 23508 28503 23511
rect 28902 23508 28908 23520
rect 28491 23480 28908 23508
rect 28491 23477 28503 23480
rect 28445 23471 28503 23477
rect 28902 23468 28908 23480
rect 28960 23468 28966 23520
rect 34238 23468 34244 23520
rect 34296 23508 34302 23520
rect 34885 23511 34943 23517
rect 34885 23508 34897 23511
rect 34296 23480 34897 23508
rect 34296 23468 34302 23480
rect 34885 23477 34897 23480
rect 34931 23477 34943 23511
rect 34885 23471 34943 23477
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 10410 23304 10416 23316
rect 10371 23276 10416 23304
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 12529 23307 12587 23313
rect 12529 23304 12541 23307
rect 12492 23276 12541 23304
rect 12492 23264 12498 23276
rect 12529 23273 12541 23276
rect 12575 23273 12587 23307
rect 15102 23304 15108 23316
rect 15063 23276 15108 23304
rect 12529 23267 12587 23273
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15286 23304 15292 23316
rect 15247 23276 15292 23304
rect 15286 23264 15292 23276
rect 15344 23264 15350 23316
rect 18785 23307 18843 23313
rect 18785 23273 18797 23307
rect 18831 23304 18843 23307
rect 18874 23304 18880 23316
rect 18831 23276 18880 23304
rect 18831 23273 18843 23276
rect 18785 23267 18843 23273
rect 18874 23264 18880 23276
rect 18932 23304 18938 23316
rect 20533 23307 20591 23313
rect 20533 23304 20545 23307
rect 18932 23276 20545 23304
rect 18932 23264 18938 23276
rect 20533 23273 20545 23276
rect 20579 23304 20591 23307
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 20579 23276 21189 23304
rect 20579 23273 20591 23276
rect 20533 23267 20591 23273
rect 21177 23273 21189 23276
rect 21223 23304 21235 23307
rect 21450 23304 21456 23316
rect 21223 23276 21456 23304
rect 21223 23273 21235 23276
rect 21177 23267 21235 23273
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 28074 23304 28080 23316
rect 28035 23276 28080 23304
rect 28074 23264 28080 23276
rect 28132 23264 28138 23316
rect 30282 23304 30288 23316
rect 30243 23276 30288 23304
rect 30282 23264 30288 23276
rect 30340 23264 30346 23316
rect 30558 23304 30564 23316
rect 30519 23276 30564 23304
rect 30558 23264 30564 23276
rect 30616 23264 30622 23316
rect 34057 23307 34115 23313
rect 34057 23273 34069 23307
rect 34103 23304 34115 23307
rect 34514 23304 34520 23316
rect 34103 23276 34520 23304
rect 34103 23273 34115 23276
rect 34057 23267 34115 23273
rect 34514 23264 34520 23276
rect 34572 23264 34578 23316
rect 35526 23264 35532 23316
rect 35584 23304 35590 23316
rect 35805 23307 35863 23313
rect 35805 23304 35817 23307
rect 35584 23276 35817 23304
rect 35584 23264 35590 23276
rect 35805 23273 35817 23276
rect 35851 23273 35863 23307
rect 35805 23267 35863 23273
rect 35986 23264 35992 23316
rect 36044 23304 36050 23316
rect 36357 23307 36415 23313
rect 36357 23304 36369 23307
rect 36044 23276 36369 23304
rect 36044 23264 36050 23276
rect 36357 23273 36369 23276
rect 36403 23273 36415 23307
rect 36357 23267 36415 23273
rect 19426 23245 19432 23248
rect 19420 23236 19432 23245
rect 19387 23208 19432 23236
rect 19420 23199 19432 23208
rect 19426 23196 19432 23199
rect 19484 23196 19490 23248
rect 24940 23239 24998 23245
rect 24940 23205 24952 23239
rect 24986 23236 24998 23239
rect 25130 23236 25136 23248
rect 24986 23208 25136 23236
rect 24986 23205 24998 23208
rect 24940 23199 24998 23205
rect 25130 23196 25136 23208
rect 25188 23196 25194 23248
rect 33594 23196 33600 23248
rect 33652 23236 33658 23248
rect 33689 23239 33747 23245
rect 33689 23236 33701 23239
rect 33652 23208 33701 23236
rect 33652 23196 33658 23208
rect 33689 23205 33701 23208
rect 33735 23236 33747 23239
rect 34238 23236 34244 23248
rect 33735 23208 34244 23236
rect 33735 23205 33747 23208
rect 33689 23199 33747 23205
rect 34238 23196 34244 23208
rect 34296 23196 34302 23248
rect 34422 23245 34428 23248
rect 34416 23236 34428 23245
rect 34383 23208 34428 23236
rect 34416 23199 34428 23208
rect 34422 23196 34428 23199
rect 34480 23196 34486 23248
rect 10502 23128 10508 23180
rect 10560 23168 10566 23180
rect 10597 23171 10655 23177
rect 10597 23168 10609 23171
rect 10560 23140 10609 23168
rect 10560 23128 10566 23140
rect 10597 23137 10609 23140
rect 10643 23168 10655 23171
rect 11054 23168 11060 23180
rect 10643 23140 11060 23168
rect 10643 23137 10655 23140
rect 10597 23131 10655 23137
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 12710 23168 12716 23180
rect 12671 23140 12716 23168
rect 12710 23128 12716 23140
rect 12768 23128 12774 23180
rect 13262 23177 13268 23180
rect 13256 23168 13268 23177
rect 13223 23140 13268 23168
rect 13256 23131 13268 23140
rect 13262 23128 13268 23131
rect 13320 23128 13326 23180
rect 15654 23168 15660 23180
rect 15615 23140 15660 23168
rect 15654 23128 15660 23140
rect 15712 23128 15718 23180
rect 17221 23171 17279 23177
rect 17221 23137 17233 23171
rect 17267 23168 17279 23171
rect 17586 23168 17592 23180
rect 17267 23140 17592 23168
rect 17267 23137 17279 23140
rect 17221 23131 17279 23137
rect 17586 23128 17592 23140
rect 17644 23128 17650 23180
rect 18598 23128 18604 23180
rect 18656 23168 18662 23180
rect 19153 23171 19211 23177
rect 19153 23168 19165 23171
rect 18656 23140 19165 23168
rect 18656 23128 18662 23140
rect 19153 23137 19165 23140
rect 19199 23137 19211 23171
rect 24670 23168 24676 23180
rect 24631 23140 24676 23168
rect 19153 23131 19211 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 27798 23128 27804 23180
rect 27856 23168 27862 23180
rect 29178 23177 29184 23180
rect 28261 23171 28319 23177
rect 28261 23168 28273 23171
rect 27856 23140 28273 23168
rect 27856 23128 27862 23140
rect 28261 23137 28273 23140
rect 28307 23137 28319 23171
rect 29172 23168 29184 23177
rect 29139 23140 29184 23168
rect 28261 23131 28319 23137
rect 29172 23131 29184 23140
rect 29178 23128 29184 23131
rect 29236 23128 29242 23180
rect 33042 23168 33048 23180
rect 33003 23140 33048 23168
rect 33042 23128 33048 23140
rect 33100 23128 33106 23180
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23069 13047 23103
rect 12989 23063 13047 23069
rect 12437 22967 12495 22973
rect 12437 22933 12449 22967
rect 12483 22964 12495 22967
rect 13004 22964 13032 23063
rect 15378 23060 15384 23112
rect 15436 23100 15442 23112
rect 15749 23103 15807 23109
rect 15749 23100 15761 23103
rect 15436 23072 15761 23100
rect 15436 23060 15442 23072
rect 15749 23069 15761 23072
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 15933 23103 15991 23109
rect 15933 23069 15945 23103
rect 15979 23069 15991 23103
rect 17310 23100 17316 23112
rect 17271 23072 17316 23100
rect 15933 23063 15991 23069
rect 14458 22992 14464 23044
rect 14516 23032 14522 23044
rect 14737 23035 14795 23041
rect 14737 23032 14749 23035
rect 14516 23004 14749 23032
rect 14516 22992 14522 23004
rect 14737 23001 14749 23004
rect 14783 23032 14795 23035
rect 15010 23032 15016 23044
rect 14783 23004 15016 23032
rect 14783 23001 14795 23004
rect 14737 22995 14795 23001
rect 15010 22992 15016 23004
rect 15068 23032 15074 23044
rect 15948 23032 15976 23063
rect 17310 23060 17316 23072
rect 17368 23060 17374 23112
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23100 17463 23103
rect 17865 23103 17923 23109
rect 17865 23100 17877 23103
rect 17451 23072 17877 23100
rect 17451 23069 17463 23072
rect 17405 23063 17463 23069
rect 17865 23069 17877 23072
rect 17911 23069 17923 23103
rect 28902 23100 28908 23112
rect 28863 23072 28908 23100
rect 17865 23063 17923 23069
rect 16022 23032 16028 23044
rect 15068 23004 16028 23032
rect 15068 22992 15074 23004
rect 16022 22992 16028 23004
rect 16080 23032 16086 23044
rect 17218 23032 17224 23044
rect 16080 23004 17224 23032
rect 16080 22992 16086 23004
rect 17218 22992 17224 23004
rect 17276 23032 17282 23044
rect 17420 23032 17448 23063
rect 28902 23060 28908 23072
rect 28960 23060 28966 23112
rect 31202 23060 31208 23112
rect 31260 23100 31266 23112
rect 34054 23100 34060 23112
rect 31260 23072 34060 23100
rect 31260 23060 31266 23072
rect 34054 23060 34060 23072
rect 34112 23100 34118 23112
rect 34149 23103 34207 23109
rect 34149 23100 34161 23103
rect 34112 23072 34161 23100
rect 34112 23060 34118 23072
rect 34149 23069 34161 23072
rect 34195 23069 34207 23103
rect 34149 23063 34207 23069
rect 17276 23004 17448 23032
rect 17276 22992 17282 23004
rect 13630 22964 13636 22976
rect 12483 22936 13636 22964
rect 12483 22933 12495 22936
rect 12437 22927 12495 22933
rect 13630 22924 13636 22936
rect 13688 22924 13694 22976
rect 14274 22924 14280 22976
rect 14332 22964 14338 22976
rect 14369 22967 14427 22973
rect 14369 22964 14381 22967
rect 14332 22936 14381 22964
rect 14332 22924 14338 22936
rect 14369 22933 14381 22936
rect 14415 22933 14427 22967
rect 16390 22964 16396 22976
rect 16351 22936 16396 22964
rect 14369 22927 14427 22933
rect 16390 22924 16396 22936
rect 16448 22924 16454 22976
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 16853 22967 16911 22973
rect 16853 22964 16865 22967
rect 16724 22936 16865 22964
rect 16724 22924 16730 22936
rect 16853 22933 16865 22936
rect 16899 22933 16911 22967
rect 18414 22964 18420 22976
rect 18375 22936 18420 22964
rect 16853 22927 16911 22933
rect 18414 22924 18420 22936
rect 18472 22924 18478 22976
rect 21542 22964 21548 22976
rect 21503 22936 21548 22964
rect 21542 22924 21548 22936
rect 21600 22924 21606 22976
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 22152 22936 22197 22964
rect 22152 22924 22158 22936
rect 24210 22924 24216 22976
rect 24268 22964 24274 22976
rect 24305 22967 24363 22973
rect 24305 22964 24317 22967
rect 24268 22936 24317 22964
rect 24268 22924 24274 22936
rect 24305 22933 24317 22936
rect 24351 22933 24363 22967
rect 24305 22927 24363 22933
rect 25866 22924 25872 22976
rect 25924 22964 25930 22976
rect 26053 22967 26111 22973
rect 26053 22964 26065 22967
rect 25924 22936 26065 22964
rect 25924 22924 25930 22936
rect 26053 22933 26065 22936
rect 26099 22933 26111 22967
rect 33226 22964 33232 22976
rect 33187 22936 33232 22964
rect 26053 22927 26111 22933
rect 33226 22924 33232 22936
rect 33284 22924 33290 22976
rect 35526 22964 35532 22976
rect 35487 22936 35532 22964
rect 35526 22924 35532 22936
rect 35584 22924 35590 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 10502 22760 10508 22772
rect 10463 22732 10508 22760
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 12253 22763 12311 22769
rect 12253 22729 12265 22763
rect 12299 22760 12311 22763
rect 12618 22760 12624 22772
rect 12299 22732 12624 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 12986 22760 12992 22772
rect 12947 22732 12992 22760
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 13909 22763 13967 22769
rect 13909 22729 13921 22763
rect 13955 22760 13967 22763
rect 15378 22760 15384 22772
rect 13955 22732 15384 22760
rect 13955 22729 13967 22732
rect 13909 22723 13967 22729
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 15654 22720 15660 22772
rect 15712 22760 15718 22772
rect 16485 22763 16543 22769
rect 16485 22760 16497 22763
rect 15712 22732 16497 22760
rect 15712 22720 15718 22732
rect 16485 22729 16497 22732
rect 16531 22729 16543 22763
rect 17310 22760 17316 22772
rect 17271 22732 17316 22760
rect 16485 22723 16543 22729
rect 17310 22720 17316 22732
rect 17368 22720 17374 22772
rect 17586 22760 17592 22772
rect 17547 22732 17592 22760
rect 17586 22720 17592 22732
rect 17644 22720 17650 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19484 22732 19717 22760
rect 19484 22720 19490 22732
rect 19705 22729 19717 22732
rect 19751 22760 19763 22763
rect 19981 22763 20039 22769
rect 19981 22760 19993 22763
rect 19751 22732 19993 22760
rect 19751 22729 19763 22732
rect 19705 22723 19763 22729
rect 19981 22729 19993 22732
rect 20027 22729 20039 22763
rect 19981 22723 20039 22729
rect 20809 22763 20867 22769
rect 20809 22729 20821 22763
rect 20855 22760 20867 22763
rect 20990 22760 20996 22772
rect 20855 22732 20996 22760
rect 20855 22729 20867 22732
rect 20809 22723 20867 22729
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 23937 22763 23995 22769
rect 23937 22729 23949 22763
rect 23983 22760 23995 22763
rect 25130 22760 25136 22772
rect 23983 22732 25136 22760
rect 23983 22729 23995 22732
rect 23937 22723 23995 22729
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 25682 22760 25688 22772
rect 25643 22732 25688 22760
rect 25682 22720 25688 22732
rect 25740 22720 25746 22772
rect 30742 22760 30748 22772
rect 30655 22732 30748 22760
rect 30742 22720 30748 22732
rect 30800 22760 30806 22772
rect 31202 22760 31208 22772
rect 30800 22732 31208 22760
rect 30800 22720 30806 22732
rect 31202 22720 31208 22732
rect 31260 22720 31266 22772
rect 31757 22763 31815 22769
rect 31757 22729 31769 22763
rect 31803 22760 31815 22763
rect 31938 22760 31944 22772
rect 31803 22732 31944 22760
rect 31803 22729 31815 22732
rect 31757 22723 31815 22729
rect 12713 22695 12771 22701
rect 12713 22661 12725 22695
rect 12759 22692 12771 22695
rect 15473 22695 15531 22701
rect 15473 22692 15485 22695
rect 12759 22664 15485 22692
rect 12759 22661 12771 22664
rect 12713 22655 12771 22661
rect 12820 22565 12848 22664
rect 15473 22661 15485 22664
rect 15519 22661 15531 22695
rect 15473 22655 15531 22661
rect 13262 22584 13268 22636
rect 13320 22624 13326 22636
rect 13449 22627 13507 22633
rect 13449 22624 13461 22627
rect 13320 22596 13461 22624
rect 13320 22584 13326 22596
rect 13449 22593 13461 22596
rect 13495 22624 13507 22627
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 13495 22596 13829 22624
rect 13495 22593 13507 22596
rect 13449 22587 13507 22593
rect 13817 22593 13829 22596
rect 13863 22624 13875 22627
rect 14366 22624 14372 22636
rect 13863 22596 14372 22624
rect 13863 22593 13875 22596
rect 13817 22587 13875 22593
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22624 14611 22627
rect 14642 22624 14648 22636
rect 14599 22596 14648 22624
rect 14599 22593 14611 22596
rect 14553 22587 14611 22593
rect 14642 22584 14648 22596
rect 14700 22624 14706 22636
rect 15102 22624 15108 22636
rect 14700 22596 15108 22624
rect 14700 22584 14706 22596
rect 15102 22584 15108 22596
rect 15160 22584 15166 22636
rect 16022 22624 16028 22636
rect 15983 22596 16028 22624
rect 16022 22584 16028 22596
rect 16080 22584 16086 22636
rect 21545 22627 21603 22633
rect 21545 22593 21557 22627
rect 21591 22624 21603 22627
rect 22649 22627 22707 22633
rect 22649 22624 22661 22627
rect 21591 22596 22661 22624
rect 21591 22593 21603 22596
rect 21545 22587 21603 22593
rect 22649 22593 22661 22596
rect 22695 22624 22707 22627
rect 23382 22624 23388 22636
rect 22695 22596 23388 22624
rect 22695 22593 22707 22596
rect 22649 22587 22707 22593
rect 23382 22584 23388 22596
rect 23440 22584 23446 22636
rect 29917 22627 29975 22633
rect 29917 22593 29929 22627
rect 29963 22624 29975 22627
rect 30098 22624 30104 22636
rect 29963 22596 30104 22624
rect 29963 22593 29975 22596
rect 29917 22587 29975 22593
rect 30098 22584 30104 22596
rect 30156 22624 30162 22636
rect 30285 22627 30343 22633
rect 30285 22624 30297 22627
rect 30156 22596 30297 22624
rect 30156 22584 30162 22596
rect 30285 22593 30297 22596
rect 30331 22593 30343 22627
rect 30285 22587 30343 22593
rect 12805 22559 12863 22565
rect 12805 22525 12817 22559
rect 12851 22525 12863 22559
rect 12805 22519 12863 22525
rect 18325 22559 18383 22565
rect 18325 22525 18337 22559
rect 18371 22525 18383 22559
rect 18325 22519 18383 22525
rect 15838 22488 15844 22500
rect 15751 22460 15844 22488
rect 15838 22448 15844 22460
rect 15896 22488 15902 22500
rect 16853 22491 16911 22497
rect 16853 22488 16865 22491
rect 15896 22460 16865 22488
rect 15896 22448 15902 22460
rect 16853 22457 16865 22460
rect 16899 22457 16911 22491
rect 16853 22451 16911 22457
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 14274 22420 14280 22432
rect 13872 22392 14280 22420
rect 13872 22380 13878 22392
rect 14274 22380 14280 22392
rect 14332 22420 14338 22432
rect 14921 22423 14979 22429
rect 14921 22420 14933 22423
rect 14332 22392 14933 22420
rect 14332 22380 14338 22392
rect 14921 22389 14933 22392
rect 14967 22389 14979 22423
rect 14921 22383 14979 22389
rect 15933 22423 15991 22429
rect 15933 22389 15945 22423
rect 15979 22420 15991 22423
rect 16298 22420 16304 22432
rect 15979 22392 16304 22420
rect 15979 22389 15991 22392
rect 15933 22383 15991 22389
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 18046 22380 18052 22432
rect 18104 22420 18110 22432
rect 18340 22420 18368 22519
rect 18414 22516 18420 22568
rect 18472 22556 18478 22568
rect 18581 22559 18639 22565
rect 18581 22556 18593 22559
rect 18472 22528 18593 22556
rect 18472 22516 18478 22528
rect 18581 22525 18593 22528
rect 18627 22525 18639 22559
rect 18581 22519 18639 22525
rect 22094 22516 22100 22568
rect 22152 22556 22158 22568
rect 22373 22559 22431 22565
rect 22373 22556 22385 22559
rect 22152 22528 22385 22556
rect 22152 22516 22158 22528
rect 22373 22525 22385 22528
rect 22419 22525 22431 22559
rect 26878 22556 26884 22568
rect 26839 22528 26884 22556
rect 22373 22519 22431 22525
rect 26878 22516 26884 22528
rect 26936 22556 26942 22568
rect 27433 22559 27491 22565
rect 27433 22556 27445 22559
rect 26936 22528 27445 22556
rect 26936 22516 26942 22528
rect 27433 22525 27445 22528
rect 27479 22525 27491 22559
rect 27433 22519 27491 22525
rect 28721 22559 28779 22565
rect 28721 22525 28733 22559
rect 28767 22556 28779 22559
rect 29178 22556 29184 22568
rect 28767 22528 29184 22556
rect 28767 22525 28779 22528
rect 28721 22519 28779 22525
rect 29178 22516 29184 22528
rect 29236 22516 29242 22568
rect 31389 22559 31447 22565
rect 31389 22525 31401 22559
rect 31435 22556 31447 22559
rect 31772 22556 31800 22723
rect 31938 22720 31944 22732
rect 31996 22720 32002 22772
rect 32769 22763 32827 22769
rect 32769 22729 32781 22763
rect 32815 22760 32827 22763
rect 33042 22760 33048 22772
rect 32815 22732 33048 22760
rect 32815 22729 32827 22732
rect 32769 22723 32827 22729
rect 33042 22720 33048 22732
rect 33100 22720 33106 22772
rect 34333 22763 34391 22769
rect 34333 22729 34345 22763
rect 34379 22760 34391 22763
rect 34422 22760 34428 22772
rect 34379 22732 34428 22760
rect 34379 22729 34391 22732
rect 34333 22723 34391 22729
rect 34422 22720 34428 22732
rect 34480 22720 34486 22772
rect 32401 22627 32459 22633
rect 32401 22593 32413 22627
rect 32447 22624 32459 22627
rect 33781 22627 33839 22633
rect 33781 22624 33793 22627
rect 32447 22596 33793 22624
rect 32447 22593 32459 22596
rect 32401 22587 32459 22593
rect 33781 22593 33793 22596
rect 33827 22624 33839 22627
rect 34609 22627 34667 22633
rect 34609 22624 34621 22627
rect 33827 22596 34621 22624
rect 33827 22593 33839 22596
rect 33781 22587 33839 22593
rect 34609 22593 34621 22596
rect 34655 22624 34667 22627
rect 34655 22596 35020 22624
rect 34655 22593 34667 22596
rect 34609 22587 34667 22593
rect 31435 22528 31800 22556
rect 33137 22559 33195 22565
rect 31435 22525 31447 22528
rect 31389 22519 31447 22525
rect 33137 22525 33149 22559
rect 33183 22556 33195 22559
rect 33689 22559 33747 22565
rect 33689 22556 33701 22559
rect 33183 22528 33701 22556
rect 33183 22525 33195 22528
rect 33137 22519 33195 22525
rect 33689 22525 33701 22528
rect 33735 22556 33747 22559
rect 34238 22556 34244 22568
rect 33735 22528 34244 22556
rect 33735 22525 33747 22528
rect 33689 22519 33747 22525
rect 34238 22516 34244 22528
rect 34296 22516 34302 22568
rect 34882 22556 34888 22568
rect 34843 22528 34888 22556
rect 34882 22516 34888 22528
rect 34940 22516 34946 22568
rect 34992 22556 35020 22596
rect 35141 22559 35199 22565
rect 35141 22556 35153 22559
rect 34992 22528 35153 22556
rect 35141 22525 35153 22528
rect 35187 22556 35199 22559
rect 35526 22556 35532 22568
rect 35187 22528 35532 22556
rect 35187 22525 35199 22528
rect 35141 22519 35199 22525
rect 35526 22516 35532 22528
rect 35584 22516 35590 22568
rect 21913 22491 21971 22497
rect 21913 22457 21925 22491
rect 21959 22488 21971 22491
rect 24397 22491 24455 22497
rect 21959 22460 22508 22488
rect 21959 22457 21971 22460
rect 21913 22451 21971 22457
rect 20346 22420 20352 22432
rect 18104 22392 20352 22420
rect 18104 22380 18110 22392
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 22002 22420 22008 22432
rect 21963 22392 22008 22420
rect 22002 22380 22008 22392
rect 22060 22380 22066 22432
rect 22480 22429 22508 22460
rect 24397 22457 24409 22491
rect 24443 22457 24455 22491
rect 24397 22451 24455 22457
rect 29089 22491 29147 22497
rect 29089 22457 29101 22491
rect 29135 22488 29147 22491
rect 29641 22491 29699 22497
rect 29641 22488 29653 22491
rect 29135 22460 29653 22488
rect 29135 22457 29147 22460
rect 29089 22451 29147 22457
rect 29641 22457 29653 22460
rect 29687 22488 29699 22491
rect 30006 22488 30012 22500
rect 29687 22460 30012 22488
rect 29687 22457 29699 22460
rect 29641 22451 29699 22457
rect 22465 22423 22523 22429
rect 22465 22389 22477 22423
rect 22511 22420 22523 22423
rect 22738 22420 22744 22432
rect 22511 22392 22744 22420
rect 22511 22389 22523 22392
rect 22465 22383 22523 22389
rect 22738 22380 22744 22392
rect 22796 22380 22802 22432
rect 23934 22380 23940 22432
rect 23992 22420 23998 22432
rect 24213 22423 24271 22429
rect 24213 22420 24225 22423
rect 23992 22392 24225 22420
rect 23992 22380 23998 22392
rect 24213 22389 24225 22392
rect 24259 22420 24271 22423
rect 24412 22420 24440 22451
rect 30006 22448 30012 22460
rect 30064 22448 30070 22500
rect 33594 22488 33600 22500
rect 33555 22460 33600 22488
rect 33594 22448 33600 22460
rect 33652 22488 33658 22500
rect 34146 22488 34152 22500
rect 33652 22460 34152 22488
rect 33652 22448 33658 22460
rect 34146 22448 34152 22460
rect 34204 22448 34210 22500
rect 34900 22488 34928 22516
rect 36541 22491 36599 22497
rect 36541 22488 36553 22491
rect 34900 22460 36553 22488
rect 36541 22457 36553 22460
rect 36587 22488 36599 22491
rect 36630 22488 36636 22500
rect 36587 22460 36636 22488
rect 36587 22457 36599 22460
rect 36541 22451 36599 22457
rect 36630 22448 36636 22460
rect 36688 22448 36694 22500
rect 24259 22392 24440 22420
rect 24259 22389 24271 22392
rect 24213 22383 24271 22389
rect 25222 22380 25228 22432
rect 25280 22420 25286 22432
rect 27065 22423 27123 22429
rect 27065 22420 27077 22423
rect 25280 22392 27077 22420
rect 25280 22380 25286 22392
rect 27065 22389 27077 22392
rect 27111 22389 27123 22423
rect 27065 22383 27123 22389
rect 27798 22380 27804 22432
rect 27856 22420 27862 22432
rect 28077 22423 28135 22429
rect 28077 22420 28089 22423
rect 27856 22392 28089 22420
rect 27856 22380 27862 22392
rect 28077 22389 28089 22392
rect 28123 22389 28135 22423
rect 29270 22420 29276 22432
rect 29231 22392 29276 22420
rect 28077 22383 28135 22389
rect 29270 22380 29276 22392
rect 29328 22380 29334 22432
rect 29730 22380 29736 22432
rect 29788 22420 29794 22432
rect 29788 22392 29833 22420
rect 29788 22380 29794 22392
rect 33134 22380 33140 22432
rect 33192 22420 33198 22432
rect 33229 22423 33287 22429
rect 33229 22420 33241 22423
rect 33192 22392 33241 22420
rect 33192 22380 33198 22392
rect 33229 22389 33241 22392
rect 33275 22389 33287 22423
rect 36262 22420 36268 22432
rect 36223 22392 36268 22420
rect 33229 22383 33287 22389
rect 36262 22380 36268 22392
rect 36320 22380 36326 22432
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 12618 22216 12624 22228
rect 12579 22188 12624 22216
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 14642 22216 14648 22228
rect 14603 22188 14648 22216
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 15010 22216 15016 22228
rect 14971 22188 15016 22216
rect 15010 22176 15016 22188
rect 15068 22176 15074 22228
rect 15289 22219 15347 22225
rect 15289 22185 15301 22219
rect 15335 22216 15347 22219
rect 15654 22216 15660 22228
rect 15335 22188 15660 22216
rect 15335 22185 15347 22188
rect 15289 22179 15347 22185
rect 15654 22176 15660 22188
rect 15712 22176 15718 22228
rect 16853 22219 16911 22225
rect 16853 22185 16865 22219
rect 16899 22216 16911 22219
rect 17310 22216 17316 22228
rect 16899 22188 17316 22216
rect 16899 22185 16911 22188
rect 16853 22179 16911 22185
rect 17310 22176 17316 22188
rect 17368 22176 17374 22228
rect 17586 22176 17592 22228
rect 17644 22216 17650 22228
rect 18417 22219 18475 22225
rect 18417 22216 18429 22219
rect 17644 22188 18429 22216
rect 17644 22176 17650 22188
rect 18417 22185 18429 22188
rect 18463 22185 18475 22219
rect 18417 22179 18475 22185
rect 18506 22176 18512 22228
rect 18564 22216 18570 22228
rect 18785 22219 18843 22225
rect 18785 22216 18797 22219
rect 18564 22188 18797 22216
rect 18564 22176 18570 22188
rect 18785 22185 18797 22188
rect 18831 22216 18843 22219
rect 19334 22216 19340 22228
rect 18831 22188 19340 22216
rect 18831 22185 18843 22188
rect 18785 22179 18843 22185
rect 19334 22176 19340 22188
rect 19392 22176 19398 22228
rect 19889 22219 19947 22225
rect 19889 22185 19901 22219
rect 19935 22216 19947 22219
rect 20346 22216 20352 22228
rect 19935 22188 20352 22216
rect 19935 22185 19947 22188
rect 19889 22179 19947 22185
rect 20346 22176 20352 22188
rect 20404 22176 20410 22228
rect 24857 22219 24915 22225
rect 24857 22185 24869 22219
rect 24903 22216 24915 22219
rect 25130 22216 25136 22228
rect 24903 22188 25136 22216
rect 24903 22185 24915 22188
rect 24857 22179 24915 22185
rect 25130 22176 25136 22188
rect 25188 22176 25194 22228
rect 29089 22219 29147 22225
rect 29089 22185 29101 22219
rect 29135 22216 29147 22219
rect 29270 22216 29276 22228
rect 29135 22188 29276 22216
rect 29135 22185 29147 22188
rect 29089 22179 29147 22185
rect 15120 22120 15700 22148
rect 11790 22040 11796 22092
rect 11848 22080 11854 22092
rect 12802 22080 12808 22092
rect 11848 22052 12572 22080
rect 12763 22052 12808 22080
rect 11848 22040 11854 22052
rect 12544 22012 12572 22052
rect 12802 22040 12808 22052
rect 12860 22040 12866 22092
rect 12986 22040 12992 22092
rect 13044 22080 13050 22092
rect 13164 22083 13222 22089
rect 13164 22080 13176 22083
rect 13044 22052 13176 22080
rect 13044 22040 13050 22052
rect 13164 22049 13176 22052
rect 13210 22080 13222 22083
rect 13722 22080 13728 22092
rect 13210 22052 13728 22080
rect 13210 22049 13222 22052
rect 13164 22043 13222 22049
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 14734 22040 14740 22092
rect 14792 22080 14798 22092
rect 15120 22080 15148 22120
rect 15672 22089 15700 22120
rect 22094 22108 22100 22160
rect 22152 22148 22158 22160
rect 27614 22148 27620 22160
rect 22152 22120 23428 22148
rect 27575 22120 27620 22148
rect 22152 22108 22158 22120
rect 14792 22052 15148 22080
rect 15657 22083 15715 22089
rect 14792 22040 14798 22052
rect 15657 22049 15669 22083
rect 15703 22080 15715 22083
rect 15930 22080 15936 22092
rect 15703 22052 15737 22080
rect 15843 22052 15936 22080
rect 15703 22049 15715 22052
rect 15657 22043 15715 22049
rect 12897 22015 12955 22021
rect 12897 22012 12909 22015
rect 12544 21984 12909 22012
rect 12544 21885 12572 21984
rect 12897 21981 12909 21984
rect 12943 21981 12955 22015
rect 15102 22012 15108 22024
rect 12897 21975 12955 21981
rect 14292 21984 15108 22012
rect 14292 21956 14320 21984
rect 15102 21972 15108 21984
rect 15160 22012 15166 22024
rect 15856 22021 15884 22052
rect 15930 22040 15936 22052
rect 15988 22080 15994 22092
rect 17221 22083 17279 22089
rect 15988 22052 16804 22080
rect 15988 22040 15994 22052
rect 15749 22015 15807 22021
rect 15749 22012 15761 22015
rect 15160 21984 15761 22012
rect 15160 21972 15166 21984
rect 15749 21981 15761 21984
rect 15795 21981 15807 22015
rect 15749 21975 15807 21981
rect 15841 22015 15899 22021
rect 15841 21981 15853 22015
rect 15887 21981 15899 22015
rect 15841 21975 15899 21981
rect 14274 21944 14280 21956
rect 14187 21916 14280 21944
rect 14274 21904 14280 21916
rect 14332 21904 14338 21956
rect 14642 21904 14648 21956
rect 14700 21944 14706 21956
rect 15856 21944 15884 21975
rect 16776 21953 16804 22052
rect 17221 22049 17233 22083
rect 17267 22080 17279 22083
rect 17678 22080 17684 22092
rect 17267 22052 17684 22080
rect 17267 22049 17279 22052
rect 17221 22043 17279 22049
rect 17678 22040 17684 22052
rect 17736 22040 17742 22092
rect 20990 22040 20996 22092
rect 21048 22080 21054 22092
rect 21157 22083 21215 22089
rect 21157 22080 21169 22083
rect 21048 22052 21169 22080
rect 21048 22040 21054 22052
rect 21157 22049 21169 22052
rect 21203 22049 21215 22083
rect 23400 22080 23428 22120
rect 27614 22108 27620 22120
rect 27672 22108 27678 22160
rect 29104 22148 29132 22179
rect 29270 22176 29276 22188
rect 29328 22176 29334 22228
rect 33229 22219 33287 22225
rect 33229 22185 33241 22219
rect 33275 22216 33287 22219
rect 33962 22216 33968 22228
rect 33275 22188 33968 22216
rect 33275 22185 33287 22188
rect 33229 22179 33287 22185
rect 33962 22176 33968 22188
rect 34020 22176 34026 22228
rect 34054 22176 34060 22228
rect 34112 22216 34118 22228
rect 34241 22219 34299 22225
rect 34241 22216 34253 22219
rect 34112 22188 34253 22216
rect 34112 22176 34118 22188
rect 34241 22185 34253 22188
rect 34287 22216 34299 22219
rect 34517 22219 34575 22225
rect 34517 22216 34529 22219
rect 34287 22188 34529 22216
rect 34287 22185 34299 22188
rect 34241 22179 34299 22185
rect 34517 22185 34529 22188
rect 34563 22216 34575 22219
rect 34609 22219 34667 22225
rect 34609 22216 34621 22219
rect 34563 22188 34621 22216
rect 34563 22185 34575 22188
rect 34517 22179 34575 22185
rect 34609 22185 34621 22188
rect 34655 22216 34667 22219
rect 34882 22216 34888 22228
rect 34655 22188 34888 22216
rect 34655 22185 34667 22188
rect 34609 22179 34667 22185
rect 34882 22176 34888 22188
rect 34940 22176 34946 22228
rect 30193 22151 30251 22157
rect 30193 22148 30205 22151
rect 28920 22120 29132 22148
rect 29196 22120 30205 22148
rect 23750 22089 23756 22092
rect 23733 22083 23756 22089
rect 23733 22080 23745 22083
rect 23400 22052 23745 22080
rect 21157 22043 21215 22049
rect 23733 22049 23745 22052
rect 23808 22080 23814 22092
rect 23808 22052 23881 22080
rect 23733 22043 23756 22049
rect 23750 22040 23756 22043
rect 23808 22040 23814 22052
rect 26234 22040 26240 22092
rect 26292 22080 26298 22092
rect 26510 22080 26516 22092
rect 26292 22052 26516 22080
rect 26292 22040 26298 22052
rect 26510 22040 26516 22052
rect 26568 22040 26574 22092
rect 28537 22083 28595 22089
rect 28537 22049 28549 22083
rect 28583 22080 28595 22083
rect 28920 22080 28948 22120
rect 28583 22052 28948 22080
rect 28997 22083 29055 22089
rect 28583 22049 28595 22052
rect 28537 22043 28595 22049
rect 28997 22049 29009 22083
rect 29043 22080 29055 22083
rect 29196 22080 29224 22120
rect 30193 22117 30205 22120
rect 30239 22117 30251 22151
rect 36262 22148 36268 22160
rect 30193 22111 30251 22117
rect 35912 22120 36268 22148
rect 29043 22052 29224 22080
rect 29043 22049 29055 22052
rect 28997 22043 29055 22049
rect 17310 22012 17316 22024
rect 17271 21984 17316 22012
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17497 22015 17555 22021
rect 17497 21981 17509 22015
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 18141 22015 18199 22021
rect 18141 21981 18153 22015
rect 18187 22012 18199 22015
rect 18874 22012 18880 22024
rect 18187 21984 18880 22012
rect 18187 21981 18199 21984
rect 18141 21975 18199 21981
rect 14700 21916 15884 21944
rect 16761 21947 16819 21953
rect 14700 21904 14706 21916
rect 16761 21913 16773 21947
rect 16807 21944 16819 21947
rect 17512 21944 17540 21975
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 19061 22015 19119 22021
rect 19061 21981 19073 22015
rect 19107 22012 19119 22015
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 19107 21984 19441 22012
rect 19107 21981 19119 21984
rect 19061 21975 19119 21981
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 21981 20959 22015
rect 20901 21975 20959 21981
rect 23477 22015 23535 22021
rect 23477 21981 23489 22015
rect 23523 21981 23535 22015
rect 23477 21975 23535 21981
rect 19076 21944 19104 21975
rect 16807 21916 19104 21944
rect 16807 21913 16819 21916
rect 16761 21907 16819 21913
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 12894 21876 12900 21888
rect 12575 21848 12900 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 16298 21876 16304 21888
rect 16259 21848 16304 21876
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 20916 21876 20944 21975
rect 21266 21876 21272 21888
rect 20916 21848 21272 21876
rect 21266 21836 21272 21848
rect 21324 21836 21330 21888
rect 21634 21836 21640 21888
rect 21692 21876 21698 21888
rect 22281 21879 22339 21885
rect 22281 21876 22293 21879
rect 21692 21848 22293 21876
rect 21692 21836 21698 21848
rect 22281 21845 22293 21848
rect 22327 21845 22339 21879
rect 22281 21839 22339 21845
rect 23106 21836 23112 21888
rect 23164 21876 23170 21888
rect 23492 21876 23520 21975
rect 28810 21972 28816 22024
rect 28868 22012 28874 22024
rect 29012 22012 29040 22043
rect 29454 22040 29460 22092
rect 29512 22080 29518 22092
rect 29730 22080 29736 22092
rect 29512 22052 29736 22080
rect 29512 22040 29518 22052
rect 29730 22040 29736 22052
rect 29788 22040 29794 22092
rect 33594 22080 33600 22092
rect 33555 22052 33600 22080
rect 33594 22040 33600 22052
rect 33652 22040 33658 22092
rect 34698 22080 34704 22092
rect 33888 22052 34704 22080
rect 29178 22012 29184 22024
rect 28868 21984 29040 22012
rect 29139 21984 29184 22012
rect 28868 21972 28874 21984
rect 29178 21972 29184 21984
rect 29236 21972 29242 22024
rect 32950 21972 32956 22024
rect 33008 22012 33014 22024
rect 33134 22012 33140 22024
rect 33008 21984 33140 22012
rect 33008 21972 33014 21984
rect 33134 21972 33140 21984
rect 33192 22012 33198 22024
rect 33888 22021 33916 22052
rect 34698 22040 34704 22052
rect 34756 22080 34762 22092
rect 35060 22083 35118 22089
rect 35060 22080 35072 22083
rect 34756 22052 35072 22080
rect 34756 22040 34762 22052
rect 35060 22049 35072 22052
rect 35106 22080 35118 22083
rect 35912 22080 35940 22120
rect 36262 22108 36268 22120
rect 36320 22108 36326 22160
rect 35106 22052 35940 22080
rect 35106 22049 35118 22052
rect 35060 22043 35118 22049
rect 33689 22015 33747 22021
rect 33689 22012 33701 22015
rect 33192 21984 33701 22012
rect 33192 21972 33198 21984
rect 33689 21981 33701 21984
rect 33735 21981 33747 22015
rect 33689 21975 33747 21981
rect 33873 22015 33931 22021
rect 33873 21981 33885 22015
rect 33919 21981 33931 22015
rect 33873 21975 33931 21981
rect 34517 22015 34575 22021
rect 34517 21981 34529 22015
rect 34563 22012 34575 22015
rect 34790 22012 34796 22024
rect 34563 21984 34796 22012
rect 34563 21981 34575 21984
rect 34517 21975 34575 21981
rect 34790 21972 34796 21984
rect 34848 21972 34854 22024
rect 24670 21876 24676 21888
rect 23164 21848 24676 21876
rect 23164 21836 23170 21848
rect 24670 21836 24676 21848
rect 24728 21876 24734 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 24728 21848 25237 21876
rect 24728 21836 24734 21848
rect 25225 21845 25237 21848
rect 25271 21876 25283 21879
rect 25498 21876 25504 21888
rect 25271 21848 25504 21876
rect 25271 21845 25283 21848
rect 25225 21839 25283 21845
rect 25498 21836 25504 21848
rect 25556 21876 25562 21888
rect 25593 21879 25651 21885
rect 25593 21876 25605 21879
rect 25556 21848 25605 21876
rect 25556 21836 25562 21848
rect 25593 21845 25605 21848
rect 25639 21845 25651 21879
rect 26694 21876 26700 21888
rect 26655 21848 26700 21876
rect 25593 21839 25651 21845
rect 26694 21836 26700 21848
rect 26752 21836 26758 21888
rect 28626 21876 28632 21888
rect 28587 21848 28632 21876
rect 28626 21836 28632 21848
rect 28684 21836 28690 21888
rect 30098 21876 30104 21888
rect 30059 21848 30104 21876
rect 30098 21836 30104 21848
rect 30156 21836 30162 21888
rect 31202 21836 31208 21888
rect 31260 21876 31266 21888
rect 31481 21879 31539 21885
rect 31481 21876 31493 21879
rect 31260 21848 31493 21876
rect 31260 21836 31266 21848
rect 31481 21845 31493 21848
rect 31527 21845 31539 21879
rect 33134 21876 33140 21888
rect 33095 21848 33140 21876
rect 31481 21839 31539 21845
rect 33134 21836 33140 21848
rect 33192 21836 33198 21888
rect 35710 21836 35716 21888
rect 35768 21876 35774 21888
rect 36173 21879 36231 21885
rect 36173 21876 36185 21879
rect 35768 21848 36185 21876
rect 35768 21836 35774 21848
rect 36173 21845 36185 21848
rect 36219 21845 36231 21879
rect 36173 21839 36231 21845
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 11790 21672 11796 21684
rect 11751 21644 11796 21672
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12897 21675 12955 21681
rect 12897 21641 12909 21675
rect 12943 21672 12955 21675
rect 12986 21672 12992 21684
rect 12943 21644 12992 21672
rect 12943 21641 12955 21644
rect 12897 21635 12955 21641
rect 12986 21632 12992 21644
rect 13044 21632 13050 21684
rect 14369 21675 14427 21681
rect 14369 21641 14381 21675
rect 14415 21672 14427 21675
rect 14734 21672 14740 21684
rect 14415 21644 14740 21672
rect 14415 21641 14427 21644
rect 14369 21635 14427 21641
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 15102 21672 15108 21684
rect 15063 21644 15108 21672
rect 15102 21632 15108 21644
rect 15160 21632 15166 21684
rect 15197 21675 15255 21681
rect 15197 21641 15209 21675
rect 15243 21672 15255 21675
rect 16298 21672 16304 21684
rect 15243 21644 16304 21672
rect 15243 21641 15255 21644
rect 15197 21635 15255 21641
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 16666 21672 16672 21684
rect 16627 21644 16672 21672
rect 16666 21632 16672 21644
rect 16724 21632 16730 21684
rect 16942 21672 16948 21684
rect 16903 21644 16948 21672
rect 16942 21632 16948 21644
rect 17000 21632 17006 21684
rect 17678 21672 17684 21684
rect 17639 21644 17684 21672
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 19429 21675 19487 21681
rect 19429 21672 19441 21675
rect 19392 21644 19441 21672
rect 19392 21632 19398 21644
rect 19429 21641 19441 21644
rect 19475 21672 19487 21675
rect 20073 21675 20131 21681
rect 20073 21672 20085 21675
rect 19475 21644 20085 21672
rect 19475 21641 19487 21644
rect 19429 21635 19487 21641
rect 20073 21641 20085 21644
rect 20119 21641 20131 21675
rect 22738 21672 22744 21684
rect 22699 21644 22744 21672
rect 20073 21635 20131 21641
rect 22738 21632 22744 21644
rect 22796 21632 22802 21684
rect 23106 21672 23112 21684
rect 23067 21644 23112 21672
rect 23106 21632 23112 21644
rect 23164 21632 23170 21684
rect 23750 21632 23756 21684
rect 23808 21672 23814 21684
rect 23845 21675 23903 21681
rect 23845 21672 23857 21675
rect 23808 21644 23857 21672
rect 23808 21632 23814 21644
rect 23845 21641 23857 21644
rect 23891 21641 23903 21675
rect 23845 21635 23903 21641
rect 24029 21675 24087 21681
rect 24029 21641 24041 21675
rect 24075 21672 24087 21675
rect 24762 21672 24768 21684
rect 24075 21644 24768 21672
rect 24075 21641 24087 21644
rect 24029 21635 24087 21641
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 26510 21632 26516 21684
rect 26568 21672 26574 21684
rect 27249 21675 27307 21681
rect 27249 21672 27261 21675
rect 26568 21644 27261 21672
rect 26568 21632 26574 21644
rect 27249 21641 27261 21644
rect 27295 21641 27307 21675
rect 28442 21672 28448 21684
rect 28403 21644 28448 21672
rect 27249 21635 27307 21641
rect 28442 21632 28448 21644
rect 28500 21632 28506 21684
rect 28810 21672 28816 21684
rect 28771 21644 28816 21672
rect 28810 21632 28816 21644
rect 28868 21632 28874 21684
rect 29178 21632 29184 21684
rect 29236 21672 29242 21684
rect 30653 21675 30711 21681
rect 30653 21672 30665 21675
rect 29236 21644 30665 21672
rect 29236 21632 29242 21644
rect 30653 21641 30665 21644
rect 30699 21641 30711 21675
rect 30653 21635 30711 21641
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21672 32827 21675
rect 33226 21672 33232 21684
rect 32815 21644 33232 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 33226 21632 33232 21644
rect 33284 21632 33290 21684
rect 34333 21675 34391 21681
rect 34333 21641 34345 21675
rect 34379 21672 34391 21675
rect 34698 21672 34704 21684
rect 34379 21644 34704 21672
rect 34379 21641 34391 21644
rect 34333 21635 34391 21641
rect 34698 21632 34704 21644
rect 34756 21632 34762 21684
rect 36630 21672 36636 21684
rect 36591 21644 36636 21672
rect 36630 21632 36636 21644
rect 36688 21632 36694 21684
rect 31481 21607 31539 21613
rect 31481 21573 31493 21607
rect 31527 21604 31539 21607
rect 34514 21604 34520 21616
rect 31527 21576 34520 21604
rect 31527 21573 31539 21576
rect 31481 21567 31539 21573
rect 34514 21564 34520 21576
rect 34572 21564 34578 21616
rect 12253 21539 12311 21545
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 15841 21539 15899 21545
rect 12299 21508 13124 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 12986 21468 12992 21480
rect 12947 21440 12992 21468
rect 12986 21428 12992 21440
rect 13044 21428 13050 21480
rect 13096 21468 13124 21508
rect 15841 21505 15853 21539
rect 15887 21536 15899 21539
rect 15930 21536 15936 21548
rect 15887 21508 15936 21536
rect 15887 21505 15899 21508
rect 15841 21499 15899 21505
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 24486 21536 24492 21548
rect 24447 21508 24492 21536
rect 24486 21496 24492 21508
rect 24544 21496 24550 21548
rect 24670 21536 24676 21548
rect 24631 21508 24676 21536
rect 24670 21496 24676 21508
rect 24728 21496 24734 21548
rect 31570 21496 31576 21548
rect 31628 21536 31634 21548
rect 32033 21539 32091 21545
rect 32033 21536 32045 21539
rect 31628 21508 32045 21536
rect 31628 21496 31634 21508
rect 32033 21505 32045 21508
rect 32079 21505 32091 21539
rect 32033 21499 32091 21505
rect 33134 21496 33140 21548
rect 33192 21536 33198 21548
rect 33781 21539 33839 21545
rect 33781 21536 33793 21539
rect 33192 21508 33793 21536
rect 33192 21496 33198 21508
rect 33781 21505 33793 21508
rect 33827 21536 33839 21539
rect 33827 21508 35112 21536
rect 33827 21505 33839 21508
rect 33781 21499 33839 21505
rect 13256 21471 13314 21477
rect 13256 21468 13268 21471
rect 13096 21440 13268 21468
rect 13256 21437 13268 21440
rect 13302 21468 13314 21471
rect 14274 21468 14280 21480
rect 13302 21440 14280 21468
rect 13302 21437 13314 21440
rect 13256 21431 13314 21437
rect 14274 21428 14280 21440
rect 14332 21428 14338 21480
rect 16666 21428 16672 21480
rect 16724 21468 16730 21480
rect 16761 21471 16819 21477
rect 16761 21468 16773 21471
rect 16724 21440 16773 21468
rect 16724 21428 16730 21440
rect 16761 21437 16773 21440
rect 16807 21437 16819 21471
rect 18046 21468 18052 21480
rect 18007 21440 18052 21468
rect 16761 21431 16819 21437
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 21358 21468 21364 21480
rect 21319 21440 21364 21468
rect 21358 21428 21364 21440
rect 21416 21428 21422 21480
rect 21634 21477 21640 21480
rect 21628 21468 21640 21477
rect 21468 21440 21640 21468
rect 15286 21360 15292 21412
rect 15344 21400 15350 21412
rect 15565 21403 15623 21409
rect 15565 21400 15577 21403
rect 15344 21372 15577 21400
rect 15344 21360 15350 21372
rect 15565 21369 15577 21372
rect 15611 21400 15623 21403
rect 16209 21403 16267 21409
rect 16209 21400 16221 21403
rect 15611 21372 16221 21400
rect 15611 21369 15623 21372
rect 15565 21363 15623 21369
rect 16209 21369 16221 21372
rect 16255 21369 16267 21403
rect 16209 21363 16267 21369
rect 18316 21403 18374 21409
rect 18316 21369 18328 21403
rect 18362 21400 18374 21403
rect 18874 21400 18880 21412
rect 18362 21372 18880 21400
rect 18362 21369 18374 21372
rect 18316 21363 18374 21369
rect 18874 21360 18880 21372
rect 18932 21400 18938 21412
rect 18932 21372 19472 21400
rect 18932 21360 18938 21372
rect 19444 21344 19472 21372
rect 19886 21360 19892 21412
rect 19944 21400 19950 21412
rect 20625 21403 20683 21409
rect 20625 21400 20637 21403
rect 19944 21372 20637 21400
rect 19944 21360 19950 21372
rect 20625 21369 20637 21372
rect 20671 21400 20683 21403
rect 21468 21400 21496 21440
rect 21628 21431 21640 21440
rect 21634 21428 21640 21431
rect 21692 21428 21698 21480
rect 25498 21428 25504 21480
rect 25556 21468 25562 21480
rect 25593 21471 25651 21477
rect 25593 21468 25605 21471
rect 25556 21440 25605 21468
rect 25556 21428 25562 21440
rect 25593 21437 25605 21440
rect 25639 21468 25651 21471
rect 26786 21468 26792 21480
rect 25639 21440 26792 21468
rect 25639 21437 25651 21440
rect 25593 21431 25651 21437
rect 26786 21428 26792 21440
rect 26844 21428 26850 21480
rect 27801 21471 27859 21477
rect 27801 21437 27813 21471
rect 27847 21468 27859 21471
rect 28442 21468 28448 21480
rect 27847 21440 28448 21468
rect 27847 21437 27859 21440
rect 27801 21431 27859 21437
rect 28442 21428 28448 21440
rect 28500 21428 28506 21480
rect 28902 21428 28908 21480
rect 28960 21468 28966 21480
rect 29273 21471 29331 21477
rect 29273 21468 29285 21471
rect 28960 21440 29285 21468
rect 28960 21428 28966 21440
rect 29273 21437 29285 21440
rect 29319 21437 29331 21471
rect 29273 21431 29331 21437
rect 29540 21471 29598 21477
rect 29540 21437 29552 21471
rect 29586 21468 29598 21471
rect 30098 21468 30104 21480
rect 29586 21440 30104 21468
rect 29586 21437 29598 21440
rect 29540 21431 29598 21437
rect 25866 21409 25872 21412
rect 25838 21403 25872 21409
rect 25838 21400 25850 21403
rect 20671 21372 21496 21400
rect 25424 21372 25850 21400
rect 20671 21369 20683 21372
rect 20625 21363 20683 21369
rect 15654 21332 15660 21344
rect 15615 21304 15660 21332
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 17310 21332 17316 21344
rect 17271 21304 17316 21332
rect 17310 21292 17316 21304
rect 17368 21292 17374 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19705 21335 19763 21341
rect 19705 21332 19717 21335
rect 19484 21304 19717 21332
rect 19484 21292 19490 21304
rect 19705 21301 19717 21304
rect 19751 21301 19763 21335
rect 20898 21332 20904 21344
rect 20859 21304 20904 21332
rect 19705 21295 19763 21301
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 23842 21332 23848 21344
rect 23523 21304 23848 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 23842 21292 23848 21304
rect 23900 21332 23906 21344
rect 24397 21335 24455 21341
rect 24397 21332 24409 21335
rect 23900 21304 24409 21332
rect 23900 21292 23906 21304
rect 24397 21301 24409 21304
rect 24443 21301 24455 21335
rect 24397 21295 24455 21301
rect 25130 21292 25136 21344
rect 25188 21332 25194 21344
rect 25424 21341 25452 21372
rect 25838 21369 25850 21372
rect 25924 21400 25930 21412
rect 27709 21403 27767 21409
rect 25924 21372 25986 21400
rect 25838 21363 25872 21369
rect 25866 21360 25872 21363
rect 25924 21360 25930 21372
rect 27709 21369 27721 21403
rect 27755 21400 27767 21403
rect 28920 21400 28948 21428
rect 27755 21372 28948 21400
rect 29288 21400 29316 21431
rect 30098 21428 30104 21440
rect 30156 21428 30162 21480
rect 31389 21471 31447 21477
rect 31389 21437 31401 21471
rect 31435 21468 31447 21471
rect 31846 21468 31852 21480
rect 31435 21440 31852 21468
rect 31435 21437 31447 21440
rect 31389 21431 31447 21437
rect 31846 21428 31852 21440
rect 31904 21428 31910 21480
rect 33226 21428 33232 21480
rect 33284 21468 33290 21480
rect 33597 21471 33655 21477
rect 33597 21468 33609 21471
rect 33284 21440 33609 21468
rect 33284 21428 33290 21440
rect 33597 21437 33609 21440
rect 33643 21468 33655 21471
rect 33962 21468 33968 21480
rect 33643 21440 33968 21468
rect 33643 21437 33655 21440
rect 33597 21431 33655 21437
rect 33962 21428 33968 21440
rect 34020 21428 34026 21480
rect 34054 21428 34060 21480
rect 34112 21428 34118 21480
rect 34514 21428 34520 21480
rect 34572 21468 34578 21480
rect 34698 21468 34704 21480
rect 34572 21440 34704 21468
rect 34572 21428 34578 21440
rect 34698 21428 34704 21440
rect 34756 21428 34762 21480
rect 34790 21428 34796 21480
rect 34848 21468 34854 21480
rect 34977 21471 35035 21477
rect 34977 21468 34989 21471
rect 34848 21440 34989 21468
rect 34848 21428 34854 21440
rect 34977 21437 34989 21440
rect 35023 21437 35035 21471
rect 35084 21468 35112 21508
rect 35233 21471 35291 21477
rect 35233 21468 35245 21471
rect 35084 21440 35245 21468
rect 34977 21431 35035 21437
rect 35233 21437 35245 21440
rect 35279 21468 35291 21471
rect 35618 21468 35624 21480
rect 35279 21440 35624 21468
rect 35279 21437 35291 21440
rect 35233 21431 35291 21437
rect 29822 21400 29828 21412
rect 29288 21372 29828 21400
rect 27755 21369 27767 21372
rect 27709 21363 27767 21369
rect 29822 21360 29828 21372
rect 29880 21400 29886 21412
rect 30742 21400 30748 21412
rect 29880 21372 30748 21400
rect 29880 21360 29886 21372
rect 30742 21360 30748 21372
rect 30800 21400 30806 21412
rect 31021 21403 31079 21409
rect 31021 21400 31033 21403
rect 30800 21372 31033 21400
rect 30800 21360 30806 21372
rect 31021 21369 31033 21372
rect 31067 21400 31079 21403
rect 31662 21400 31668 21412
rect 31067 21372 31668 21400
rect 31067 21369 31079 21372
rect 31021 21363 31079 21369
rect 31662 21360 31668 21372
rect 31720 21360 31726 21412
rect 33137 21403 33195 21409
rect 33137 21369 33149 21403
rect 33183 21400 33195 21403
rect 34072 21400 34100 21428
rect 34606 21400 34612 21412
rect 33183 21372 33732 21400
rect 34072 21372 34612 21400
rect 33183 21369 33195 21372
rect 33137 21363 33195 21369
rect 25409 21335 25467 21341
rect 25409 21332 25421 21335
rect 25188 21304 25421 21332
rect 25188 21292 25194 21304
rect 25409 21301 25421 21304
rect 25455 21301 25467 21335
rect 25409 21295 25467 21301
rect 26973 21335 27031 21341
rect 26973 21301 26985 21335
rect 27019 21332 27031 21335
rect 27062 21332 27068 21344
rect 27019 21304 27068 21332
rect 27019 21301 27031 21304
rect 26973 21295 27031 21301
rect 27062 21292 27068 21304
rect 27120 21292 27126 21344
rect 27982 21332 27988 21344
rect 27943 21304 27988 21332
rect 27982 21292 27988 21304
rect 28040 21292 28046 21344
rect 31202 21292 31208 21344
rect 31260 21332 31266 21344
rect 31941 21335 31999 21341
rect 31941 21332 31953 21335
rect 31260 21304 31953 21332
rect 31260 21292 31266 21304
rect 31941 21301 31953 21304
rect 31987 21301 31999 21335
rect 33226 21332 33232 21344
rect 33187 21304 33232 21332
rect 31941 21295 31999 21301
rect 33226 21292 33232 21304
rect 33284 21292 33290 21344
rect 33704 21341 33732 21372
rect 34606 21360 34612 21372
rect 34664 21360 34670 21412
rect 34992 21400 35020 21431
rect 35618 21428 35624 21440
rect 35676 21428 35682 21480
rect 35434 21400 35440 21412
rect 34992 21372 35440 21400
rect 35434 21360 35440 21372
rect 35492 21360 35498 21412
rect 33689 21335 33747 21341
rect 33689 21301 33701 21335
rect 33735 21332 33747 21335
rect 33870 21332 33876 21344
rect 33735 21304 33876 21332
rect 33735 21301 33747 21304
rect 33689 21295 33747 21301
rect 33870 21292 33876 21304
rect 33928 21332 33934 21344
rect 35158 21332 35164 21344
rect 33928 21304 35164 21332
rect 33928 21292 33934 21304
rect 35158 21292 35164 21304
rect 35216 21292 35222 21344
rect 35894 21292 35900 21344
rect 35952 21332 35958 21344
rect 36357 21335 36415 21341
rect 36357 21332 36369 21335
rect 35952 21304 36369 21332
rect 35952 21292 35958 21304
rect 36357 21301 36369 21304
rect 36403 21301 36415 21335
rect 36357 21295 36415 21301
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 12713 21131 12771 21137
rect 12713 21097 12725 21131
rect 12759 21128 12771 21131
rect 12802 21128 12808 21140
rect 12759 21100 12808 21128
rect 12759 21097 12771 21100
rect 12713 21091 12771 21097
rect 12802 21088 12808 21100
rect 12860 21088 12866 21140
rect 14182 21088 14188 21140
rect 14240 21128 14246 21140
rect 14369 21131 14427 21137
rect 14369 21128 14381 21131
rect 14240 21100 14381 21128
rect 14240 21088 14246 21100
rect 14369 21097 14381 21100
rect 14415 21128 14427 21131
rect 15565 21131 15623 21137
rect 15565 21128 15577 21131
rect 14415 21100 15577 21128
rect 14415 21097 14427 21100
rect 14369 21091 14427 21097
rect 15565 21097 15577 21100
rect 15611 21128 15623 21131
rect 15654 21128 15660 21140
rect 15611 21100 15660 21128
rect 15611 21097 15623 21100
rect 15565 21091 15623 21097
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 15930 21128 15936 21140
rect 15891 21100 15936 21128
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 17589 21131 17647 21137
rect 17589 21097 17601 21131
rect 17635 21128 17647 21131
rect 17678 21128 17684 21140
rect 17635 21100 17684 21128
rect 17635 21097 17647 21100
rect 17589 21091 17647 21097
rect 17678 21088 17684 21100
rect 17736 21128 17742 21140
rect 18049 21131 18107 21137
rect 18049 21128 18061 21131
rect 17736 21100 18061 21128
rect 17736 21088 17742 21100
rect 18049 21097 18061 21100
rect 18095 21128 18107 21131
rect 18138 21128 18144 21140
rect 18095 21100 18144 21128
rect 18095 21097 18107 21100
rect 18049 21091 18107 21097
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 23661 21131 23719 21137
rect 23661 21097 23673 21131
rect 23707 21128 23719 21131
rect 23750 21128 23756 21140
rect 23707 21100 23756 21128
rect 23707 21097 23719 21100
rect 23661 21091 23719 21097
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 24026 21088 24032 21140
rect 24084 21128 24090 21140
rect 24121 21131 24179 21137
rect 24121 21128 24133 21131
rect 24084 21100 24133 21128
rect 24084 21088 24090 21100
rect 24121 21097 24133 21100
rect 24167 21128 24179 21131
rect 24486 21128 24492 21140
rect 24167 21100 24492 21128
rect 24167 21097 24179 21100
rect 24121 21091 24179 21097
rect 24486 21088 24492 21100
rect 24544 21088 24550 21140
rect 25222 21128 25228 21140
rect 25183 21100 25228 21128
rect 25222 21088 25228 21100
rect 25280 21088 25286 21140
rect 25317 21131 25375 21137
rect 25317 21097 25329 21131
rect 25363 21128 25375 21131
rect 25590 21128 25596 21140
rect 25363 21100 25596 21128
rect 25363 21097 25375 21100
rect 25317 21091 25375 21097
rect 25590 21088 25596 21100
rect 25648 21088 25654 21140
rect 28626 21088 28632 21140
rect 28684 21128 28690 21140
rect 29273 21131 29331 21137
rect 29273 21128 29285 21131
rect 28684 21100 29285 21128
rect 28684 21088 28690 21100
rect 29273 21097 29285 21100
rect 29319 21128 29331 21131
rect 29730 21128 29736 21140
rect 29319 21100 29736 21128
rect 29319 21097 29331 21100
rect 29273 21091 29331 21097
rect 29730 21088 29736 21100
rect 29788 21088 29794 21140
rect 30098 21088 30104 21140
rect 30156 21128 30162 21140
rect 31021 21131 31079 21137
rect 31021 21128 31033 21131
rect 30156 21100 31033 21128
rect 30156 21088 30162 21100
rect 31021 21097 31033 21100
rect 31067 21097 31079 21131
rect 31570 21128 31576 21140
rect 31531 21100 31576 21128
rect 31021 21091 31079 21097
rect 31570 21088 31576 21100
rect 31628 21088 31634 21140
rect 31846 21088 31852 21140
rect 31904 21128 31910 21140
rect 32125 21131 32183 21137
rect 32125 21128 32137 21131
rect 31904 21100 32137 21128
rect 31904 21088 31910 21100
rect 32125 21097 32137 21100
rect 32171 21097 32183 21131
rect 32950 21128 32956 21140
rect 32911 21100 32956 21128
rect 32125 21091 32183 21097
rect 32950 21088 32956 21100
rect 33008 21088 33014 21140
rect 33321 21131 33379 21137
rect 33321 21097 33333 21131
rect 33367 21128 33379 21131
rect 33594 21128 33600 21140
rect 33367 21100 33600 21128
rect 33367 21097 33379 21100
rect 33321 21091 33379 21097
rect 33594 21088 33600 21100
rect 33652 21128 33658 21140
rect 33652 21100 34928 21128
rect 33652 21088 33658 21100
rect 13078 21020 13084 21072
rect 13136 21060 13142 21072
rect 13256 21063 13314 21069
rect 13256 21060 13268 21063
rect 13136 21032 13268 21060
rect 13136 21020 13142 21032
rect 13256 21029 13268 21032
rect 13302 21060 13314 21063
rect 14734 21060 14740 21072
rect 13302 21032 14740 21060
rect 13302 21029 13314 21032
rect 13256 21023 13314 21029
rect 14734 21020 14740 21032
rect 14792 21020 14798 21072
rect 15105 21063 15163 21069
rect 15105 21029 15117 21063
rect 15151 21060 15163 21063
rect 15948 21060 15976 21088
rect 15151 21032 15976 21060
rect 22548 21063 22606 21069
rect 15151 21029 15163 21032
rect 15105 21023 15163 21029
rect 22548 21029 22560 21063
rect 22594 21060 22606 21063
rect 22738 21060 22744 21072
rect 22594 21032 22744 21060
rect 22594 21029 22606 21032
rect 22548 21023 22606 21029
rect 22738 21020 22744 21032
rect 22796 21020 22802 21072
rect 28721 21063 28779 21069
rect 28721 21029 28733 21063
rect 28767 21060 28779 21063
rect 29178 21060 29184 21072
rect 28767 21032 29184 21060
rect 28767 21029 28779 21032
rect 28721 21023 28779 21029
rect 29178 21020 29184 21032
rect 29236 21020 29242 21072
rect 29908 21063 29966 21069
rect 29908 21029 29920 21063
rect 29954 21060 29966 21063
rect 31588 21060 31616 21088
rect 29954 21032 31616 21060
rect 34900 21060 34928 21100
rect 35158 21088 35164 21140
rect 35216 21128 35222 21140
rect 35345 21131 35403 21137
rect 35345 21128 35357 21131
rect 35216 21100 35357 21128
rect 35216 21088 35222 21100
rect 35345 21097 35357 21100
rect 35391 21097 35403 21131
rect 35618 21128 35624 21140
rect 35579 21100 35624 21128
rect 35345 21091 35403 21097
rect 35618 21088 35624 21100
rect 35676 21088 35682 21140
rect 36173 21063 36231 21069
rect 36173 21060 36185 21063
rect 34900 21032 36185 21060
rect 29954 21029 29966 21032
rect 29908 21023 29966 21029
rect 36173 21029 36185 21032
rect 36219 21029 36231 21063
rect 36173 21023 36231 21029
rect 16476 20995 16534 21001
rect 16476 20961 16488 20995
rect 16522 20992 16534 20995
rect 17310 20992 17316 21004
rect 16522 20964 17316 20992
rect 16522 20961 16534 20964
rect 16476 20955 16534 20961
rect 17310 20952 17316 20964
rect 17368 20952 17374 21004
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18417 20995 18475 21001
rect 18417 20992 18429 20995
rect 18012 20964 18429 20992
rect 18012 20952 18018 20964
rect 18417 20961 18429 20964
rect 18463 20961 18475 20995
rect 21174 20992 21180 21004
rect 21135 20964 21180 20992
rect 18417 20955 18475 20961
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 22189 20995 22247 21001
rect 22189 20992 22201 20995
rect 21744 20964 22201 20992
rect 12986 20924 12992 20936
rect 12947 20896 12992 20924
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 16206 20924 16212 20936
rect 16167 20896 16212 20924
rect 16206 20884 16212 20896
rect 16264 20884 16270 20936
rect 20162 20924 20168 20936
rect 20123 20896 20168 20924
rect 20162 20884 20168 20896
rect 20220 20884 20226 20936
rect 20346 20884 20352 20936
rect 20404 20924 20410 20936
rect 20533 20927 20591 20933
rect 20533 20924 20545 20927
rect 20404 20896 20545 20924
rect 20404 20884 20410 20896
rect 20533 20893 20545 20896
rect 20579 20924 20591 20927
rect 21358 20924 21364 20936
rect 20579 20896 21364 20924
rect 20579 20893 20591 20896
rect 20533 20887 20591 20893
rect 21358 20884 21364 20896
rect 21416 20924 21422 20936
rect 21744 20933 21772 20964
rect 22189 20961 22201 20964
rect 22235 20992 22247 20995
rect 22281 20995 22339 21001
rect 22281 20992 22293 20995
rect 22235 20964 22293 20992
rect 22235 20961 22247 20964
rect 22189 20955 22247 20961
rect 22281 20961 22293 20964
rect 22327 20992 22339 20995
rect 23106 20992 23112 21004
rect 22327 20964 23112 20992
rect 22327 20961 22339 20964
rect 22281 20955 22339 20961
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 24489 20995 24547 21001
rect 24489 20961 24501 20995
rect 24535 20992 24547 20995
rect 24670 20992 24676 21004
rect 24535 20964 24676 20992
rect 24535 20961 24547 20964
rect 24489 20955 24547 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 27062 21001 27068 21004
rect 27056 20992 27068 21001
rect 27023 20964 27068 20992
rect 27056 20955 27068 20964
rect 27062 20952 27068 20955
rect 27120 20952 27126 21004
rect 34238 20992 34244 21004
rect 34199 20964 34244 20992
rect 34238 20952 34244 20964
rect 34296 20952 34302 21004
rect 21729 20927 21787 20933
rect 21729 20924 21741 20927
rect 21416 20896 21741 20924
rect 21416 20884 21422 20896
rect 21729 20893 21741 20896
rect 21775 20893 21787 20927
rect 21729 20887 21787 20893
rect 25130 20884 25136 20936
rect 25188 20924 25194 20936
rect 25409 20927 25467 20933
rect 25409 20924 25421 20927
rect 25188 20896 25421 20924
rect 25188 20884 25194 20896
rect 25409 20893 25421 20896
rect 25455 20893 25467 20927
rect 26786 20924 26792 20936
rect 26747 20896 26792 20924
rect 25409 20887 25467 20893
rect 26786 20884 26792 20896
rect 26844 20884 26850 20936
rect 29641 20927 29699 20933
rect 29641 20893 29653 20927
rect 29687 20893 29699 20927
rect 29641 20887 29699 20893
rect 21358 20788 21364 20800
rect 21319 20760 21364 20788
rect 21358 20748 21364 20760
rect 21416 20748 21422 20800
rect 24857 20791 24915 20797
rect 24857 20757 24869 20791
rect 24903 20788 24915 20791
rect 26053 20791 26111 20797
rect 26053 20788 26065 20791
rect 24903 20760 26065 20788
rect 24903 20757 24915 20760
rect 24857 20751 24915 20757
rect 26053 20757 26065 20760
rect 26099 20788 26111 20791
rect 26234 20788 26240 20800
rect 26099 20760 26240 20788
rect 26099 20757 26111 20760
rect 26053 20751 26111 20757
rect 26234 20748 26240 20760
rect 26292 20748 26298 20800
rect 27890 20748 27896 20800
rect 27948 20788 27954 20800
rect 28169 20791 28227 20797
rect 28169 20788 28181 20791
rect 27948 20760 28181 20788
rect 27948 20748 27954 20760
rect 28169 20757 28181 20760
rect 28215 20757 28227 20791
rect 29656 20788 29684 20887
rect 33134 20884 33140 20936
rect 33192 20924 33198 20936
rect 33505 20927 33563 20933
rect 33505 20924 33517 20927
rect 33192 20896 33517 20924
rect 33192 20884 33198 20896
rect 33505 20893 33517 20896
rect 33551 20893 33563 20927
rect 33505 20887 33563 20893
rect 33686 20884 33692 20936
rect 33744 20924 33750 20936
rect 33828 20927 33886 20933
rect 33828 20924 33840 20927
rect 33744 20896 33840 20924
rect 33744 20884 33750 20896
rect 33828 20893 33840 20896
rect 33874 20893 33886 20927
rect 33828 20887 33886 20893
rect 33962 20884 33968 20936
rect 34020 20924 34026 20936
rect 34020 20896 34065 20924
rect 34020 20884 34026 20896
rect 29822 20788 29828 20800
rect 29656 20760 29828 20788
rect 28169 20751 28227 20757
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 12986 20544 12992 20596
rect 13044 20584 13050 20596
rect 13357 20587 13415 20593
rect 13357 20584 13369 20587
rect 13044 20556 13369 20584
rect 13044 20544 13050 20556
rect 13357 20553 13369 20556
rect 13403 20553 13415 20587
rect 15286 20584 15292 20596
rect 15247 20556 15292 20584
rect 13357 20547 13415 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 15896 20556 16129 20584
rect 15896 20544 15902 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 16206 20544 16212 20596
rect 16264 20584 16270 20596
rect 17681 20587 17739 20593
rect 17681 20584 17693 20587
rect 16264 20556 17693 20584
rect 16264 20544 16270 20556
rect 17681 20553 17693 20556
rect 17727 20584 17739 20587
rect 18046 20584 18052 20596
rect 17727 20556 18052 20584
rect 17727 20553 17739 20556
rect 17681 20547 17739 20553
rect 18046 20544 18052 20556
rect 18104 20544 18110 20596
rect 19426 20584 19432 20596
rect 19387 20556 19432 20584
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20898 20584 20904 20596
rect 20036 20556 20904 20584
rect 20036 20544 20042 20556
rect 20898 20544 20904 20556
rect 20956 20584 20962 20596
rect 21913 20587 21971 20593
rect 21913 20584 21925 20587
rect 20956 20556 21925 20584
rect 20956 20544 20962 20556
rect 21913 20553 21925 20556
rect 21959 20553 21971 20587
rect 21913 20547 21971 20553
rect 22373 20587 22431 20593
rect 22373 20553 22385 20587
rect 22419 20584 22431 20587
rect 22738 20584 22744 20596
rect 22419 20556 22744 20584
rect 22419 20553 22431 20556
rect 22373 20547 22431 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 24949 20587 25007 20593
rect 24949 20553 24961 20587
rect 24995 20584 25007 20587
rect 25222 20584 25228 20596
rect 24995 20556 25228 20584
rect 24995 20553 25007 20556
rect 24949 20547 25007 20553
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 25317 20587 25375 20593
rect 25317 20553 25329 20587
rect 25363 20584 25375 20587
rect 25590 20584 25596 20596
rect 25363 20556 25596 20584
rect 25363 20553 25375 20556
rect 25317 20547 25375 20553
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 27614 20584 27620 20596
rect 27575 20556 27620 20584
rect 27614 20544 27620 20556
rect 27672 20544 27678 20596
rect 28718 20544 28724 20596
rect 28776 20584 28782 20596
rect 28776 20556 29132 20584
rect 28776 20544 28782 20556
rect 13078 20516 13084 20528
rect 13039 20488 13084 20516
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 17221 20519 17279 20525
rect 17221 20485 17233 20519
rect 17267 20516 17279 20519
rect 17310 20516 17316 20528
rect 17267 20488 17316 20516
rect 17267 20485 17279 20488
rect 17221 20479 17279 20485
rect 17310 20476 17316 20488
rect 17368 20516 17374 20528
rect 17862 20516 17868 20528
rect 17368 20488 17868 20516
rect 17368 20476 17374 20488
rect 17862 20476 17868 20488
rect 17920 20476 17926 20528
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20448 13875 20451
rect 13863 20420 14044 20448
rect 13863 20417 13875 20420
rect 13817 20411 13875 20417
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 13906 20380 13912 20392
rect 13688 20352 13912 20380
rect 13688 20340 13694 20352
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 14016 20380 14044 20420
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 15988 20420 16681 20448
rect 15988 20408 15994 20420
rect 16669 20417 16681 20420
rect 16715 20448 16727 20451
rect 16942 20448 16948 20460
rect 16715 20420 16948 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 18064 20457 18092 20544
rect 19518 20516 19524 20528
rect 19479 20488 19524 20516
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 20070 20448 20076 20460
rect 20031 20420 20076 20448
rect 18049 20411 18107 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 23109 20451 23167 20457
rect 23109 20417 23121 20451
rect 23155 20448 23167 20451
rect 24302 20448 24308 20460
rect 23155 20420 24308 20448
rect 23155 20417 23167 20420
rect 23109 20411 23167 20417
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 26234 20408 26240 20460
rect 26292 20448 26298 20460
rect 26513 20451 26571 20457
rect 26513 20448 26525 20451
rect 26292 20420 26525 20448
rect 26292 20408 26298 20420
rect 26513 20417 26525 20420
rect 26559 20417 26571 20451
rect 26513 20411 26571 20417
rect 26602 20408 26608 20460
rect 26660 20448 26666 20460
rect 27062 20448 27068 20460
rect 26660 20420 27068 20448
rect 26660 20408 26666 20420
rect 27062 20408 27068 20420
rect 27120 20408 27126 20460
rect 27522 20408 27528 20460
rect 27580 20408 27586 20460
rect 28261 20451 28319 20457
rect 28261 20417 28273 20451
rect 28307 20417 28319 20451
rect 28261 20411 28319 20417
rect 14182 20389 14188 20392
rect 14176 20380 14188 20389
rect 14016 20352 14188 20380
rect 14176 20343 14188 20352
rect 14182 20340 14188 20343
rect 14240 20340 14246 20392
rect 17402 20340 17408 20392
rect 17460 20380 17466 20392
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 17460 20352 17877 20380
rect 17460 20340 17466 20352
rect 17865 20349 17877 20352
rect 17911 20349 17923 20383
rect 17865 20343 17923 20349
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 18305 20383 18363 20389
rect 18305 20380 18317 20383
rect 18196 20352 18317 20380
rect 18196 20340 18202 20352
rect 18305 20349 18317 20352
rect 18351 20349 18363 20383
rect 19886 20380 19892 20392
rect 19847 20352 19892 20380
rect 18305 20343 18363 20349
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 20346 20340 20352 20392
rect 20404 20380 20410 20392
rect 20533 20383 20591 20389
rect 20533 20380 20545 20383
rect 20404 20352 20545 20380
rect 20404 20340 20410 20352
rect 20533 20349 20545 20352
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 23658 20340 23664 20392
rect 23716 20380 23722 20392
rect 24029 20383 24087 20389
rect 24029 20380 24041 20383
rect 23716 20352 24041 20380
rect 23716 20340 23722 20352
rect 24029 20349 24041 20352
rect 24075 20349 24087 20383
rect 24029 20343 24087 20349
rect 25961 20383 26019 20389
rect 25961 20349 25973 20383
rect 26007 20380 26019 20383
rect 26421 20383 26479 20389
rect 26421 20380 26433 20383
rect 26007 20352 26433 20380
rect 26007 20349 26019 20352
rect 25961 20343 26019 20349
rect 26421 20349 26433 20352
rect 26467 20380 26479 20383
rect 27540 20380 27568 20408
rect 26467 20352 27568 20380
rect 28276 20380 28304 20411
rect 28721 20383 28779 20389
rect 28721 20380 28733 20383
rect 28276 20352 28733 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 28721 20349 28733 20352
rect 28767 20380 28779 20383
rect 28994 20380 29000 20392
rect 28767 20352 29000 20380
rect 28767 20349 28779 20352
rect 28721 20343 28779 20349
rect 28994 20340 29000 20352
rect 29052 20340 29058 20392
rect 16022 20312 16028 20324
rect 15935 20284 16028 20312
rect 16022 20272 16028 20284
rect 16080 20312 16086 20324
rect 16577 20315 16635 20321
rect 16577 20312 16589 20315
rect 16080 20284 16589 20312
rect 16080 20272 16086 20284
rect 16577 20281 16589 20284
rect 16623 20281 16635 20315
rect 17954 20312 17960 20324
rect 16577 20275 16635 20281
rect 17512 20284 17960 20312
rect 17512 20256 17540 20284
rect 17954 20272 17960 20284
rect 18012 20272 18018 20324
rect 20778 20315 20836 20321
rect 20778 20312 20790 20315
rect 20548 20284 20790 20312
rect 20548 20256 20576 20284
rect 20778 20281 20790 20284
rect 20824 20281 20836 20315
rect 20778 20275 20836 20281
rect 22741 20315 22799 20321
rect 22741 20281 22753 20315
rect 22787 20312 22799 20315
rect 23106 20312 23112 20324
rect 22787 20284 23112 20312
rect 22787 20281 22799 20284
rect 22741 20275 22799 20281
rect 23106 20272 23112 20284
rect 23164 20272 23170 20324
rect 24121 20315 24179 20321
rect 24121 20312 24133 20315
rect 23492 20284 24133 20312
rect 23492 20256 23520 20284
rect 24121 20281 24133 20284
rect 24167 20281 24179 20315
rect 24121 20275 24179 20281
rect 27525 20315 27583 20321
rect 27525 20281 27537 20315
rect 27571 20312 27583 20315
rect 27985 20315 28043 20321
rect 27985 20312 27997 20315
rect 27571 20284 27997 20312
rect 27571 20281 27583 20284
rect 27525 20275 27583 20281
rect 27985 20281 27997 20284
rect 28031 20312 28043 20315
rect 28166 20312 28172 20324
rect 28031 20284 28172 20312
rect 28031 20281 28043 20284
rect 27985 20275 28043 20281
rect 28166 20272 28172 20284
rect 28224 20272 28230 20324
rect 15657 20247 15715 20253
rect 15657 20213 15669 20247
rect 15703 20244 15715 20247
rect 16485 20247 16543 20253
rect 16485 20244 16497 20247
rect 15703 20216 16497 20244
rect 15703 20213 15715 20216
rect 15657 20207 15715 20213
rect 16485 20213 16497 20216
rect 16531 20244 16543 20247
rect 16666 20244 16672 20256
rect 16531 20216 16672 20244
rect 16531 20213 16543 20216
rect 16485 20207 16543 20213
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 17494 20244 17500 20256
rect 17455 20216 17500 20244
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 19978 20204 19984 20256
rect 20036 20244 20042 20256
rect 20036 20216 20081 20244
rect 20036 20204 20042 20216
rect 20530 20204 20536 20256
rect 20588 20204 20594 20256
rect 23474 20244 23480 20256
rect 23435 20216 23480 20244
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 23661 20247 23719 20253
rect 23661 20213 23673 20247
rect 23707 20244 23719 20247
rect 23750 20244 23756 20256
rect 23707 20216 23756 20244
rect 23707 20213 23719 20216
rect 23661 20207 23719 20213
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 26050 20244 26056 20256
rect 26011 20216 26056 20244
rect 26050 20204 26056 20216
rect 26108 20204 26114 20256
rect 28074 20244 28080 20256
rect 28035 20216 28080 20244
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 29104 20253 29132 20556
rect 29270 20544 29276 20596
rect 29328 20584 29334 20596
rect 31389 20587 31447 20593
rect 31389 20584 31401 20587
rect 29328 20556 31401 20584
rect 29328 20544 29334 20556
rect 31389 20553 31401 20556
rect 31435 20584 31447 20587
rect 31573 20587 31631 20593
rect 31573 20584 31585 20587
rect 31435 20556 31585 20584
rect 31435 20553 31447 20556
rect 31389 20547 31447 20553
rect 31573 20553 31585 20556
rect 31619 20553 31631 20587
rect 33686 20584 33692 20596
rect 33647 20556 33692 20584
rect 31573 20547 31631 20553
rect 33686 20544 33692 20556
rect 33744 20544 33750 20596
rect 33962 20584 33968 20596
rect 33923 20556 33968 20584
rect 33962 20544 33968 20556
rect 34020 20544 34026 20596
rect 34238 20544 34244 20596
rect 34296 20584 34302 20596
rect 34333 20587 34391 20593
rect 34333 20584 34345 20587
rect 34296 20556 34345 20584
rect 34296 20544 34302 20556
rect 34333 20553 34345 20556
rect 34379 20553 34391 20587
rect 34333 20547 34391 20553
rect 34790 20544 34796 20596
rect 34848 20584 34854 20596
rect 36078 20584 36084 20596
rect 34848 20556 36084 20584
rect 34848 20544 34854 20556
rect 36078 20544 36084 20556
rect 36136 20544 36142 20596
rect 29730 20408 29736 20460
rect 29788 20448 29794 20460
rect 29788 20420 29833 20448
rect 29788 20408 29794 20420
rect 31662 20408 31668 20460
rect 31720 20448 31726 20460
rect 31846 20448 31852 20460
rect 31720 20420 31852 20448
rect 31720 20408 31726 20420
rect 31846 20408 31852 20420
rect 31904 20448 31910 20460
rect 31948 20451 32006 20457
rect 31948 20448 31960 20451
rect 31904 20420 31960 20448
rect 31904 20408 31910 20420
rect 31948 20417 31960 20420
rect 31994 20417 32006 20451
rect 31948 20411 32006 20417
rect 29270 20380 29276 20392
rect 29231 20352 29276 20380
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 29362 20340 29368 20392
rect 29420 20380 29426 20392
rect 30006 20380 30012 20392
rect 29420 20352 30012 20380
rect 29420 20340 29426 20352
rect 30006 20340 30012 20352
rect 30064 20340 30070 20392
rect 35069 20383 35127 20389
rect 35069 20349 35081 20383
rect 35115 20349 35127 20383
rect 35069 20343 35127 20349
rect 31754 20272 31760 20324
rect 31812 20312 31818 20324
rect 32186 20315 32244 20321
rect 32186 20312 32198 20315
rect 31812 20284 32198 20312
rect 31812 20272 31818 20284
rect 32186 20281 32198 20284
rect 32232 20281 32244 20315
rect 35084 20312 35112 20343
rect 35158 20340 35164 20392
rect 35216 20380 35222 20392
rect 35336 20383 35394 20389
rect 35336 20380 35348 20383
rect 35216 20352 35348 20380
rect 35216 20340 35222 20352
rect 35336 20349 35348 20352
rect 35382 20380 35394 20383
rect 35894 20380 35900 20392
rect 35382 20352 35900 20380
rect 35382 20349 35394 20352
rect 35336 20343 35394 20349
rect 35894 20340 35900 20352
rect 35952 20340 35958 20392
rect 35434 20312 35440 20324
rect 35084 20284 35440 20312
rect 32186 20275 32244 20281
rect 35434 20272 35440 20284
rect 35492 20312 35498 20324
rect 36725 20315 36783 20321
rect 36725 20312 36737 20315
rect 35492 20284 36737 20312
rect 35492 20272 35498 20284
rect 36725 20281 36737 20284
rect 36771 20281 36783 20315
rect 36725 20275 36783 20281
rect 29089 20247 29147 20253
rect 29089 20213 29101 20247
rect 29135 20244 29147 20247
rect 29730 20244 29736 20256
rect 29788 20253 29794 20256
rect 29135 20216 29736 20244
rect 29135 20213 29147 20216
rect 29089 20207 29147 20213
rect 29730 20204 29736 20216
rect 29788 20244 29797 20253
rect 31110 20244 31116 20256
rect 29788 20216 29833 20244
rect 31071 20216 31116 20244
rect 29788 20207 29797 20216
rect 29788 20204 29794 20207
rect 31110 20204 31116 20216
rect 31168 20204 31174 20256
rect 31573 20247 31631 20253
rect 31573 20213 31585 20247
rect 31619 20244 31631 20247
rect 32950 20244 32956 20256
rect 31619 20216 32956 20244
rect 31619 20213 31631 20216
rect 31573 20207 31631 20213
rect 32950 20204 32956 20216
rect 33008 20204 33014 20256
rect 33318 20244 33324 20256
rect 33279 20216 33324 20244
rect 33318 20204 33324 20216
rect 33376 20204 33382 20256
rect 36078 20204 36084 20256
rect 36136 20244 36142 20256
rect 36449 20247 36507 20253
rect 36449 20244 36461 20247
rect 36136 20216 36461 20244
rect 36136 20204 36142 20216
rect 36449 20213 36461 20216
rect 36495 20213 36507 20247
rect 37274 20244 37280 20256
rect 37235 20216 37280 20244
rect 36449 20207 36507 20213
rect 37274 20204 37280 20216
rect 37332 20204 37338 20256
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 13906 20040 13912 20052
rect 13867 20012 13912 20040
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 16942 20040 16948 20052
rect 16903 20012 16948 20040
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 17402 20040 17408 20052
rect 17363 20012 17408 20040
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 18877 20043 18935 20049
rect 18877 20040 18889 20043
rect 17920 20012 18889 20040
rect 17920 20000 17926 20012
rect 18877 20009 18889 20012
rect 18923 20009 18935 20043
rect 18877 20003 18935 20009
rect 19613 20043 19671 20049
rect 19613 20009 19625 20043
rect 19659 20040 19671 20043
rect 19978 20040 19984 20052
rect 19659 20012 19984 20040
rect 19659 20009 19671 20012
rect 19613 20003 19671 20009
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 21174 20040 21180 20052
rect 21135 20012 21180 20040
rect 21174 20000 21180 20012
rect 21232 20040 21238 20052
rect 21913 20043 21971 20049
rect 21913 20040 21925 20043
rect 21232 20012 21925 20040
rect 21232 20000 21238 20012
rect 21913 20009 21925 20012
rect 21959 20009 21971 20043
rect 23658 20040 23664 20052
rect 23619 20012 23664 20040
rect 21913 20003 21971 20009
rect 23658 20000 23664 20012
rect 23716 20000 23722 20052
rect 24026 20040 24032 20052
rect 23987 20012 24032 20040
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 25130 20040 25136 20052
rect 25091 20012 25136 20040
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 26145 20043 26203 20049
rect 26145 20009 26157 20043
rect 26191 20040 26203 20043
rect 26602 20040 26608 20052
rect 26191 20012 26608 20040
rect 26191 20009 26203 20012
rect 26145 20003 26203 20009
rect 26602 20000 26608 20012
rect 26660 20000 26666 20052
rect 28994 20040 29000 20052
rect 28955 20012 29000 20040
rect 28994 20000 29000 20012
rect 29052 20000 29058 20052
rect 29733 20043 29791 20049
rect 29733 20009 29745 20043
rect 29779 20040 29791 20043
rect 31205 20043 31263 20049
rect 31205 20040 31217 20043
rect 29779 20012 31217 20040
rect 29779 20009 29791 20012
rect 29733 20003 29791 20009
rect 31205 20009 31217 20012
rect 31251 20040 31263 20043
rect 31570 20040 31576 20052
rect 31251 20012 31576 20040
rect 31251 20009 31263 20012
rect 31205 20003 31263 20009
rect 31570 20000 31576 20012
rect 31628 20000 31634 20052
rect 31846 20000 31852 20052
rect 31904 20040 31910 20052
rect 32309 20043 32367 20049
rect 32309 20040 32321 20043
rect 31904 20012 32321 20040
rect 31904 20000 31910 20012
rect 32309 20009 32321 20012
rect 32355 20009 32367 20043
rect 32309 20003 32367 20009
rect 33226 20000 33232 20052
rect 33284 20040 33290 20052
rect 33419 20043 33477 20049
rect 33419 20040 33431 20043
rect 33284 20012 33431 20040
rect 33284 20000 33290 20012
rect 33419 20009 33431 20012
rect 33465 20040 33477 20043
rect 33686 20040 33692 20052
rect 33465 20012 33692 20040
rect 33465 20009 33477 20012
rect 33419 20003 33477 20009
rect 33686 20000 33692 20012
rect 33744 20000 33750 20052
rect 34330 20000 34336 20052
rect 34388 20040 34394 20052
rect 34793 20043 34851 20049
rect 34793 20040 34805 20043
rect 34388 20012 34805 20040
rect 34388 20000 34394 20012
rect 34793 20009 34805 20012
rect 34839 20009 34851 20043
rect 35158 20040 35164 20052
rect 35119 20012 35164 20040
rect 34793 20003 34851 20009
rect 35158 20000 35164 20012
rect 35216 20000 35222 20052
rect 15556 19975 15614 19981
rect 15556 19941 15568 19975
rect 15602 19972 15614 19975
rect 16022 19972 16028 19984
rect 15602 19944 16028 19972
rect 15602 19941 15614 19944
rect 15556 19935 15614 19941
rect 16022 19932 16028 19944
rect 16080 19932 16086 19984
rect 16206 19932 16212 19984
rect 16264 19932 16270 19984
rect 16684 19972 16712 20000
rect 17586 19972 17592 19984
rect 16684 19944 17592 19972
rect 17586 19932 17592 19944
rect 17644 19972 17650 19984
rect 17742 19975 17800 19981
rect 17742 19972 17754 19975
rect 17644 19944 17754 19972
rect 17644 19932 17650 19944
rect 17742 19941 17754 19944
rect 17788 19941 17800 19975
rect 19886 19972 19892 19984
rect 19847 19944 19892 19972
rect 17742 19935 17800 19941
rect 19886 19932 19892 19944
rect 19944 19932 19950 19984
rect 23385 19975 23443 19981
rect 23385 19941 23397 19975
rect 23431 19972 23443 19975
rect 24302 19972 24308 19984
rect 23431 19944 24308 19972
rect 23431 19941 23443 19944
rect 23385 19935 23443 19941
rect 24302 19932 24308 19944
rect 24360 19972 24366 19984
rect 27525 19975 27583 19981
rect 24360 19944 24624 19972
rect 24360 19932 24366 19944
rect 16224 19904 16252 19932
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 16224 19876 17509 19904
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 22094 19864 22100 19916
rect 22152 19904 22158 19916
rect 22278 19904 22284 19916
rect 22152 19876 22284 19904
rect 22152 19864 22158 19876
rect 22278 19864 22284 19876
rect 22336 19864 22342 19916
rect 24394 19904 24400 19916
rect 24355 19876 24400 19904
rect 24394 19864 24400 19876
rect 24452 19864 24458 19916
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 15289 19839 15347 19845
rect 15289 19836 15301 19839
rect 14608 19808 15301 19836
rect 14608 19796 14614 19808
rect 15289 19805 15301 19808
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19836 21879 19839
rect 21867 19808 22140 19836
rect 21867 19805 21879 19808
rect 21821 19799 21879 19805
rect 22112 19768 22140 19808
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 22244 19808 22385 19836
rect 22244 19796 22250 19808
rect 22373 19805 22385 19808
rect 22419 19805 22431 19839
rect 22554 19836 22560 19848
rect 22373 19799 22431 19805
rect 22480 19808 22560 19836
rect 22480 19768 22508 19808
rect 22554 19796 22560 19808
rect 22612 19796 22618 19848
rect 24026 19796 24032 19848
rect 24084 19836 24090 19848
rect 24596 19845 24624 19944
rect 27525 19941 27537 19975
rect 27571 19972 27583 19975
rect 28074 19972 28080 19984
rect 27571 19944 28080 19972
rect 27571 19941 27583 19944
rect 27525 19935 27583 19941
rect 28074 19932 28080 19944
rect 28132 19932 28138 19984
rect 30098 19981 30104 19984
rect 30092 19972 30104 19981
rect 30059 19944 30104 19972
rect 30092 19935 30104 19944
rect 30098 19932 30104 19935
rect 30156 19932 30162 19984
rect 26510 19904 26516 19916
rect 26471 19876 26516 19904
rect 26510 19864 26516 19876
rect 26568 19864 26574 19916
rect 27890 19913 27896 19916
rect 27884 19904 27896 19913
rect 27851 19876 27896 19904
rect 27884 19867 27896 19876
rect 27890 19864 27896 19867
rect 27948 19864 27954 19916
rect 29822 19904 29828 19916
rect 29783 19876 29828 19904
rect 29822 19864 29828 19876
rect 29880 19864 29886 19916
rect 35986 19904 35992 19916
rect 33612 19876 35664 19904
rect 35947 19876 35992 19904
rect 24489 19839 24547 19845
rect 24489 19836 24501 19839
rect 24084 19808 24501 19836
rect 24084 19796 24090 19808
rect 24489 19805 24501 19808
rect 24535 19805 24547 19839
rect 24489 19799 24547 19805
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 26786 19796 26792 19848
rect 26844 19836 26850 19848
rect 27157 19839 27215 19845
rect 27157 19836 27169 19839
rect 26844 19808 27169 19836
rect 26844 19796 26850 19808
rect 27157 19805 27169 19808
rect 27203 19836 27215 19839
rect 27614 19836 27620 19848
rect 27203 19808 27620 19836
rect 27203 19805 27215 19808
rect 27157 19799 27215 19805
rect 27614 19796 27620 19808
rect 27672 19796 27678 19848
rect 32953 19839 33011 19845
rect 32953 19805 32965 19839
rect 32999 19805 33011 19839
rect 33410 19836 33416 19848
rect 33369 19808 33416 19836
rect 32953 19799 33011 19805
rect 22112 19740 22508 19768
rect 32968 19712 32996 19799
rect 33410 19796 33416 19808
rect 33468 19845 33474 19848
rect 33468 19839 33517 19845
rect 33468 19805 33471 19839
rect 33505 19836 33517 19839
rect 33612 19836 33640 19876
rect 33505 19808 33640 19836
rect 33505 19805 33517 19808
rect 33468 19799 33517 19805
rect 33468 19796 33474 19799
rect 33686 19796 33692 19848
rect 33744 19836 33750 19848
rect 33744 19808 33789 19836
rect 33744 19796 33750 19808
rect 34422 19728 34428 19780
rect 34480 19768 34486 19780
rect 35636 19777 35664 19876
rect 35986 19864 35992 19876
rect 36044 19864 36050 19916
rect 36081 19839 36139 19845
rect 36081 19805 36093 19839
rect 36127 19805 36139 19839
rect 36081 19799 36139 19805
rect 36265 19839 36323 19845
rect 36265 19805 36277 19839
rect 36311 19836 36323 19839
rect 36906 19836 36912 19848
rect 36311 19808 36912 19836
rect 36311 19805 36323 19808
rect 36265 19799 36323 19805
rect 35437 19771 35495 19777
rect 35437 19768 35449 19771
rect 34480 19740 35449 19768
rect 34480 19728 34486 19740
rect 35437 19737 35449 19740
rect 35483 19737 35495 19771
rect 35437 19731 35495 19737
rect 35621 19771 35679 19777
rect 35621 19737 35633 19771
rect 35667 19737 35679 19771
rect 35621 19731 35679 19737
rect 19245 19703 19303 19709
rect 19245 19669 19257 19703
rect 19291 19700 19303 19703
rect 19978 19700 19984 19712
rect 19291 19672 19984 19700
rect 19291 19669 19303 19672
rect 19245 19663 19303 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 20530 19700 20536 19712
rect 20491 19672 20536 19700
rect 20530 19660 20536 19672
rect 20588 19660 20594 19712
rect 26234 19660 26240 19712
rect 26292 19700 26298 19712
rect 26697 19703 26755 19709
rect 26697 19700 26709 19703
rect 26292 19672 26709 19700
rect 26292 19660 26298 19672
rect 26697 19669 26709 19672
rect 26743 19669 26755 19703
rect 29362 19700 29368 19712
rect 29323 19672 29368 19700
rect 26697 19663 26755 19669
rect 29362 19660 29368 19672
rect 29420 19660 29426 19712
rect 32861 19703 32919 19709
rect 32861 19669 32873 19703
rect 32907 19700 32919 19703
rect 32950 19700 32956 19712
rect 32907 19672 32956 19700
rect 32907 19669 32919 19672
rect 32861 19663 32919 19669
rect 32950 19660 32956 19672
rect 33008 19660 33014 19712
rect 35452 19700 35480 19731
rect 36096 19700 36124 19799
rect 36906 19796 36912 19808
rect 36964 19796 36970 19848
rect 35452 19672 36124 19700
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 15933 19499 15991 19505
rect 15933 19465 15945 19499
rect 15979 19496 15991 19499
rect 16022 19496 16028 19508
rect 15979 19468 16028 19496
rect 15979 19465 15991 19468
rect 15933 19459 15991 19465
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 17586 19496 17592 19508
rect 17547 19468 17592 19496
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 18046 19456 18052 19508
rect 18104 19496 18110 19508
rect 18233 19499 18291 19505
rect 18233 19496 18245 19499
rect 18104 19468 18245 19496
rect 18104 19456 18110 19468
rect 18233 19465 18245 19468
rect 18279 19496 18291 19499
rect 18601 19499 18659 19505
rect 18601 19496 18613 19499
rect 18279 19468 18613 19496
rect 18279 19465 18291 19468
rect 18233 19459 18291 19465
rect 18601 19465 18613 19468
rect 18647 19465 18659 19499
rect 20346 19496 20352 19508
rect 18601 19459 18659 19465
rect 19996 19468 20352 19496
rect 13906 19320 13912 19372
rect 13964 19360 13970 19372
rect 14550 19360 14556 19372
rect 13964 19332 14556 19360
rect 13964 19320 13970 19332
rect 14550 19320 14556 19332
rect 14608 19320 14614 19372
rect 19996 19369 20024 19468
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 22005 19499 22063 19505
rect 22005 19465 22017 19499
rect 22051 19496 22063 19499
rect 22186 19496 22192 19508
rect 22051 19468 22192 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 22186 19456 22192 19468
rect 22244 19456 22250 19508
rect 26510 19496 26516 19508
rect 26471 19468 26516 19496
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 27890 19496 27896 19508
rect 27851 19468 27896 19496
rect 27890 19456 27896 19468
rect 27948 19456 27954 19508
rect 33042 19496 33048 19508
rect 32600 19468 33048 19496
rect 19521 19363 19579 19369
rect 19521 19329 19533 19363
rect 19567 19360 19579 19363
rect 19981 19363 20039 19369
rect 19981 19360 19993 19363
rect 19567 19332 19993 19360
rect 19567 19329 19579 19332
rect 19521 19323 19579 19329
rect 19981 19329 19993 19332
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 22554 19320 22560 19372
rect 22612 19360 22618 19372
rect 24765 19363 24823 19369
rect 24765 19360 24777 19363
rect 22612 19332 24777 19360
rect 22612 19320 22618 19332
rect 24765 19329 24777 19332
rect 24811 19329 24823 19363
rect 28166 19360 28172 19372
rect 28127 19332 28172 19360
rect 24765 19323 24823 19329
rect 14820 19295 14878 19301
rect 14820 19292 14832 19295
rect 14752 19264 14832 19292
rect 14461 19227 14519 19233
rect 14461 19193 14473 19227
rect 14507 19224 14519 19227
rect 14752 19224 14780 19264
rect 14820 19261 14832 19264
rect 14866 19292 14878 19295
rect 15102 19292 15108 19304
rect 14866 19264 15108 19292
rect 14866 19261 14878 19264
rect 14820 19255 14878 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 22002 19252 22008 19304
rect 22060 19292 22066 19304
rect 22189 19295 22247 19301
rect 22189 19292 22201 19295
rect 22060 19264 22201 19292
rect 22060 19252 22066 19264
rect 22189 19261 22201 19264
rect 22235 19292 22247 19295
rect 22741 19295 22799 19301
rect 22741 19292 22753 19295
rect 22235 19264 22753 19292
rect 22235 19261 22247 19264
rect 22189 19255 22247 19261
rect 22741 19261 22753 19264
rect 22787 19261 22799 19295
rect 22741 19255 22799 19261
rect 24118 19252 24124 19304
rect 24176 19292 24182 19304
rect 24578 19292 24584 19304
rect 24176 19264 24584 19292
rect 24176 19252 24182 19264
rect 24578 19252 24584 19264
rect 24636 19252 24642 19304
rect 24780 19292 24808 19323
rect 28166 19320 28172 19332
rect 28224 19320 28230 19372
rect 29730 19320 29736 19372
rect 29788 19360 29794 19372
rect 30282 19369 30288 19372
rect 29825 19363 29883 19369
rect 29825 19360 29837 19363
rect 29788 19332 29837 19360
rect 29788 19320 29794 19332
rect 29825 19329 29837 19332
rect 29871 19360 29883 19363
rect 30240 19363 30288 19369
rect 30240 19360 30252 19363
rect 29871 19332 30252 19360
rect 29871 19329 29883 19332
rect 29825 19323 29883 19329
rect 30240 19329 30252 19332
rect 30286 19329 30288 19363
rect 30240 19323 30288 19329
rect 30282 19320 30288 19323
rect 30340 19320 30346 19372
rect 30466 19369 30472 19372
rect 30423 19363 30472 19369
rect 30423 19329 30435 19363
rect 30469 19329 30472 19363
rect 30423 19323 30472 19329
rect 30466 19320 30472 19323
rect 30524 19320 30530 19372
rect 30653 19363 30711 19369
rect 30653 19329 30665 19363
rect 30699 19360 30711 19363
rect 31110 19360 31116 19372
rect 30699 19332 31116 19360
rect 30699 19329 30711 19332
rect 30653 19323 30711 19329
rect 25774 19292 25780 19304
rect 24780 19264 25360 19292
rect 25735 19264 25780 19292
rect 19886 19224 19892 19236
rect 14507 19196 14780 19224
rect 19799 19196 19892 19224
rect 14507 19193 14519 19196
rect 14461 19187 14519 19193
rect 19886 19184 19892 19196
rect 19944 19224 19950 19236
rect 20248 19227 20306 19233
rect 20248 19224 20260 19227
rect 19944 19196 20260 19224
rect 19944 19184 19950 19196
rect 20248 19193 20260 19196
rect 20294 19224 20306 19227
rect 21174 19224 21180 19236
rect 20294 19196 21180 19224
rect 20294 19193 20306 19196
rect 20248 19187 20306 19193
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 25332 19233 25360 19264
rect 25774 19252 25780 19264
rect 25832 19252 25838 19304
rect 26878 19292 26884 19304
rect 26791 19264 26884 19292
rect 26878 19252 26884 19264
rect 26936 19292 26942 19304
rect 27433 19295 27491 19301
rect 27433 19292 27445 19295
rect 26936 19264 27445 19292
rect 26936 19252 26942 19264
rect 27433 19261 27445 19264
rect 27479 19261 27491 19295
rect 29270 19292 29276 19304
rect 27433 19255 27491 19261
rect 28644 19264 29276 19292
rect 23477 19227 23535 19233
rect 23477 19193 23489 19227
rect 23523 19224 23535 19227
rect 25317 19227 25375 19233
rect 23523 19196 24532 19224
rect 23523 19193 23535 19196
rect 23477 19187 23535 19193
rect 24504 19168 24532 19196
rect 25317 19193 25329 19227
rect 25363 19224 25375 19227
rect 25363 19196 26004 19224
rect 25363 19193 25375 19196
rect 25317 19187 25375 19193
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 16206 19156 16212 19168
rect 14608 19128 16212 19156
rect 14608 19116 14614 19128
rect 16206 19116 16212 19128
rect 16264 19156 16270 19168
rect 16577 19159 16635 19165
rect 16577 19156 16589 19159
rect 16264 19128 16589 19156
rect 16264 19116 16270 19128
rect 16577 19125 16589 19128
rect 16623 19125 16635 19159
rect 16577 19119 16635 19125
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 21361 19159 21419 19165
rect 21361 19156 21373 19159
rect 20588 19128 21373 19156
rect 20588 19116 20594 19128
rect 21361 19125 21373 19128
rect 21407 19125 21419 19159
rect 21361 19119 21419 19125
rect 22373 19159 22431 19165
rect 22373 19125 22385 19159
rect 22419 19156 22431 19159
rect 23290 19156 23296 19168
rect 22419 19128 23296 19156
rect 22419 19125 22431 19128
rect 22373 19119 22431 19125
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 24026 19156 24032 19168
rect 23987 19128 24032 19156
rect 24026 19116 24032 19128
rect 24084 19116 24090 19168
rect 24210 19156 24216 19168
rect 24171 19128 24216 19156
rect 24210 19116 24216 19128
rect 24268 19116 24274 19168
rect 24486 19116 24492 19168
rect 24544 19156 24550 19168
rect 24581 19159 24639 19165
rect 24581 19156 24593 19159
rect 24544 19128 24593 19156
rect 24544 19116 24550 19128
rect 24581 19125 24593 19128
rect 24627 19125 24639 19159
rect 24581 19119 24639 19125
rect 24670 19116 24676 19168
rect 24728 19156 24734 19168
rect 25685 19159 25743 19165
rect 24728 19128 24773 19156
rect 24728 19116 24734 19128
rect 25685 19125 25697 19159
rect 25731 19156 25743 19159
rect 25774 19156 25780 19168
rect 25731 19128 25780 19156
rect 25731 19125 25743 19128
rect 25685 19119 25743 19125
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 25976 19165 26004 19196
rect 28644 19168 28672 19264
rect 29270 19252 29276 19264
rect 29328 19292 29334 19304
rect 29917 19295 29975 19301
rect 29917 19292 29929 19295
rect 29328 19264 29929 19292
rect 29328 19252 29334 19264
rect 29917 19261 29929 19264
rect 29963 19261 29975 19295
rect 30668 19292 30696 19323
rect 31110 19320 31116 19332
rect 31168 19320 31174 19372
rect 29917 19255 29975 19261
rect 30015 19264 30696 19292
rect 29089 19227 29147 19233
rect 29089 19193 29101 19227
rect 29135 19224 29147 19227
rect 29178 19224 29184 19236
rect 29135 19196 29184 19224
rect 29135 19193 29147 19196
rect 29089 19187 29147 19193
rect 29178 19184 29184 19196
rect 29236 19224 29242 19236
rect 30015 19224 30043 19264
rect 30742 19252 30748 19304
rect 30800 19292 30806 19304
rect 32600 19292 32628 19468
rect 33042 19456 33048 19468
rect 33100 19496 33106 19508
rect 33226 19496 33232 19508
rect 33100 19468 33232 19496
rect 33100 19456 33106 19468
rect 33226 19456 33232 19468
rect 33284 19456 33290 19508
rect 33410 19360 33416 19372
rect 33060 19332 33416 19360
rect 30800 19264 32628 19292
rect 32677 19295 32735 19301
rect 30800 19252 30806 19264
rect 32677 19261 32689 19295
rect 32723 19292 32735 19295
rect 33060 19292 33088 19332
rect 33410 19320 33416 19332
rect 33468 19320 33474 19372
rect 34701 19363 34759 19369
rect 34701 19329 34713 19363
rect 34747 19360 34759 19363
rect 35434 19360 35440 19372
rect 34747 19332 35440 19360
rect 34747 19329 34759 19332
rect 34701 19323 34759 19329
rect 35434 19320 35440 19332
rect 35492 19320 35498 19372
rect 32723 19264 33088 19292
rect 35704 19295 35762 19301
rect 32723 19261 32735 19264
rect 32677 19255 32735 19261
rect 35704 19261 35716 19295
rect 35750 19261 35762 19295
rect 35704 19255 35762 19261
rect 33778 19224 33784 19236
rect 29236 19196 30043 19224
rect 31772 19196 33456 19224
rect 33739 19196 33784 19224
rect 29236 19184 29242 19196
rect 25961 19159 26019 19165
rect 25961 19125 25973 19159
rect 26007 19125 26019 19159
rect 27062 19156 27068 19168
rect 27023 19128 27068 19156
rect 25961 19119 26019 19125
rect 27062 19116 27068 19128
rect 27120 19116 27126 19168
rect 28626 19156 28632 19168
rect 28587 19128 28632 19156
rect 28626 19116 28632 19128
rect 28684 19116 28690 19168
rect 30282 19116 30288 19168
rect 30340 19156 30346 19168
rect 30742 19156 30748 19168
rect 30340 19128 30748 19156
rect 30340 19116 30346 19128
rect 30742 19116 30748 19128
rect 30800 19116 30806 19168
rect 30926 19116 30932 19168
rect 30984 19156 30990 19168
rect 31772 19165 31800 19196
rect 33428 19165 33456 19196
rect 33778 19184 33784 19196
rect 33836 19184 33842 19236
rect 35719 19224 35747 19255
rect 35986 19252 35992 19304
rect 36044 19292 36050 19304
rect 37093 19295 37151 19301
rect 37093 19292 37105 19295
rect 36044 19264 37105 19292
rect 36044 19252 36050 19264
rect 37093 19261 37105 19264
rect 37139 19261 37151 19295
rect 37093 19255 37151 19261
rect 36078 19224 36084 19236
rect 35719 19196 36084 19224
rect 36078 19184 36084 19196
rect 36136 19184 36142 19236
rect 31757 19159 31815 19165
rect 31757 19156 31769 19159
rect 30984 19128 31769 19156
rect 30984 19116 30990 19128
rect 31757 19125 31769 19128
rect 31803 19125 31815 19159
rect 31757 19119 31815 19125
rect 33413 19159 33471 19165
rect 33413 19125 33425 19159
rect 33459 19156 33471 19159
rect 33686 19156 33692 19168
rect 33459 19128 33692 19156
rect 33459 19125 33471 19128
rect 33413 19119 33471 19125
rect 33686 19116 33692 19128
rect 33744 19156 33750 19168
rect 34054 19156 34060 19168
rect 33744 19128 34060 19156
rect 33744 19116 33750 19128
rect 34054 19116 34060 19128
rect 34112 19116 34118 19168
rect 35345 19159 35403 19165
rect 35345 19125 35357 19159
rect 35391 19156 35403 19159
rect 36817 19159 36875 19165
rect 36817 19156 36829 19159
rect 35391 19128 36829 19156
rect 35391 19125 35403 19128
rect 35345 19119 35403 19125
rect 36817 19125 36829 19128
rect 36863 19156 36875 19159
rect 36906 19156 36912 19168
rect 36863 19128 36912 19156
rect 36863 19125 36875 19128
rect 36817 19119 36875 19125
rect 36906 19116 36912 19128
rect 36964 19116 36970 19168
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 14550 18952 14556 18964
rect 14511 18924 14556 18952
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 15565 18955 15623 18961
rect 15565 18921 15577 18955
rect 15611 18952 15623 18955
rect 16022 18952 16028 18964
rect 15611 18924 16028 18952
rect 15611 18921 15623 18924
rect 15565 18915 15623 18921
rect 16022 18912 16028 18924
rect 16080 18912 16086 18964
rect 22278 18912 22284 18964
rect 22336 18952 22342 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 22336 18924 22569 18952
rect 22336 18912 22342 18924
rect 22557 18921 22569 18924
rect 22603 18921 22615 18955
rect 22557 18915 22615 18921
rect 23382 18912 23388 18964
rect 23440 18952 23446 18964
rect 24213 18955 24271 18961
rect 24213 18952 24225 18955
rect 23440 18924 24225 18952
rect 23440 18912 23446 18924
rect 24213 18921 24225 18924
rect 24259 18952 24271 18955
rect 24394 18952 24400 18964
rect 24259 18924 24400 18952
rect 24259 18921 24271 18924
rect 24213 18915 24271 18921
rect 24394 18912 24400 18924
rect 24452 18912 24458 18964
rect 24581 18955 24639 18961
rect 24581 18921 24593 18955
rect 24627 18952 24639 18955
rect 24670 18952 24676 18964
rect 24627 18924 24676 18952
rect 24627 18921 24639 18924
rect 24581 18915 24639 18921
rect 24670 18912 24676 18924
rect 24728 18952 24734 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 24728 18924 24777 18952
rect 24728 18912 24734 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 25961 18955 26019 18961
rect 25961 18952 25973 18955
rect 25740 18924 25973 18952
rect 25740 18912 25746 18924
rect 25961 18921 25973 18924
rect 26007 18921 26019 18955
rect 26694 18952 26700 18964
rect 26655 18924 26700 18952
rect 25961 18915 26019 18921
rect 26694 18912 26700 18924
rect 26752 18912 26758 18964
rect 27617 18955 27675 18961
rect 27617 18921 27629 18955
rect 27663 18952 27675 18955
rect 27798 18952 27804 18964
rect 27663 18924 27804 18952
rect 27663 18921 27675 18924
rect 27617 18915 27675 18921
rect 27798 18912 27804 18924
rect 27856 18912 27862 18964
rect 28074 18912 28080 18964
rect 28132 18952 28138 18964
rect 28721 18955 28779 18961
rect 28721 18952 28733 18955
rect 28132 18924 28733 18952
rect 28132 18912 28138 18924
rect 28721 18921 28733 18924
rect 28767 18921 28779 18955
rect 29178 18952 29184 18964
rect 29139 18924 29184 18952
rect 28721 18915 28779 18921
rect 29178 18912 29184 18924
rect 29236 18912 29242 18964
rect 29914 18952 29920 18964
rect 29875 18924 29920 18952
rect 29914 18912 29920 18924
rect 29972 18952 29978 18964
rect 30466 18952 30472 18964
rect 29972 18924 30472 18952
rect 29972 18912 29978 18924
rect 30466 18912 30472 18924
rect 30524 18952 30530 18964
rect 30745 18955 30803 18961
rect 30745 18952 30757 18955
rect 30524 18924 30757 18952
rect 30524 18912 30530 18924
rect 30745 18921 30757 18924
rect 30791 18921 30803 18955
rect 30745 18915 30803 18921
rect 30837 18955 30895 18961
rect 30837 18921 30849 18955
rect 30883 18952 30895 18955
rect 30926 18952 30932 18964
rect 30883 18924 30932 18952
rect 30883 18921 30895 18924
rect 30837 18915 30895 18921
rect 30926 18912 30932 18924
rect 30984 18912 30990 18964
rect 31481 18955 31539 18961
rect 31481 18921 31493 18955
rect 31527 18952 31539 18955
rect 31662 18952 31668 18964
rect 31527 18924 31668 18952
rect 31527 18921 31539 18924
rect 31481 18915 31539 18921
rect 31662 18912 31668 18924
rect 31720 18912 31726 18964
rect 33137 18955 33195 18961
rect 33137 18921 33149 18955
rect 33183 18952 33195 18955
rect 33226 18952 33232 18964
rect 33183 18924 33232 18952
rect 33183 18921 33195 18924
rect 33137 18915 33195 18921
rect 33226 18912 33232 18924
rect 33284 18912 33290 18964
rect 34146 18912 34152 18964
rect 34204 18952 34210 18964
rect 34517 18955 34575 18961
rect 34517 18952 34529 18955
rect 34204 18924 34529 18952
rect 34204 18912 34210 18924
rect 34517 18921 34529 18924
rect 34563 18921 34575 18955
rect 34517 18915 34575 18921
rect 35710 18912 35716 18964
rect 35768 18952 35774 18964
rect 35989 18955 36047 18961
rect 35989 18952 36001 18955
rect 35768 18924 36001 18952
rect 35768 18912 35774 18924
rect 35989 18921 36001 18924
rect 36035 18952 36047 18955
rect 37182 18952 37188 18964
rect 36035 18924 37188 18952
rect 36035 18921 36047 18924
rect 35989 18915 36047 18921
rect 37182 18912 37188 18924
rect 37240 18912 37246 18964
rect 19334 18844 19340 18896
rect 19392 18884 19398 18896
rect 19705 18887 19763 18893
rect 19705 18884 19717 18887
rect 19392 18856 19717 18884
rect 19392 18844 19398 18856
rect 19705 18853 19717 18856
rect 19751 18884 19763 18887
rect 19886 18884 19892 18896
rect 19751 18856 19892 18884
rect 19751 18853 19763 18856
rect 19705 18847 19763 18853
rect 19886 18844 19892 18856
rect 19944 18844 19950 18896
rect 29089 18887 29147 18893
rect 29089 18853 29101 18887
rect 29135 18884 29147 18887
rect 29454 18884 29460 18896
rect 29135 18856 29460 18884
rect 29135 18853 29147 18856
rect 29089 18847 29147 18853
rect 29454 18844 29460 18856
rect 29512 18844 29518 18896
rect 36081 18887 36139 18893
rect 36081 18853 36093 18887
rect 36127 18884 36139 18887
rect 36170 18884 36176 18896
rect 36127 18856 36176 18884
rect 36127 18853 36139 18856
rect 36081 18847 36139 18853
rect 36170 18844 36176 18856
rect 36228 18844 36234 18896
rect 19610 18816 19616 18828
rect 19571 18788 19616 18816
rect 19610 18776 19616 18788
rect 19668 18816 19674 18828
rect 20530 18816 20536 18828
rect 19668 18788 20536 18816
rect 19668 18776 19674 18788
rect 20530 18776 20536 18788
rect 20588 18776 20594 18828
rect 21168 18819 21226 18825
rect 21168 18785 21180 18819
rect 21214 18816 21226 18819
rect 21542 18816 21548 18828
rect 21214 18788 21548 18816
rect 21214 18785 21226 18788
rect 21168 18779 21226 18785
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 23477 18819 23535 18825
rect 23477 18785 23489 18819
rect 23523 18816 23535 18819
rect 23842 18816 23848 18828
rect 23523 18788 23848 18816
rect 23523 18785 23535 18788
rect 23477 18779 23535 18785
rect 23842 18776 23848 18788
rect 23900 18776 23906 18828
rect 25130 18816 25136 18828
rect 25091 18788 25136 18816
rect 25130 18776 25136 18788
rect 25188 18776 25194 18828
rect 26510 18816 26516 18828
rect 26471 18788 26516 18816
rect 26510 18776 26516 18788
rect 26568 18776 26574 18828
rect 27706 18776 27712 18828
rect 27764 18816 27770 18828
rect 27801 18819 27859 18825
rect 27801 18816 27813 18819
rect 27764 18788 27813 18816
rect 27764 18776 27770 18788
rect 27801 18785 27813 18788
rect 27847 18785 27859 18819
rect 27801 18779 27859 18785
rect 34054 18776 34060 18828
rect 34112 18816 34118 18828
rect 34425 18819 34483 18825
rect 34425 18816 34437 18819
rect 34112 18788 34437 18816
rect 34112 18776 34118 18788
rect 34425 18785 34437 18788
rect 34471 18785 34483 18819
rect 34425 18779 34483 18785
rect 35894 18776 35900 18828
rect 35952 18816 35958 18828
rect 35952 18788 36216 18816
rect 35952 18776 35958 18788
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18748 19947 18751
rect 19978 18748 19984 18760
rect 19935 18720 19984 18748
rect 19935 18717 19947 18720
rect 19889 18711 19947 18717
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20898 18748 20904 18760
rect 20859 18720 20904 18748
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 23566 18748 23572 18760
rect 23527 18720 23572 18748
rect 23566 18708 23572 18720
rect 23624 18708 23630 18760
rect 23658 18708 23664 18760
rect 23716 18748 23722 18760
rect 25222 18748 25228 18760
rect 23716 18720 23761 18748
rect 25183 18720 25228 18748
rect 23716 18708 23722 18720
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 25317 18751 25375 18757
rect 25317 18717 25329 18751
rect 25363 18748 25375 18751
rect 26142 18748 26148 18760
rect 25363 18720 26148 18748
rect 25363 18717 25375 18720
rect 25317 18711 25375 18717
rect 22462 18640 22468 18692
rect 22520 18680 22526 18692
rect 23109 18683 23167 18689
rect 23109 18680 23121 18683
rect 22520 18652 23121 18680
rect 22520 18640 22526 18652
rect 23109 18649 23121 18652
rect 23155 18649 23167 18683
rect 23676 18680 23704 18708
rect 25332 18680 25360 18711
rect 26142 18708 26148 18720
rect 26200 18708 26206 18760
rect 27614 18708 27620 18760
rect 27672 18748 27678 18760
rect 28077 18751 28135 18757
rect 28077 18748 28089 18751
rect 27672 18720 28089 18748
rect 27672 18708 27678 18720
rect 28077 18717 28089 18720
rect 28123 18717 28135 18751
rect 28077 18711 28135 18717
rect 29273 18751 29331 18757
rect 29273 18717 29285 18751
rect 29319 18717 29331 18751
rect 31018 18748 31024 18760
rect 30979 18720 31024 18748
rect 29273 18711 29331 18717
rect 23676 18652 25360 18680
rect 23109 18643 23167 18649
rect 27890 18640 27896 18692
rect 27948 18680 27954 18692
rect 29288 18680 29316 18711
rect 31018 18708 31024 18720
rect 31076 18708 31082 18760
rect 33778 18708 33784 18760
rect 33836 18748 33842 18760
rect 34609 18751 34667 18757
rect 34609 18748 34621 18751
rect 33836 18720 34621 18748
rect 33836 18708 33842 18720
rect 34609 18717 34621 18720
rect 34655 18748 34667 18751
rect 35437 18751 35495 18757
rect 35437 18748 35449 18751
rect 34655 18720 35449 18748
rect 34655 18717 34667 18720
rect 34609 18711 34667 18717
rect 35437 18717 35449 18720
rect 35483 18748 35495 18751
rect 36078 18748 36084 18760
rect 35483 18720 36084 18748
rect 35483 18717 35495 18720
rect 35437 18711 35495 18717
rect 36078 18708 36084 18720
rect 36136 18708 36142 18760
rect 36188 18757 36216 18788
rect 36173 18751 36231 18757
rect 36173 18717 36185 18751
rect 36219 18717 36231 18751
rect 36173 18711 36231 18717
rect 27948 18652 29316 18680
rect 30377 18683 30435 18689
rect 27948 18640 27954 18652
rect 30377 18649 30389 18683
rect 30423 18680 30435 18683
rect 31202 18680 31208 18692
rect 30423 18652 31208 18680
rect 30423 18649 30435 18652
rect 30377 18643 30435 18649
rect 31202 18640 31208 18652
rect 31260 18640 31266 18692
rect 34057 18683 34115 18689
rect 34057 18649 34069 18683
rect 34103 18680 34115 18683
rect 34422 18680 34428 18692
rect 34103 18652 34428 18680
rect 34103 18649 34115 18652
rect 34057 18643 34115 18649
rect 34422 18640 34428 18652
rect 34480 18640 34486 18692
rect 19242 18612 19248 18624
rect 19203 18584 19248 18612
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 22152 18584 22293 18612
rect 22152 18572 22158 18584
rect 22281 18581 22293 18584
rect 22327 18581 22339 18615
rect 32766 18612 32772 18624
rect 32727 18584 32772 18612
rect 22281 18575 22339 18581
rect 32766 18572 32772 18584
rect 32824 18572 32830 18624
rect 35618 18612 35624 18624
rect 35579 18584 35624 18612
rect 35618 18572 35624 18584
rect 35676 18612 35682 18624
rect 37090 18612 37096 18624
rect 35676 18584 37096 18612
rect 35676 18572 35682 18584
rect 37090 18572 37096 18584
rect 37148 18572 37154 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 19334 18408 19340 18420
rect 19295 18380 19340 18408
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 19610 18408 19616 18420
rect 19571 18380 19616 18408
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 21174 18408 21180 18420
rect 21135 18380 21180 18408
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 22002 18408 22008 18420
rect 21963 18380 22008 18408
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 22278 18368 22284 18420
rect 22336 18408 22342 18420
rect 23201 18411 23259 18417
rect 23201 18408 23213 18411
rect 22336 18380 23213 18408
rect 22336 18368 22342 18380
rect 23201 18377 23213 18380
rect 23247 18408 23259 18411
rect 23566 18408 23572 18420
rect 23247 18380 23572 18408
rect 23247 18377 23259 18380
rect 23201 18371 23259 18377
rect 23566 18368 23572 18380
rect 23624 18368 23630 18420
rect 24857 18411 24915 18417
rect 24857 18377 24869 18411
rect 24903 18408 24915 18411
rect 25222 18408 25228 18420
rect 24903 18380 25228 18408
rect 24903 18377 24915 18380
rect 24857 18371 24915 18377
rect 25222 18368 25228 18380
rect 25280 18408 25286 18420
rect 26234 18408 26240 18420
rect 25280 18380 26240 18408
rect 25280 18368 25286 18380
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 27706 18368 27712 18420
rect 27764 18368 27770 18420
rect 27890 18368 27896 18420
rect 27948 18408 27954 18420
rect 28353 18411 28411 18417
rect 28353 18408 28365 18411
rect 27948 18380 28365 18408
rect 27948 18368 27954 18380
rect 28353 18377 28365 18380
rect 28399 18377 28411 18411
rect 28353 18371 28411 18377
rect 28813 18411 28871 18417
rect 28813 18377 28825 18411
rect 28859 18408 28871 18411
rect 29178 18408 29184 18420
rect 28859 18380 29184 18408
rect 28859 18377 28871 18380
rect 28813 18371 28871 18377
rect 29178 18368 29184 18380
rect 29236 18368 29242 18420
rect 29454 18408 29460 18420
rect 29415 18380 29460 18408
rect 29454 18368 29460 18380
rect 29512 18368 29518 18420
rect 30469 18411 30527 18417
rect 30469 18377 30481 18411
rect 30515 18408 30527 18411
rect 30926 18408 30932 18420
rect 30515 18380 30932 18408
rect 30515 18377 30527 18380
rect 30469 18371 30527 18377
rect 30926 18368 30932 18380
rect 30984 18368 30990 18420
rect 31018 18368 31024 18420
rect 31076 18408 31082 18420
rect 31113 18411 31171 18417
rect 31113 18408 31125 18411
rect 31076 18380 31125 18408
rect 31076 18368 31082 18380
rect 31113 18377 31125 18380
rect 31159 18377 31171 18411
rect 33778 18408 33784 18420
rect 33739 18380 33784 18408
rect 31113 18371 31171 18377
rect 33778 18368 33784 18380
rect 33836 18368 33842 18420
rect 34054 18408 34060 18420
rect 34015 18380 34060 18408
rect 34054 18368 34060 18380
rect 34112 18368 34118 18420
rect 34146 18368 34152 18420
rect 34204 18408 34210 18420
rect 34425 18411 34483 18417
rect 34425 18408 34437 18411
rect 34204 18380 34437 18408
rect 34204 18368 34210 18380
rect 34425 18377 34437 18380
rect 34471 18377 34483 18411
rect 35710 18408 35716 18420
rect 35671 18380 35716 18408
rect 34425 18371 34483 18377
rect 35710 18368 35716 18380
rect 35768 18368 35774 18420
rect 35894 18368 35900 18420
rect 35952 18408 35958 18420
rect 35989 18411 36047 18417
rect 35989 18408 36001 18411
rect 35952 18380 36001 18408
rect 35952 18368 35958 18380
rect 35989 18377 36001 18380
rect 36035 18377 36047 18411
rect 35989 18371 36047 18377
rect 36170 18368 36176 18420
rect 36228 18408 36234 18420
rect 36357 18411 36415 18417
rect 36357 18408 36369 18411
rect 36228 18380 36369 18408
rect 36228 18368 36234 18380
rect 36357 18377 36369 18380
rect 36403 18377 36415 18411
rect 36357 18371 36415 18377
rect 24210 18300 24216 18352
rect 24268 18340 24274 18352
rect 25777 18343 25835 18349
rect 25777 18340 25789 18343
rect 24268 18312 25789 18340
rect 24268 18300 24274 18312
rect 25777 18309 25789 18312
rect 25823 18340 25835 18343
rect 26510 18340 26516 18352
rect 25823 18312 26516 18340
rect 25823 18309 25835 18312
rect 25777 18303 25835 18309
rect 26510 18300 26516 18312
rect 26568 18300 26574 18352
rect 27724 18340 27752 18368
rect 27985 18343 28043 18349
rect 27985 18340 27997 18343
rect 27724 18312 27997 18340
rect 27985 18309 27997 18312
rect 28031 18309 28043 18343
rect 27985 18303 28043 18309
rect 29917 18343 29975 18349
rect 29917 18309 29929 18343
rect 29963 18340 29975 18343
rect 31036 18340 31064 18368
rect 29963 18312 31064 18340
rect 29963 18309 29975 18312
rect 29917 18303 29975 18309
rect 21913 18275 21971 18281
rect 21913 18241 21925 18275
rect 21959 18272 21971 18275
rect 22462 18272 22468 18284
rect 21959 18244 22468 18272
rect 21959 18241 21971 18244
rect 21913 18235 21971 18241
rect 22462 18232 22468 18244
rect 22520 18232 22526 18284
rect 22554 18232 22560 18284
rect 22612 18272 22618 18284
rect 27709 18275 27767 18281
rect 22612 18244 22657 18272
rect 22612 18232 22618 18244
rect 27709 18241 27721 18275
rect 27755 18272 27767 18275
rect 28626 18272 28632 18284
rect 27755 18244 28632 18272
rect 27755 18241 27767 18244
rect 27709 18235 27767 18241
rect 28626 18232 28632 18244
rect 28684 18232 28690 18284
rect 30466 18232 30472 18284
rect 30524 18272 30530 18284
rect 30745 18275 30803 18281
rect 30745 18272 30757 18275
rect 30524 18244 30757 18272
rect 30524 18232 30530 18244
rect 30745 18241 30757 18244
rect 30791 18241 30803 18275
rect 30745 18235 30803 18241
rect 32217 18275 32275 18281
rect 32217 18241 32229 18275
rect 32263 18272 32275 18275
rect 32398 18272 32404 18284
rect 32263 18244 32404 18272
rect 32263 18241 32275 18244
rect 32217 18235 32275 18241
rect 32398 18232 32404 18244
rect 32456 18272 32462 18284
rect 33229 18275 33287 18281
rect 33229 18272 33241 18275
rect 32456 18244 33241 18272
rect 32456 18232 32462 18244
rect 33229 18241 33241 18244
rect 33275 18241 33287 18275
rect 33229 18235 33287 18241
rect 19797 18207 19855 18213
rect 19797 18173 19809 18207
rect 19843 18204 19855 18207
rect 19886 18204 19892 18216
rect 19843 18176 19892 18204
rect 19843 18173 19855 18176
rect 19797 18167 19855 18173
rect 19886 18164 19892 18176
rect 19944 18164 19950 18216
rect 22370 18204 22376 18216
rect 22331 18176 22376 18204
rect 22370 18164 22376 18176
rect 22428 18164 22434 18216
rect 23842 18204 23848 18216
rect 23803 18176 23848 18204
rect 23842 18164 23848 18176
rect 23900 18164 23906 18216
rect 25682 18164 25688 18216
rect 25740 18204 25746 18216
rect 25961 18207 26019 18213
rect 25961 18204 25973 18207
rect 25740 18176 25973 18204
rect 25740 18164 25746 18176
rect 25961 18173 25973 18176
rect 26007 18173 26019 18207
rect 25961 18167 26019 18173
rect 32766 18164 32772 18216
rect 32824 18204 32830 18216
rect 33045 18207 33103 18213
rect 33045 18204 33057 18207
rect 32824 18176 33057 18204
rect 32824 18164 32830 18176
rect 33045 18173 33057 18176
rect 33091 18173 33103 18207
rect 33045 18167 33103 18173
rect 20070 18145 20076 18148
rect 18969 18139 19027 18145
rect 18969 18105 18981 18139
rect 19015 18136 19027 18139
rect 20064 18136 20076 18145
rect 19015 18108 20076 18136
rect 19015 18105 19027 18108
rect 18969 18099 19027 18105
rect 20064 18099 20076 18108
rect 20070 18096 20076 18099
rect 20128 18096 20134 18148
rect 23658 18096 23664 18148
rect 23716 18136 23722 18148
rect 24394 18136 24400 18148
rect 23716 18108 24400 18136
rect 23716 18096 23722 18108
rect 24394 18096 24400 18108
rect 24452 18096 24458 18148
rect 32585 18139 32643 18145
rect 32585 18105 32597 18139
rect 32631 18136 32643 18139
rect 33137 18139 33195 18145
rect 33137 18136 33149 18139
rect 32631 18108 33149 18136
rect 32631 18105 32643 18108
rect 32585 18099 32643 18105
rect 33137 18105 33149 18108
rect 33183 18136 33195 18139
rect 33410 18136 33416 18148
rect 33183 18108 33416 18136
rect 33183 18105 33195 18108
rect 33137 18099 33195 18105
rect 33410 18096 33416 18108
rect 33468 18096 33474 18148
rect 34146 18096 34152 18148
rect 34204 18136 34210 18148
rect 34698 18136 34704 18148
rect 34204 18108 34704 18136
rect 34204 18096 34210 18108
rect 34698 18096 34704 18108
rect 34756 18096 34762 18148
rect 18598 18068 18604 18080
rect 18559 18040 18604 18068
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 21542 18068 21548 18080
rect 21503 18040 21548 18068
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 25222 18068 25228 18080
rect 25183 18040 25228 18068
rect 25222 18028 25228 18040
rect 25280 18028 25286 18080
rect 32674 18068 32680 18080
rect 32635 18040 32680 18068
rect 32674 18028 32680 18040
rect 32732 18028 32738 18080
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 22278 17864 22284 17876
rect 22239 17836 22284 17864
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 22370 17824 22376 17876
rect 22428 17864 22434 17876
rect 22557 17867 22615 17873
rect 22557 17864 22569 17867
rect 22428 17836 22569 17864
rect 22428 17824 22434 17836
rect 22557 17833 22569 17836
rect 22603 17833 22615 17867
rect 22557 17827 22615 17833
rect 23293 17867 23351 17873
rect 23293 17833 23305 17867
rect 23339 17864 23351 17867
rect 23382 17864 23388 17876
rect 23339 17836 23388 17864
rect 23339 17833 23351 17836
rect 23293 17827 23351 17833
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 23658 17864 23664 17876
rect 23619 17836 23664 17864
rect 23658 17824 23664 17836
rect 23716 17824 23722 17876
rect 27890 17864 27896 17876
rect 27851 17836 27896 17864
rect 27890 17824 27896 17836
rect 27948 17824 27954 17876
rect 34238 17824 34244 17876
rect 34296 17864 34302 17876
rect 34793 17867 34851 17873
rect 34793 17864 34805 17867
rect 34296 17836 34805 17864
rect 34296 17824 34302 17836
rect 34793 17833 34805 17836
rect 34839 17833 34851 17867
rect 34793 17827 34851 17833
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 19613 17799 19671 17805
rect 19613 17796 19625 17799
rect 19024 17768 19625 17796
rect 19024 17756 19030 17768
rect 19613 17765 19625 17768
rect 19659 17796 19671 17799
rect 21168 17799 21226 17805
rect 21168 17796 21180 17799
rect 19659 17768 21180 17796
rect 19659 17765 19671 17768
rect 19613 17759 19671 17765
rect 21168 17765 21180 17768
rect 21214 17796 21226 17799
rect 21358 17796 21364 17808
rect 21214 17768 21364 17796
rect 21214 17765 21226 17768
rect 21168 17759 21226 17765
rect 21358 17756 21364 17768
rect 21416 17756 21422 17808
rect 24489 17799 24547 17805
rect 24489 17765 24501 17799
rect 24535 17796 24547 17799
rect 24848 17799 24906 17805
rect 24848 17796 24860 17799
rect 24535 17768 24860 17796
rect 24535 17765 24547 17768
rect 24489 17759 24547 17765
rect 24848 17765 24860 17768
rect 24894 17796 24906 17799
rect 25222 17796 25228 17808
rect 24894 17768 25228 17796
rect 24894 17765 24906 17768
rect 24848 17759 24906 17765
rect 25222 17756 25228 17768
rect 25280 17756 25286 17808
rect 26234 17756 26240 17808
rect 26292 17796 26298 17808
rect 26694 17796 26700 17808
rect 26292 17768 26700 17796
rect 26292 17756 26298 17768
rect 26694 17756 26700 17768
rect 26752 17805 26758 17808
rect 26752 17799 26816 17805
rect 26752 17765 26770 17799
rect 26804 17765 26816 17799
rect 26752 17759 26816 17765
rect 26752 17756 26758 17759
rect 22554 17688 22560 17740
rect 22612 17728 22618 17740
rect 22925 17731 22983 17737
rect 22925 17728 22937 17731
rect 22612 17700 22937 17728
rect 22612 17688 22618 17700
rect 22925 17697 22937 17700
rect 22971 17697 22983 17731
rect 23106 17728 23112 17740
rect 23067 17700 23112 17728
rect 22925 17691 22983 17697
rect 23106 17688 23112 17700
rect 23164 17688 23170 17740
rect 24302 17688 24308 17740
rect 24360 17728 24366 17740
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 24360 17700 24593 17728
rect 24360 17688 24366 17700
rect 24581 17697 24593 17700
rect 24627 17728 24639 17731
rect 26513 17731 26571 17737
rect 26513 17728 26525 17731
rect 24627 17700 26525 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 26513 17697 26525 17700
rect 26559 17728 26571 17731
rect 27062 17728 27068 17740
rect 26559 17700 27068 17728
rect 26559 17697 26571 17700
rect 26513 17691 26571 17697
rect 27062 17688 27068 17700
rect 27120 17688 27126 17740
rect 32490 17728 32496 17740
rect 32451 17700 32496 17728
rect 32490 17688 32496 17700
rect 32548 17688 32554 17740
rect 32585 17731 32643 17737
rect 32585 17697 32597 17731
rect 32631 17728 32643 17731
rect 32858 17728 32864 17740
rect 32631 17700 32864 17728
rect 32631 17697 32643 17700
rect 32585 17691 32643 17697
rect 32858 17688 32864 17700
rect 32916 17688 32922 17740
rect 33318 17688 33324 17740
rect 33376 17728 33382 17740
rect 34701 17731 34759 17737
rect 34701 17728 34713 17731
rect 33376 17700 34713 17728
rect 33376 17688 33382 17700
rect 34701 17697 34713 17700
rect 34747 17697 34759 17731
rect 34701 17691 34759 17697
rect 35897 17731 35955 17737
rect 35897 17697 35909 17731
rect 35943 17728 35955 17731
rect 36538 17728 36544 17740
rect 35943 17700 36544 17728
rect 35943 17697 35955 17700
rect 35897 17691 35955 17697
rect 36538 17688 36544 17700
rect 36596 17688 36602 17740
rect 19610 17620 19616 17672
rect 19668 17660 19674 17672
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19668 17632 19717 17660
rect 19668 17620 19674 17632
rect 19705 17629 19717 17632
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 19978 17660 19984 17672
rect 19935 17632 19984 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20898 17660 20904 17672
rect 20640 17632 20904 17660
rect 19242 17524 19248 17536
rect 19203 17496 19248 17524
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 19886 17484 19892 17536
rect 19944 17524 19950 17536
rect 20640 17533 20668 17632
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 30285 17663 30343 17669
rect 30285 17629 30297 17663
rect 30331 17660 30343 17663
rect 30374 17660 30380 17672
rect 30331 17632 30380 17660
rect 30331 17629 30343 17632
rect 30285 17623 30343 17629
rect 30374 17620 30380 17632
rect 30432 17620 30438 17672
rect 32674 17620 32680 17672
rect 32732 17660 32738 17672
rect 32732 17632 32777 17660
rect 32732 17620 32738 17632
rect 34882 17620 34888 17672
rect 34940 17660 34946 17672
rect 34940 17632 34985 17660
rect 34940 17620 34946 17632
rect 29365 17595 29423 17601
rect 29365 17561 29377 17595
rect 29411 17592 29423 17595
rect 29914 17592 29920 17604
rect 29411 17564 29920 17592
rect 29411 17561 29423 17564
rect 29365 17555 29423 17561
rect 29914 17552 29920 17564
rect 29972 17552 29978 17604
rect 20257 17527 20315 17533
rect 20257 17524 20269 17527
rect 19944 17496 20269 17524
rect 19944 17484 19950 17496
rect 20257 17493 20269 17496
rect 20303 17524 20315 17527
rect 20625 17527 20683 17533
rect 20625 17524 20637 17527
rect 20303 17496 20637 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 20625 17493 20637 17496
rect 20671 17493 20683 17527
rect 20625 17487 20683 17493
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 24912 17496 25973 17524
rect 24912 17484 24918 17496
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 29730 17524 29736 17536
rect 29691 17496 29736 17524
rect 25961 17487 26019 17493
rect 29730 17484 29736 17496
rect 29788 17484 29794 17536
rect 31662 17524 31668 17536
rect 31623 17496 31668 17524
rect 31662 17484 31668 17496
rect 31720 17484 31726 17536
rect 32122 17524 32128 17536
rect 32083 17496 32128 17524
rect 32122 17484 32128 17496
rect 32180 17484 32186 17536
rect 34330 17524 34336 17536
rect 34291 17496 34336 17524
rect 34330 17484 34336 17496
rect 34388 17484 34394 17536
rect 35342 17484 35348 17536
rect 35400 17524 35406 17536
rect 35529 17527 35587 17533
rect 35529 17524 35541 17527
rect 35400 17496 35541 17524
rect 35400 17484 35406 17496
rect 35529 17493 35541 17496
rect 35575 17524 35587 17527
rect 35986 17524 35992 17536
rect 35575 17496 35992 17524
rect 35575 17493 35587 17496
rect 35529 17487 35587 17493
rect 35986 17484 35992 17496
rect 36044 17484 36050 17536
rect 36078 17484 36084 17536
rect 36136 17524 36142 17536
rect 36136 17496 36181 17524
rect 36136 17484 36142 17496
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 18966 17320 18972 17332
rect 18927 17292 18972 17320
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 21082 17320 21088 17332
rect 21043 17292 21088 17320
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 25222 17320 25228 17332
rect 25183 17292 25228 17320
rect 25222 17280 25228 17292
rect 25280 17280 25286 17332
rect 26694 17320 26700 17332
rect 26655 17292 26700 17320
rect 26694 17280 26700 17292
rect 26752 17320 26758 17332
rect 26973 17323 27031 17329
rect 26973 17320 26985 17323
rect 26752 17292 26985 17320
rect 26752 17280 26758 17292
rect 26973 17289 26985 17292
rect 27019 17289 27031 17323
rect 28718 17320 28724 17332
rect 28679 17292 28724 17320
rect 26973 17283 27031 17289
rect 28718 17280 28724 17292
rect 28776 17280 28782 17332
rect 34238 17280 34244 17332
rect 34296 17320 34302 17332
rect 34333 17323 34391 17329
rect 34333 17320 34345 17323
rect 34296 17292 34345 17320
rect 34296 17280 34302 17292
rect 34333 17289 34345 17292
rect 34379 17289 34391 17323
rect 34333 17283 34391 17289
rect 34606 17280 34612 17332
rect 34664 17280 34670 17332
rect 36538 17320 36544 17332
rect 36499 17292 36544 17320
rect 36538 17280 36544 17292
rect 36596 17280 36602 17332
rect 21913 17255 21971 17261
rect 21913 17221 21925 17255
rect 21959 17252 21971 17255
rect 23106 17252 23112 17264
rect 21959 17224 23112 17252
rect 21959 17221 21971 17224
rect 21913 17215 21971 17221
rect 23106 17212 23112 17224
rect 23164 17212 23170 17264
rect 29273 17255 29331 17261
rect 29273 17221 29285 17255
rect 29319 17252 29331 17255
rect 30466 17252 30472 17264
rect 29319 17224 30472 17252
rect 29319 17221 29331 17224
rect 29273 17215 29331 17221
rect 30466 17212 30472 17224
rect 30524 17212 30530 17264
rect 34624 17252 34652 17280
rect 35158 17252 35164 17264
rect 34624 17224 35164 17252
rect 35158 17212 35164 17224
rect 35216 17212 35222 17264
rect 22554 17184 22560 17196
rect 22515 17156 22560 17184
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 29730 17144 29736 17196
rect 29788 17184 29794 17196
rect 29825 17187 29883 17193
rect 29825 17184 29837 17187
rect 29788 17156 29837 17184
rect 29788 17144 29794 17156
rect 29825 17153 29837 17156
rect 29871 17153 29883 17187
rect 29825 17147 29883 17153
rect 34330 17144 34336 17196
rect 34388 17184 34394 17196
rect 35897 17187 35955 17193
rect 35897 17184 35909 17187
rect 34388 17156 35909 17184
rect 34388 17144 34394 17156
rect 35897 17153 35909 17156
rect 35943 17153 35955 17187
rect 35897 17147 35955 17153
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 19972 17119 20030 17125
rect 19751 17088 19932 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 19904 17060 19932 17088
rect 19972 17085 19984 17119
rect 20018 17116 20030 17119
rect 20346 17116 20352 17128
rect 20018 17088 20352 17116
rect 20018 17085 20030 17088
rect 19972 17079 20030 17085
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 22278 17116 22284 17128
rect 22239 17088 22284 17116
rect 22278 17076 22284 17088
rect 22336 17116 22342 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22336 17088 22937 17116
rect 22336 17076 22342 17088
rect 22925 17085 22937 17088
rect 22971 17085 22983 17119
rect 23842 17116 23848 17128
rect 23803 17088 23848 17116
rect 22925 17079 22983 17085
rect 23842 17076 23848 17088
rect 23900 17076 23906 17128
rect 25317 17119 25375 17125
rect 25317 17085 25329 17119
rect 25363 17116 25375 17119
rect 25958 17116 25964 17128
rect 25363 17088 25964 17116
rect 25363 17085 25375 17088
rect 25317 17079 25375 17085
rect 25958 17076 25964 17088
rect 26016 17076 26022 17128
rect 27893 17119 27951 17125
rect 27893 17085 27905 17119
rect 27939 17116 27951 17119
rect 28166 17116 28172 17128
rect 27939 17088 28172 17116
rect 27939 17085 27951 17088
rect 27893 17079 27951 17085
rect 28166 17076 28172 17088
rect 28224 17076 28230 17128
rect 28353 17119 28411 17125
rect 28353 17085 28365 17119
rect 28399 17116 28411 17119
rect 28902 17116 28908 17128
rect 28399 17088 28908 17116
rect 28399 17085 28411 17088
rect 28353 17079 28411 17085
rect 28902 17076 28908 17088
rect 28960 17076 28966 17128
rect 31573 17119 31631 17125
rect 31573 17116 31585 17119
rect 31128 17088 31585 17116
rect 19610 17008 19616 17060
rect 19668 17008 19674 17060
rect 19886 17008 19892 17060
rect 19944 17008 19950 17060
rect 21726 17048 21732 17060
rect 21687 17020 21732 17048
rect 21726 17008 21732 17020
rect 21784 17048 21790 17060
rect 22373 17051 22431 17057
rect 22373 17048 22385 17051
rect 21784 17020 22385 17048
rect 21784 17008 21790 17020
rect 22373 17017 22385 17020
rect 22419 17017 22431 17051
rect 22373 17011 22431 17017
rect 23477 17051 23535 17057
rect 23477 17017 23489 17051
rect 23523 17048 23535 17051
rect 24112 17051 24170 17057
rect 24112 17048 24124 17051
rect 23523 17020 24124 17048
rect 23523 17017 23535 17020
rect 23477 17011 23535 17017
rect 24112 17017 24124 17020
rect 24158 17048 24170 17051
rect 24854 17048 24860 17060
rect 24158 17020 24860 17048
rect 24158 17017 24170 17020
rect 24112 17011 24170 17017
rect 24854 17008 24860 17020
rect 24912 17008 24918 17060
rect 25498 17008 25504 17060
rect 25556 17057 25562 17060
rect 25556 17051 25620 17057
rect 25556 17017 25574 17051
rect 25608 17017 25620 17051
rect 25556 17011 25620 17017
rect 27985 17051 28043 17057
rect 27985 17017 27997 17051
rect 28031 17048 28043 17051
rect 28718 17048 28724 17060
rect 28031 17020 28724 17048
rect 28031 17017 28043 17020
rect 27985 17011 28043 17017
rect 25556 17008 25562 17011
rect 28718 17008 28724 17020
rect 28776 17008 28782 17060
rect 29641 17051 29699 17057
rect 29641 17048 29653 17051
rect 29012 17020 29653 17048
rect 18598 16980 18604 16992
rect 18559 16952 18604 16980
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 19337 16983 19395 16989
rect 19337 16949 19349 16983
rect 19383 16980 19395 16983
rect 19628 16980 19656 17008
rect 29012 16992 29040 17020
rect 29641 17017 29653 17020
rect 29687 17017 29699 17051
rect 29641 17011 29699 17017
rect 31128 16992 31156 17088
rect 31573 17085 31585 17088
rect 31619 17085 31631 17119
rect 35912 17116 35940 17147
rect 35986 17144 35992 17196
rect 36044 17184 36050 17196
rect 36044 17156 36089 17184
rect 36044 17144 36050 17156
rect 36817 17119 36875 17125
rect 36817 17116 36829 17119
rect 35912 17088 36829 17116
rect 31573 17079 31631 17085
rect 36817 17085 36829 17088
rect 36863 17085 36875 17119
rect 36817 17079 36875 17085
rect 31386 17048 31392 17060
rect 31347 17020 31392 17048
rect 31386 17008 31392 17020
rect 31444 17008 31450 17060
rect 31662 17008 31668 17060
rect 31720 17048 31726 17060
rect 31846 17057 31852 17060
rect 31840 17048 31852 17057
rect 31720 17020 31852 17048
rect 31720 17008 31726 17020
rect 31840 17011 31852 17020
rect 31846 17008 31852 17011
rect 31904 17008 31910 17060
rect 32858 17008 32864 17060
rect 32916 17048 32922 17060
rect 33229 17051 33287 17057
rect 33229 17048 33241 17051
rect 32916 17020 33241 17048
rect 32916 17008 32922 17020
rect 33229 17017 33241 17020
rect 33275 17017 33287 17051
rect 33229 17011 33287 17017
rect 33781 17051 33839 17057
rect 33781 17017 33793 17051
rect 33827 17048 33839 17051
rect 34422 17048 34428 17060
rect 33827 17020 34428 17048
rect 33827 17017 33839 17020
rect 33781 17011 33839 17017
rect 34422 17008 34428 17020
rect 34480 17008 34486 17060
rect 35345 17051 35403 17057
rect 35345 17017 35357 17051
rect 35391 17048 35403 17051
rect 35391 17020 35848 17048
rect 35391 17017 35403 17020
rect 35345 17011 35403 17017
rect 20254 16980 20260 16992
rect 19383 16952 20260 16980
rect 19383 16949 19395 16952
rect 19337 16943 19395 16949
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 21358 16980 21364 16992
rect 21319 16952 21364 16980
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 27062 16940 27068 16992
rect 27120 16980 27126 16992
rect 27341 16983 27399 16989
rect 27341 16980 27353 16983
rect 27120 16952 27353 16980
rect 27120 16940 27126 16952
rect 27341 16949 27353 16952
rect 27387 16949 27399 16983
rect 28994 16980 29000 16992
rect 28955 16952 29000 16980
rect 27341 16943 27399 16949
rect 28994 16940 29000 16952
rect 29052 16940 29058 16992
rect 29733 16983 29791 16989
rect 29733 16949 29745 16983
rect 29779 16980 29791 16983
rect 29914 16980 29920 16992
rect 29779 16952 29920 16980
rect 29779 16949 29791 16952
rect 29733 16943 29791 16949
rect 29914 16940 29920 16952
rect 29972 16940 29978 16992
rect 31110 16980 31116 16992
rect 31071 16952 31116 16980
rect 31110 16940 31116 16952
rect 31168 16940 31174 16992
rect 31404 16980 31432 17008
rect 32674 16980 32680 16992
rect 31404 16952 32680 16980
rect 32674 16940 32680 16952
rect 32732 16980 32738 16992
rect 32953 16983 33011 16989
rect 32953 16980 32965 16983
rect 32732 16952 32965 16980
rect 32732 16940 32738 16952
rect 32953 16949 32965 16952
rect 32999 16949 33011 16983
rect 32953 16943 33011 16949
rect 33318 16940 33324 16992
rect 33376 16980 33382 16992
rect 33597 16983 33655 16989
rect 33597 16980 33609 16983
rect 33376 16952 33609 16980
rect 33376 16940 33382 16952
rect 33597 16949 33609 16952
rect 33643 16949 33655 16983
rect 35434 16980 35440 16992
rect 35395 16952 35440 16980
rect 33597 16943 33655 16949
rect 35434 16940 35440 16952
rect 35492 16940 35498 16992
rect 35820 16989 35848 17020
rect 35805 16983 35863 16989
rect 35805 16949 35817 16983
rect 35851 16980 35863 16983
rect 35894 16980 35900 16992
rect 35851 16952 35900 16980
rect 35851 16949 35863 16952
rect 35805 16943 35863 16949
rect 35894 16940 35900 16952
rect 35952 16940 35958 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 22278 16776 22284 16788
rect 22239 16748 22284 16776
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 22554 16776 22560 16788
rect 22515 16748 22560 16776
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 23106 16776 23112 16788
rect 23067 16748 23112 16776
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 23842 16736 23848 16788
rect 23900 16776 23906 16788
rect 23937 16779 23995 16785
rect 23937 16776 23949 16779
rect 23900 16748 23949 16776
rect 23900 16736 23906 16748
rect 23937 16745 23949 16748
rect 23983 16776 23995 16779
rect 24302 16776 24308 16788
rect 23983 16748 24308 16776
rect 23983 16745 23995 16748
rect 23937 16739 23995 16745
rect 24302 16736 24308 16748
rect 24360 16736 24366 16788
rect 24397 16779 24455 16785
rect 24397 16745 24409 16779
rect 24443 16776 24455 16779
rect 24486 16776 24492 16788
rect 24443 16748 24492 16776
rect 24443 16745 24455 16748
rect 24397 16739 24455 16745
rect 24486 16736 24492 16748
rect 24544 16736 24550 16788
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25498 16776 25504 16788
rect 25459 16748 25504 16776
rect 25498 16736 25504 16748
rect 25556 16736 25562 16788
rect 25869 16779 25927 16785
rect 25869 16745 25881 16779
rect 25915 16776 25927 16779
rect 25958 16776 25964 16788
rect 25915 16748 25964 16776
rect 25915 16745 25927 16748
rect 25869 16739 25927 16745
rect 25958 16736 25964 16748
rect 26016 16776 26022 16788
rect 27062 16776 27068 16788
rect 26016 16748 27068 16776
rect 26016 16736 26022 16748
rect 27062 16736 27068 16748
rect 27120 16736 27126 16788
rect 27430 16776 27436 16788
rect 27391 16748 27436 16776
rect 27430 16736 27436 16748
rect 27488 16736 27494 16788
rect 29730 16776 29736 16788
rect 29691 16748 29736 16776
rect 29730 16736 29736 16748
rect 29788 16736 29794 16788
rect 31941 16779 31999 16785
rect 31941 16745 31953 16779
rect 31987 16776 31999 16779
rect 32122 16776 32128 16788
rect 31987 16748 32128 16776
rect 31987 16745 31999 16748
rect 31941 16739 31999 16745
rect 32122 16736 32128 16748
rect 32180 16736 32186 16788
rect 32401 16779 32459 16785
rect 32401 16745 32413 16779
rect 32447 16776 32459 16779
rect 32490 16776 32496 16788
rect 32447 16748 32496 16776
rect 32447 16745 32459 16748
rect 32401 16739 32459 16745
rect 32490 16736 32496 16748
rect 32548 16776 32554 16788
rect 33042 16776 33048 16788
rect 32548 16748 33048 16776
rect 32548 16736 32554 16748
rect 33042 16736 33048 16748
rect 33100 16736 33106 16788
rect 33134 16736 33140 16788
rect 33192 16776 33198 16788
rect 33235 16779 33293 16785
rect 33235 16776 33247 16779
rect 33192 16748 33247 16776
rect 33192 16736 33198 16748
rect 33235 16745 33247 16748
rect 33281 16745 33293 16779
rect 33235 16739 33293 16745
rect 34238 16736 34244 16788
rect 34296 16776 34302 16788
rect 34609 16779 34667 16785
rect 34609 16776 34621 16779
rect 34296 16748 34621 16776
rect 34296 16736 34302 16748
rect 34609 16745 34621 16748
rect 34655 16745 34667 16779
rect 34609 16739 34667 16745
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 34885 16779 34943 16785
rect 34885 16776 34897 16779
rect 34848 16748 34897 16776
rect 34848 16736 34854 16748
rect 34885 16745 34897 16748
rect 34931 16745 34943 16779
rect 34885 16739 34943 16745
rect 19153 16711 19211 16717
rect 19153 16677 19165 16711
rect 19199 16708 19211 16711
rect 19886 16708 19892 16720
rect 19199 16680 19892 16708
rect 19199 16677 19211 16680
rect 19153 16671 19211 16677
rect 19886 16668 19892 16680
rect 19944 16668 19950 16720
rect 24765 16711 24823 16717
rect 24765 16677 24777 16711
rect 24811 16708 24823 16711
rect 25222 16708 25228 16720
rect 24811 16680 25228 16708
rect 24811 16677 24823 16680
rect 24765 16671 24823 16677
rect 25222 16668 25228 16680
rect 25280 16668 25286 16720
rect 28166 16668 28172 16720
rect 28224 16708 28230 16720
rect 28598 16711 28656 16717
rect 28598 16708 28610 16711
rect 28224 16680 28610 16708
rect 28224 16668 28230 16680
rect 28598 16677 28610 16680
rect 28644 16677 28656 16711
rect 34900 16708 34928 16739
rect 35986 16736 35992 16788
rect 36044 16776 36050 16788
rect 36817 16779 36875 16785
rect 36817 16776 36829 16779
rect 36044 16748 36829 16776
rect 36044 16736 36050 16748
rect 36817 16745 36829 16748
rect 36863 16745 36875 16779
rect 36817 16739 36875 16745
rect 35710 16717 35716 16720
rect 35682 16711 35716 16717
rect 35682 16708 35694 16711
rect 34900 16680 35694 16708
rect 28598 16671 28656 16677
rect 35682 16677 35694 16680
rect 35768 16708 35774 16720
rect 35768 16680 35830 16708
rect 35682 16671 35716 16677
rect 35710 16668 35716 16671
rect 35768 16668 35774 16680
rect 19610 16640 19616 16652
rect 19523 16612 19616 16640
rect 19610 16600 19616 16612
rect 19668 16640 19674 16652
rect 21168 16643 21226 16649
rect 21168 16640 21180 16643
rect 19668 16612 21180 16640
rect 19668 16600 19674 16612
rect 21168 16609 21180 16612
rect 21214 16640 21226 16643
rect 21726 16640 21732 16652
rect 21214 16612 21732 16640
rect 21214 16609 21226 16612
rect 21168 16603 21226 16609
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 27249 16643 27307 16649
rect 27249 16609 27261 16643
rect 27295 16640 27307 16643
rect 27522 16640 27528 16652
rect 27295 16612 27528 16640
rect 27295 16609 27307 16612
rect 27249 16603 27307 16609
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 28353 16643 28411 16649
rect 28353 16609 28365 16643
rect 28399 16640 28411 16643
rect 28994 16640 29000 16652
rect 28399 16612 29000 16640
rect 28399 16609 28411 16612
rect 28353 16603 28411 16609
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 30558 16640 30564 16652
rect 30471 16612 30564 16640
rect 30558 16600 30564 16612
rect 30616 16640 30622 16652
rect 31113 16643 31171 16649
rect 31113 16640 31125 16643
rect 30616 16612 31125 16640
rect 30616 16600 30622 16612
rect 31113 16609 31125 16612
rect 31159 16609 31171 16643
rect 31113 16603 31171 16609
rect 32030 16600 32036 16652
rect 32088 16640 32094 16652
rect 32769 16643 32827 16649
rect 32769 16640 32781 16643
rect 32088 16612 32781 16640
rect 32088 16600 32094 16612
rect 32769 16609 32781 16612
rect 32815 16640 32827 16643
rect 33134 16640 33140 16652
rect 32815 16612 33140 16640
rect 32815 16609 32827 16612
rect 32769 16603 32827 16609
rect 33134 16600 33140 16612
rect 33192 16600 33198 16652
rect 33410 16600 33416 16652
rect 33468 16640 33474 16652
rect 33505 16643 33563 16649
rect 33505 16640 33517 16643
rect 33468 16612 33517 16640
rect 33468 16600 33474 16612
rect 33505 16609 33517 16612
rect 33551 16609 33563 16643
rect 33505 16603 33563 16609
rect 35250 16600 35256 16652
rect 35308 16640 35314 16652
rect 35986 16640 35992 16652
rect 35308 16612 35992 16640
rect 35308 16600 35314 16612
rect 35986 16600 35992 16612
rect 36044 16600 36050 16652
rect 19334 16532 19340 16584
rect 19392 16572 19398 16584
rect 19705 16575 19763 16581
rect 19705 16572 19717 16575
rect 19392 16544 19717 16572
rect 19392 16532 19398 16544
rect 19705 16541 19717 16544
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16572 19947 16575
rect 19978 16572 19984 16584
rect 19935 16544 19984 16572
rect 19935 16541 19947 16544
rect 19889 16535 19947 16541
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20824 16544 20913 16572
rect 20824 16448 20852 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 24394 16532 24400 16584
rect 24452 16572 24458 16584
rect 24949 16575 25007 16581
rect 24949 16572 24961 16575
rect 24452 16544 24961 16572
rect 24452 16532 24458 16544
rect 24949 16541 24961 16544
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 33226 16532 33232 16584
rect 33284 16572 33290 16584
rect 35437 16575 35495 16581
rect 33284 16544 33329 16572
rect 33284 16532 33290 16544
rect 35437 16541 35449 16575
rect 35483 16541 35495 16575
rect 35437 16535 35495 16541
rect 35452 16448 35480 16535
rect 20717 16439 20775 16445
rect 20717 16405 20729 16439
rect 20763 16436 20775 16439
rect 20806 16436 20812 16448
rect 20763 16408 20812 16436
rect 20763 16405 20775 16408
rect 20717 16399 20775 16405
rect 20806 16396 20812 16408
rect 20864 16396 20870 16448
rect 30745 16439 30803 16445
rect 30745 16405 30757 16439
rect 30791 16436 30803 16439
rect 33226 16436 33232 16448
rect 30791 16408 33232 16436
rect 30791 16405 30803 16408
rect 30745 16399 30803 16405
rect 33226 16396 33232 16408
rect 33284 16396 33290 16448
rect 35345 16439 35403 16445
rect 35345 16405 35357 16439
rect 35391 16436 35403 16439
rect 35434 16436 35440 16448
rect 35391 16408 35440 16436
rect 35391 16405 35403 16408
rect 35345 16399 35403 16405
rect 35434 16396 35440 16408
rect 35492 16396 35498 16448
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 19334 16232 19340 16244
rect 19295 16204 19340 16232
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 19610 16232 19616 16244
rect 19571 16204 19616 16232
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 21358 16232 21364 16244
rect 21319 16204 21364 16232
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 24121 16235 24179 16241
rect 24121 16201 24133 16235
rect 24167 16232 24179 16235
rect 24213 16235 24271 16241
rect 24213 16232 24225 16235
rect 24167 16204 24225 16232
rect 24167 16201 24179 16204
rect 24121 16195 24179 16201
rect 24213 16201 24225 16204
rect 24259 16232 24271 16235
rect 24394 16232 24400 16244
rect 24259 16204 24400 16232
rect 24259 16201 24271 16204
rect 24213 16195 24271 16201
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 24489 16235 24547 16241
rect 24489 16201 24501 16235
rect 24535 16232 24547 16235
rect 24762 16232 24768 16244
rect 24535 16204 24768 16232
rect 24535 16201 24547 16204
rect 24489 16195 24547 16201
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 25222 16232 25228 16244
rect 25183 16204 25228 16232
rect 25222 16192 25228 16204
rect 25280 16192 25286 16244
rect 28166 16192 28172 16244
rect 28224 16232 28230 16244
rect 28353 16235 28411 16241
rect 28353 16232 28365 16235
rect 28224 16204 28365 16232
rect 28224 16192 28230 16204
rect 28353 16201 28365 16204
rect 28399 16232 28411 16235
rect 28629 16235 28687 16241
rect 28629 16232 28641 16235
rect 28399 16204 28641 16232
rect 28399 16201 28411 16204
rect 28353 16195 28411 16201
rect 28629 16201 28641 16204
rect 28675 16201 28687 16235
rect 28629 16195 28687 16201
rect 31941 16235 31999 16241
rect 31941 16201 31953 16235
rect 31987 16232 31999 16235
rect 32490 16232 32496 16244
rect 31987 16204 32496 16232
rect 31987 16201 31999 16204
rect 31941 16195 31999 16201
rect 32490 16192 32496 16204
rect 32548 16232 32554 16244
rect 32950 16232 32956 16244
rect 32548 16204 32956 16232
rect 32548 16192 32554 16204
rect 32950 16192 32956 16204
rect 33008 16192 33014 16244
rect 33410 16192 33416 16244
rect 33468 16232 33474 16244
rect 33873 16235 33931 16241
rect 33873 16232 33885 16235
rect 33468 16204 33885 16232
rect 33468 16192 33474 16204
rect 33873 16201 33885 16204
rect 33919 16232 33931 16235
rect 34517 16235 34575 16241
rect 34517 16232 34529 16235
rect 33919 16204 34529 16232
rect 33919 16201 33931 16204
rect 33873 16195 33931 16201
rect 34517 16201 34529 16204
rect 34563 16201 34575 16235
rect 35342 16232 35348 16244
rect 35303 16204 35348 16232
rect 34517 16195 34575 16201
rect 35342 16192 35348 16204
rect 35400 16192 35406 16244
rect 20990 16056 20996 16108
rect 21048 16096 21054 16108
rect 22186 16096 22192 16108
rect 21048 16068 22192 16096
rect 21048 16056 21054 16068
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 32030 16096 32036 16108
rect 31991 16068 32036 16096
rect 32030 16056 32036 16068
rect 32088 16056 32094 16108
rect 32214 16056 32220 16108
rect 32272 16096 32278 16108
rect 32496 16099 32554 16105
rect 32496 16096 32508 16099
rect 32272 16068 32508 16096
rect 32272 16056 32278 16068
rect 32496 16065 32508 16068
rect 32542 16065 32554 16099
rect 32496 16059 32554 16065
rect 33226 16056 33232 16108
rect 33284 16096 33290 16108
rect 34149 16099 34207 16105
rect 34149 16096 34161 16099
rect 33284 16068 34161 16096
rect 33284 16056 33290 16068
rect 34149 16065 34161 16068
rect 34195 16065 34207 16099
rect 35360 16096 35388 16192
rect 35360 16068 35572 16096
rect 34149 16059 34207 16065
rect 19886 15988 19892 16040
rect 19944 16028 19950 16040
rect 20254 16037 20260 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19944 16000 19993 16028
rect 19944 15988 19950 16000
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 20248 16028 20260 16037
rect 20215 16000 20260 16028
rect 19981 15991 20039 15997
rect 20248 15991 20260 16000
rect 19996 15960 20024 15991
rect 20254 15988 20260 15991
rect 20312 15988 20318 16040
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 25501 16031 25559 16037
rect 25501 16028 25513 16031
rect 24912 16000 25513 16028
rect 24912 15988 24918 16000
rect 25501 15997 25513 16000
rect 25547 16028 25559 16031
rect 26053 16031 26111 16037
rect 26053 16028 26065 16031
rect 25547 16000 26065 16028
rect 25547 15997 25559 16000
rect 25501 15991 25559 15997
rect 26053 15997 26065 16000
rect 26099 15997 26111 16031
rect 26053 15991 26111 15997
rect 26973 16031 27031 16037
rect 26973 15997 26985 16031
rect 27019 16028 27031 16031
rect 27062 16028 27068 16040
rect 27019 16000 27068 16028
rect 27019 15997 27031 16000
rect 26973 15991 27031 15997
rect 27062 15988 27068 16000
rect 27120 15988 27126 16040
rect 28994 15988 29000 16040
rect 29052 16028 29058 16040
rect 29089 16031 29147 16037
rect 29089 16028 29101 16031
rect 29052 16000 29101 16028
rect 29052 15988 29058 16000
rect 29089 15997 29101 16000
rect 29135 16028 29147 16031
rect 29546 16028 29552 16040
rect 29135 16000 29552 16028
rect 29135 15997 29147 16000
rect 29089 15991 29147 15997
rect 29546 15988 29552 16000
rect 29604 15988 29610 16040
rect 32582 15988 32588 16040
rect 32640 16028 32646 16040
rect 32769 16031 32827 16037
rect 32769 16028 32781 16031
rect 32640 16000 32781 16028
rect 32640 15988 32646 16000
rect 32769 15997 32781 16000
rect 32815 15997 32827 16031
rect 32769 15991 32827 15997
rect 34330 15988 34336 16040
rect 34388 16028 34394 16040
rect 35434 16028 35440 16040
rect 34388 16000 35440 16028
rect 34388 15988 34394 16000
rect 35434 15988 35440 16000
rect 35492 15988 35498 16040
rect 35544 16028 35572 16068
rect 35693 16031 35751 16037
rect 35693 16028 35705 16031
rect 35544 16000 35705 16028
rect 35693 15997 35705 16000
rect 35739 15997 35751 16031
rect 35693 15991 35751 15997
rect 20806 15960 20812 15972
rect 19996 15932 20812 15960
rect 20806 15920 20812 15932
rect 20864 15920 20870 15972
rect 24213 15963 24271 15969
rect 24213 15960 24225 15963
rect 21008 15932 24225 15960
rect 18598 15852 18604 15904
rect 18656 15892 18662 15904
rect 18969 15895 19027 15901
rect 18969 15892 18981 15895
rect 18656 15864 18981 15892
rect 18656 15852 18662 15864
rect 18969 15861 18981 15864
rect 19015 15892 19027 15895
rect 19978 15892 19984 15904
rect 19015 15864 19984 15892
rect 19015 15861 19027 15864
rect 18969 15855 19027 15861
rect 19978 15852 19984 15864
rect 20036 15892 20042 15904
rect 21008 15892 21036 15932
rect 24213 15929 24225 15932
rect 24259 15929 24271 15963
rect 27218 15963 27276 15969
rect 27218 15960 27230 15963
rect 24213 15923 24271 15929
rect 26804 15932 27230 15960
rect 26804 15904 26832 15932
rect 27218 15929 27230 15932
rect 27264 15929 27276 15963
rect 27218 15923 27276 15929
rect 29730 15920 29736 15972
rect 29788 15969 29794 15972
rect 29788 15963 29852 15969
rect 29788 15929 29806 15963
rect 29840 15929 29852 15963
rect 35452 15960 35480 15988
rect 37093 15963 37151 15969
rect 37093 15960 37105 15963
rect 35452 15932 37105 15960
rect 29788 15923 29852 15929
rect 37093 15929 37105 15932
rect 37139 15929 37151 15963
rect 37093 15923 37151 15929
rect 29788 15920 29794 15923
rect 21726 15892 21732 15904
rect 20036 15864 21036 15892
rect 21687 15864 21732 15892
rect 20036 15852 20042 15864
rect 21726 15852 21732 15864
rect 21784 15852 21790 15904
rect 22097 15895 22155 15901
rect 22097 15861 22109 15895
rect 22143 15892 22155 15895
rect 22186 15892 22192 15904
rect 22143 15864 22192 15892
rect 22143 15861 22155 15864
rect 22097 15855 22155 15861
rect 22186 15852 22192 15864
rect 22244 15892 22250 15904
rect 24302 15892 24308 15904
rect 22244 15864 24308 15892
rect 22244 15852 22250 15864
rect 24302 15852 24308 15864
rect 24360 15852 24366 15904
rect 24949 15895 25007 15901
rect 24949 15861 24961 15895
rect 24995 15892 25007 15895
rect 25406 15892 25412 15904
rect 24995 15864 25412 15892
rect 24995 15861 25007 15864
rect 24949 15855 25007 15861
rect 25406 15852 25412 15864
rect 25464 15852 25470 15904
rect 25682 15892 25688 15904
rect 25643 15864 25688 15892
rect 25682 15852 25688 15864
rect 25740 15852 25746 15904
rect 26786 15892 26792 15904
rect 26747 15864 26792 15892
rect 26786 15852 26792 15864
rect 26844 15852 26850 15904
rect 30926 15892 30932 15904
rect 30887 15864 30932 15892
rect 30926 15852 30932 15864
rect 30984 15852 30990 15904
rect 31202 15852 31208 15904
rect 31260 15892 31266 15904
rect 31573 15895 31631 15901
rect 31573 15892 31585 15895
rect 31260 15864 31585 15892
rect 31260 15852 31266 15864
rect 31573 15861 31585 15864
rect 31619 15892 31631 15895
rect 32490 15892 32496 15904
rect 32548 15901 32554 15904
rect 31619 15864 32496 15892
rect 31619 15861 31631 15864
rect 31573 15855 31631 15861
rect 32490 15852 32496 15864
rect 32548 15892 32557 15901
rect 36814 15892 36820 15904
rect 32548 15864 32593 15892
rect 36775 15864 36820 15892
rect 32548 15855 32557 15864
rect 32548 15852 32554 15855
rect 36814 15852 36820 15864
rect 36872 15852 36878 15904
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 20073 15691 20131 15697
rect 20073 15657 20085 15691
rect 20119 15688 20131 15691
rect 20254 15688 20260 15700
rect 20119 15660 20260 15688
rect 20119 15657 20131 15660
rect 20073 15651 20131 15657
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 21726 15648 21732 15700
rect 21784 15688 21790 15700
rect 22281 15691 22339 15697
rect 22281 15688 22293 15691
rect 21784 15660 22293 15688
rect 21784 15648 21790 15660
rect 22281 15657 22293 15660
rect 22327 15657 22339 15691
rect 22281 15651 22339 15657
rect 23937 15691 23995 15697
rect 23937 15657 23949 15691
rect 23983 15688 23995 15691
rect 24302 15688 24308 15700
rect 23983 15660 24308 15688
rect 23983 15657 23995 15660
rect 23937 15651 23995 15657
rect 24302 15648 24308 15660
rect 24360 15648 24366 15700
rect 24854 15688 24860 15700
rect 24815 15660 24860 15688
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 25682 15648 25688 15700
rect 25740 15688 25746 15700
rect 26694 15688 26700 15700
rect 25740 15660 26700 15688
rect 25740 15648 25746 15660
rect 26694 15648 26700 15660
rect 26752 15688 26758 15700
rect 26881 15691 26939 15697
rect 26881 15688 26893 15691
rect 26752 15660 26893 15688
rect 26752 15648 26758 15660
rect 26881 15657 26893 15660
rect 26927 15657 26939 15691
rect 27614 15688 27620 15700
rect 27575 15660 27620 15688
rect 26881 15651 26939 15657
rect 27614 15648 27620 15660
rect 27672 15688 27678 15700
rect 28718 15688 28724 15700
rect 27672 15660 28724 15688
rect 27672 15648 27678 15660
rect 28718 15648 28724 15660
rect 28776 15648 28782 15700
rect 29641 15691 29699 15697
rect 29641 15657 29653 15691
rect 29687 15688 29699 15691
rect 29730 15688 29736 15700
rect 29687 15660 29736 15688
rect 29687 15657 29699 15660
rect 29641 15651 29699 15657
rect 29730 15648 29736 15660
rect 29788 15648 29794 15700
rect 30374 15648 30380 15700
rect 30432 15688 30438 15700
rect 30653 15691 30711 15697
rect 30653 15688 30665 15691
rect 30432 15660 30665 15688
rect 30432 15648 30438 15660
rect 30653 15657 30665 15660
rect 30699 15657 30711 15691
rect 30653 15651 30711 15657
rect 31018 15648 31024 15700
rect 31076 15688 31082 15700
rect 31573 15691 31631 15697
rect 31573 15688 31585 15691
rect 31076 15660 31585 15688
rect 31076 15648 31082 15660
rect 31573 15657 31585 15660
rect 31619 15688 31631 15691
rect 32030 15688 32036 15700
rect 31619 15660 32036 15688
rect 31619 15657 31631 15660
rect 31573 15651 31631 15657
rect 32030 15648 32036 15660
rect 32088 15648 32094 15700
rect 35710 15648 35716 15700
rect 35768 15688 35774 15700
rect 35805 15691 35863 15697
rect 35805 15688 35817 15691
rect 35768 15660 35817 15688
rect 35768 15648 35774 15660
rect 35805 15657 35817 15660
rect 35851 15657 35863 15691
rect 35805 15651 35863 15657
rect 19334 15580 19340 15632
rect 19392 15620 19398 15632
rect 20898 15620 20904 15632
rect 19392 15592 20904 15620
rect 19392 15580 19398 15592
rect 20898 15580 20904 15592
rect 20956 15620 20962 15632
rect 21146 15623 21204 15629
rect 21146 15620 21158 15623
rect 20956 15592 21158 15620
rect 20956 15580 20962 15592
rect 21146 15589 21158 15592
rect 21192 15620 21204 15623
rect 22002 15620 22008 15632
rect 21192 15592 22008 15620
rect 21192 15589 21204 15592
rect 21146 15583 21204 15589
rect 22002 15580 22008 15592
rect 22060 15580 22066 15632
rect 25958 15620 25964 15632
rect 25919 15592 25964 15620
rect 25958 15580 25964 15592
rect 26016 15580 26022 15632
rect 26973 15623 27031 15629
rect 26973 15589 26985 15623
rect 27019 15620 27031 15623
rect 27062 15620 27068 15632
rect 27019 15592 27068 15620
rect 27019 15589 27031 15592
rect 26973 15583 27031 15589
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 28626 15620 28632 15632
rect 28587 15592 28632 15620
rect 28626 15580 28632 15592
rect 28684 15580 28690 15632
rect 30466 15580 30472 15632
rect 30524 15620 30530 15632
rect 30745 15623 30803 15629
rect 30745 15620 30757 15623
rect 30524 15592 30757 15620
rect 30524 15580 30530 15592
rect 30745 15589 30757 15592
rect 30791 15589 30803 15623
rect 30745 15583 30803 15589
rect 32398 15580 32404 15632
rect 32456 15629 32462 15632
rect 32456 15623 32520 15629
rect 32456 15589 32474 15623
rect 32508 15589 32520 15623
rect 35820 15620 35848 15651
rect 35894 15648 35900 15700
rect 35952 15688 35958 15700
rect 36633 15691 36691 15697
rect 36633 15688 36645 15691
rect 35952 15660 36645 15688
rect 35952 15648 35958 15660
rect 36633 15657 36645 15660
rect 36679 15657 36691 15691
rect 36633 15651 36691 15657
rect 36081 15623 36139 15629
rect 36081 15620 36093 15623
rect 35820 15592 36093 15620
rect 32456 15583 32520 15589
rect 36081 15589 36093 15592
rect 36127 15589 36139 15623
rect 36081 15583 36139 15589
rect 32456 15580 32462 15583
rect 23845 15555 23903 15561
rect 23845 15521 23857 15555
rect 23891 15552 23903 15555
rect 24121 15555 24179 15561
rect 24121 15552 24133 15555
rect 23891 15524 24133 15552
rect 23891 15521 23903 15524
rect 23845 15515 23903 15521
rect 24121 15521 24133 15524
rect 24167 15552 24179 15555
rect 24670 15552 24676 15564
rect 24167 15524 24676 15552
rect 24167 15521 24179 15524
rect 24121 15515 24179 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 24765 15555 24823 15561
rect 24765 15521 24777 15555
rect 24811 15552 24823 15555
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 24811 15524 25237 15552
rect 24811 15521 24823 15524
rect 24765 15515 24823 15521
rect 25225 15521 25237 15524
rect 25271 15552 25283 15555
rect 25866 15552 25872 15564
rect 25271 15524 25872 15552
rect 25271 15521 25283 15524
rect 25225 15515 25283 15521
rect 25866 15512 25872 15524
rect 25924 15512 25930 15564
rect 32217 15555 32275 15561
rect 32217 15521 32229 15555
rect 32263 15552 32275 15555
rect 32263 15524 33916 15552
rect 32263 15521 32275 15524
rect 32217 15515 32275 15521
rect 33888 15496 33916 15524
rect 34238 15512 34244 15564
rect 34296 15552 34302 15564
rect 34681 15555 34739 15561
rect 34681 15552 34693 15555
rect 34296 15524 34693 15552
rect 34296 15512 34302 15524
rect 34681 15521 34693 15524
rect 34727 15521 34739 15555
rect 34681 15515 34739 15521
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15484 20499 15487
rect 20806 15484 20812 15496
rect 20487 15456 20812 15484
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 20806 15444 20812 15456
rect 20864 15484 20870 15496
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 20864 15456 20913 15484
rect 20864 15444 20870 15456
rect 20901 15453 20913 15456
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 24946 15444 24952 15496
rect 25004 15484 25010 15496
rect 25317 15487 25375 15493
rect 25317 15484 25329 15487
rect 25004 15456 25329 15484
rect 25004 15444 25010 15456
rect 25317 15453 25329 15456
rect 25363 15453 25375 15487
rect 25317 15447 25375 15453
rect 25406 15444 25412 15496
rect 25464 15484 25470 15496
rect 25501 15487 25559 15493
rect 25501 15484 25513 15487
rect 25464 15456 25513 15484
rect 25464 15444 25470 15456
rect 25501 15453 25513 15456
rect 25547 15484 25559 15487
rect 26142 15484 26148 15496
rect 25547 15456 26148 15484
rect 25547 15453 25559 15456
rect 25501 15447 25559 15453
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15484 27215 15487
rect 27706 15484 27712 15496
rect 27203 15456 27712 15484
rect 27203 15453 27215 15456
rect 27157 15447 27215 15453
rect 27706 15444 27712 15456
rect 27764 15444 27770 15496
rect 28905 15487 28963 15493
rect 28905 15453 28917 15487
rect 28951 15484 28963 15487
rect 28994 15484 29000 15496
rect 28951 15456 29000 15484
rect 28951 15453 28963 15456
rect 28905 15447 28963 15453
rect 28994 15444 29000 15456
rect 29052 15444 29058 15496
rect 30926 15484 30932 15496
rect 30887 15456 30932 15484
rect 30926 15444 30932 15456
rect 30984 15444 30990 15496
rect 33870 15444 33876 15496
rect 33928 15484 33934 15496
rect 34330 15484 34336 15496
rect 33928 15456 34336 15484
rect 33928 15444 33934 15456
rect 34330 15444 34336 15456
rect 34388 15484 34394 15496
rect 34425 15487 34483 15493
rect 34425 15484 34437 15487
rect 34388 15456 34437 15484
rect 34388 15444 34394 15456
rect 34425 15453 34437 15456
rect 34471 15453 34483 15487
rect 34425 15447 34483 15453
rect 26513 15419 26571 15425
rect 26513 15385 26525 15419
rect 26559 15416 26571 15419
rect 28626 15416 28632 15428
rect 26559 15388 28632 15416
rect 26559 15385 26571 15388
rect 26513 15379 26571 15385
rect 28626 15376 28632 15388
rect 28684 15376 28690 15428
rect 29546 15376 29552 15428
rect 29604 15416 29610 15428
rect 30009 15419 30067 15425
rect 30009 15416 30021 15419
rect 29604 15388 30021 15416
rect 29604 15376 29610 15388
rect 30009 15385 30021 15388
rect 30055 15416 30067 15419
rect 31110 15416 31116 15428
rect 30055 15388 31116 15416
rect 30055 15385 30067 15388
rect 30009 15379 30067 15385
rect 31110 15376 31116 15388
rect 31168 15376 31174 15428
rect 28261 15351 28319 15357
rect 28261 15317 28273 15351
rect 28307 15348 28319 15351
rect 28810 15348 28816 15360
rect 28307 15320 28816 15348
rect 28307 15317 28319 15320
rect 28261 15311 28319 15317
rect 28810 15308 28816 15320
rect 28868 15308 28874 15360
rect 30282 15348 30288 15360
rect 30243 15320 30288 15348
rect 30282 15308 30288 15320
rect 30340 15308 30346 15360
rect 31941 15351 31999 15357
rect 31941 15317 31953 15351
rect 31987 15348 31999 15351
rect 32582 15348 32588 15360
rect 31987 15320 32588 15348
rect 31987 15317 31999 15320
rect 31941 15311 31999 15317
rect 32582 15308 32588 15320
rect 32640 15308 32646 15360
rect 33597 15351 33655 15357
rect 33597 15317 33609 15351
rect 33643 15348 33655 15351
rect 34238 15348 34244 15360
rect 33643 15320 34244 15348
rect 33643 15317 33655 15320
rect 33597 15311 33655 15317
rect 34238 15308 34244 15320
rect 34296 15308 34302 15360
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 20898 15144 20904 15156
rect 20859 15116 20904 15144
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 23845 15147 23903 15153
rect 23845 15113 23857 15147
rect 23891 15144 23903 15147
rect 24946 15144 24952 15156
rect 23891 15116 24952 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 24946 15104 24952 15116
rect 25004 15104 25010 15156
rect 27525 15147 27583 15153
rect 27525 15113 27537 15147
rect 27571 15144 27583 15147
rect 27706 15144 27712 15156
rect 27571 15116 27712 15144
rect 27571 15113 27583 15116
rect 27525 15107 27583 15113
rect 27706 15104 27712 15116
rect 27764 15104 27770 15156
rect 28442 15144 28448 15156
rect 28403 15116 28448 15144
rect 28442 15104 28448 15116
rect 28500 15104 28506 15156
rect 28718 15144 28724 15156
rect 28679 15116 28724 15144
rect 28718 15104 28724 15116
rect 28776 15104 28782 15156
rect 28994 15104 29000 15156
rect 29052 15144 29058 15156
rect 29457 15147 29515 15153
rect 29457 15144 29469 15147
rect 29052 15116 29469 15144
rect 29052 15104 29058 15116
rect 29457 15113 29469 15116
rect 29503 15144 29515 15147
rect 29825 15147 29883 15153
rect 29825 15144 29837 15147
rect 29503 15116 29837 15144
rect 29503 15113 29515 15116
rect 29457 15107 29515 15113
rect 29825 15113 29837 15116
rect 29871 15113 29883 15147
rect 30374 15144 30380 15156
rect 30335 15116 30380 15144
rect 29825 15107 29883 15113
rect 30374 15104 30380 15116
rect 30432 15104 30438 15156
rect 30745 15147 30803 15153
rect 30745 15113 30757 15147
rect 30791 15144 30803 15147
rect 30926 15144 30932 15156
rect 30791 15116 30932 15144
rect 30791 15113 30803 15116
rect 30745 15107 30803 15113
rect 30926 15104 30932 15116
rect 30984 15144 30990 15156
rect 31021 15147 31079 15153
rect 31021 15144 31033 15147
rect 30984 15116 31033 15144
rect 30984 15104 30990 15116
rect 31021 15113 31033 15116
rect 31067 15113 31079 15147
rect 31021 15107 31079 15113
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 21269 15079 21327 15085
rect 21269 15076 21281 15079
rect 20864 15048 21281 15076
rect 20864 15036 20870 15048
rect 21269 15045 21281 15048
rect 21315 15045 21327 15079
rect 21269 15039 21327 15045
rect 24397 15011 24455 15017
rect 24397 15008 24409 15011
rect 23032 14980 24409 15008
rect 22094 14764 22100 14816
rect 22152 14804 22158 14816
rect 23032 14813 23060 14980
rect 24397 14977 24409 14980
rect 24443 15008 24455 15011
rect 25314 15008 25320 15020
rect 24443 14980 25320 15008
rect 24443 14977 24455 14980
rect 24397 14971 24455 14977
rect 25314 14968 25320 14980
rect 25372 14968 25378 15020
rect 31036 15008 31064 15107
rect 32398 15104 32404 15156
rect 32456 15144 32462 15156
rect 32585 15147 32643 15153
rect 32585 15144 32597 15147
rect 32456 15116 32597 15144
rect 32456 15104 32462 15116
rect 32585 15113 32597 15116
rect 32631 15144 32643 15147
rect 32861 15147 32919 15153
rect 32861 15144 32873 15147
rect 32631 15116 32873 15144
rect 32631 15113 32643 15116
rect 32585 15107 32643 15113
rect 32861 15113 32873 15116
rect 32907 15113 32919 15147
rect 32861 15107 32919 15113
rect 33134 15104 33140 15156
rect 33192 15144 33198 15156
rect 33229 15147 33287 15153
rect 33229 15144 33241 15147
rect 33192 15116 33241 15144
rect 33192 15104 33198 15116
rect 33229 15113 33241 15116
rect 33275 15113 33287 15147
rect 34238 15144 34244 15156
rect 34199 15116 34244 15144
rect 33229 15107 33287 15113
rect 34238 15104 34244 15116
rect 34296 15104 34302 15156
rect 34422 15104 34428 15156
rect 34480 15144 34486 15156
rect 34517 15147 34575 15153
rect 34517 15144 34529 15147
rect 34480 15116 34529 15144
rect 34480 15104 34486 15116
rect 34517 15113 34529 15116
rect 34563 15144 34575 15147
rect 34609 15147 34667 15153
rect 34609 15144 34621 15147
rect 34563 15116 34621 15144
rect 34563 15113 34575 15116
rect 34517 15107 34575 15113
rect 34609 15113 34621 15116
rect 34655 15113 34667 15147
rect 34609 15107 34667 15113
rect 31036 14980 31340 15008
rect 25406 14940 25412 14952
rect 25319 14912 25412 14940
rect 25406 14900 25412 14912
rect 25464 14940 25470 14952
rect 25958 14940 25964 14952
rect 25464 14912 25964 14940
rect 25464 14900 25470 14912
rect 25958 14900 25964 14912
rect 26016 14900 26022 14952
rect 27801 14943 27859 14949
rect 27801 14909 27813 14943
rect 27847 14940 27859 14943
rect 28442 14940 28448 14952
rect 27847 14912 28448 14940
rect 27847 14909 27859 14912
rect 27801 14903 27859 14909
rect 28442 14900 28448 14912
rect 28500 14900 28506 14952
rect 28994 14900 29000 14952
rect 29052 14940 29058 14952
rect 29273 14943 29331 14949
rect 29273 14940 29285 14943
rect 29052 14912 29285 14940
rect 29052 14900 29058 14912
rect 29273 14909 29285 14912
rect 29319 14909 29331 14943
rect 29273 14903 29331 14909
rect 31110 14900 31116 14952
rect 31168 14940 31174 14952
rect 31205 14943 31263 14949
rect 31205 14940 31217 14943
rect 31168 14912 31217 14940
rect 31168 14900 31174 14912
rect 31205 14909 31217 14912
rect 31251 14909 31263 14943
rect 31312 14940 31340 14980
rect 33042 14968 33048 15020
rect 33100 15008 33106 15020
rect 33413 15011 33471 15017
rect 33413 15008 33425 15011
rect 33100 14980 33425 15008
rect 33100 14968 33106 14980
rect 33413 14977 33425 14980
rect 33459 14977 33471 15011
rect 33413 14971 33471 14977
rect 34238 14968 34244 15020
rect 34296 15008 34302 15020
rect 35437 15011 35495 15017
rect 35437 15008 35449 15011
rect 34296 14980 35449 15008
rect 34296 14968 34302 14980
rect 35437 14977 35449 14980
rect 35483 14977 35495 15011
rect 35437 14971 35495 14977
rect 31461 14943 31519 14949
rect 31461 14940 31473 14943
rect 31312 14912 31473 14940
rect 31205 14903 31263 14909
rect 31461 14909 31473 14912
rect 31507 14909 31519 14943
rect 31461 14903 31519 14909
rect 34517 14943 34575 14949
rect 34517 14909 34529 14943
rect 34563 14940 34575 14943
rect 35253 14943 35311 14949
rect 35253 14940 35265 14943
rect 34563 14912 35265 14940
rect 34563 14909 34575 14912
rect 34517 14903 34575 14909
rect 35253 14909 35265 14912
rect 35299 14909 35311 14943
rect 35253 14903 35311 14909
rect 24305 14875 24363 14881
rect 24305 14872 24317 14875
rect 23492 14844 24317 14872
rect 23492 14816 23520 14844
rect 24305 14841 24317 14844
rect 24351 14841 24363 14875
rect 24305 14835 24363 14841
rect 25317 14875 25375 14881
rect 25317 14841 25329 14875
rect 25363 14872 25375 14875
rect 25590 14872 25596 14884
rect 25363 14844 25596 14872
rect 25363 14841 25375 14844
rect 25317 14835 25375 14841
rect 25590 14832 25596 14844
rect 25648 14881 25654 14884
rect 25648 14875 25712 14881
rect 25648 14841 25666 14875
rect 25700 14841 25712 14875
rect 25648 14835 25712 14841
rect 25648 14832 25654 14835
rect 23017 14807 23075 14813
rect 23017 14804 23029 14807
rect 22152 14776 23029 14804
rect 22152 14764 22158 14776
rect 23017 14773 23029 14776
rect 23063 14773 23075 14807
rect 23474 14804 23480 14816
rect 23435 14776 23480 14804
rect 23017 14767 23075 14773
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 24210 14804 24216 14816
rect 24171 14776 24216 14804
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 26234 14764 26240 14816
rect 26292 14804 26298 14816
rect 26786 14804 26792 14816
rect 26292 14776 26792 14804
rect 26292 14764 26298 14776
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 27062 14804 27068 14816
rect 27023 14776 27068 14804
rect 27062 14764 27068 14776
rect 27120 14764 27126 14816
rect 27614 14764 27620 14816
rect 27672 14804 27678 14816
rect 27985 14807 28043 14813
rect 27985 14804 27997 14807
rect 27672 14776 27997 14804
rect 27672 14764 27678 14776
rect 27985 14773 27997 14776
rect 28031 14773 28043 14807
rect 31220 14804 31248 14903
rect 34698 14832 34704 14884
rect 34756 14872 34762 14884
rect 35158 14872 35164 14884
rect 34756 14844 35164 14872
rect 34756 14832 34762 14844
rect 35158 14832 35164 14844
rect 35216 14872 35222 14884
rect 35345 14875 35403 14881
rect 35345 14872 35357 14875
rect 35216 14844 35357 14872
rect 35216 14832 35222 14844
rect 35345 14841 35357 14844
rect 35391 14841 35403 14875
rect 35345 14835 35403 14841
rect 31478 14804 31484 14816
rect 31220 14776 31484 14804
rect 27985 14767 28043 14773
rect 31478 14764 31484 14776
rect 31536 14764 31542 14816
rect 33870 14804 33876 14816
rect 33831 14776 33876 14804
rect 33870 14764 33876 14776
rect 33928 14764 33934 14816
rect 34885 14807 34943 14813
rect 34885 14773 34897 14807
rect 34931 14804 34943 14807
rect 35526 14804 35532 14816
rect 34931 14776 35532 14804
rect 34931 14773 34943 14776
rect 34885 14767 34943 14773
rect 35526 14764 35532 14776
rect 35584 14804 35590 14816
rect 35986 14804 35992 14816
rect 35584 14776 35992 14804
rect 35584 14764 35590 14776
rect 35986 14764 35992 14776
rect 36044 14764 36050 14816
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 23290 14600 23296 14612
rect 23251 14572 23296 14600
rect 23290 14560 23296 14572
rect 23348 14560 23354 14612
rect 23937 14603 23995 14609
rect 23937 14569 23949 14603
rect 23983 14600 23995 14603
rect 24210 14600 24216 14612
rect 23983 14572 24216 14600
rect 23983 14569 23995 14572
rect 23937 14563 23995 14569
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 25590 14600 25596 14612
rect 25551 14572 25596 14600
rect 25590 14560 25596 14572
rect 25648 14560 25654 14612
rect 26694 14600 26700 14612
rect 26655 14572 26700 14600
rect 26694 14560 26700 14572
rect 26752 14560 26758 14612
rect 27065 14603 27123 14609
rect 27065 14569 27077 14603
rect 27111 14600 27123 14603
rect 27522 14600 27528 14612
rect 27111 14572 27528 14600
rect 27111 14569 27123 14572
rect 27065 14563 27123 14569
rect 27522 14560 27528 14572
rect 27580 14560 27586 14612
rect 28353 14603 28411 14609
rect 28353 14569 28365 14603
rect 28399 14600 28411 14603
rect 28626 14600 28632 14612
rect 28399 14572 28632 14600
rect 28399 14569 28411 14572
rect 28353 14563 28411 14569
rect 28626 14560 28632 14572
rect 28684 14560 28690 14612
rect 28994 14560 29000 14612
rect 29052 14600 29058 14612
rect 29273 14603 29331 14609
rect 29273 14600 29285 14603
rect 29052 14572 29285 14600
rect 29052 14560 29058 14572
rect 29273 14569 29285 14572
rect 29319 14569 29331 14603
rect 29914 14600 29920 14612
rect 29875 14572 29920 14600
rect 29273 14563 29331 14569
rect 29914 14560 29920 14572
rect 29972 14560 29978 14612
rect 30466 14560 30472 14612
rect 30524 14600 30530 14612
rect 30653 14603 30711 14609
rect 30653 14600 30665 14603
rect 30524 14572 30665 14600
rect 30524 14560 30530 14572
rect 30653 14569 30665 14572
rect 30699 14569 30711 14603
rect 30653 14563 30711 14569
rect 32217 14603 32275 14609
rect 32217 14569 32229 14603
rect 32263 14600 32275 14603
rect 32858 14600 32864 14612
rect 32263 14572 32864 14600
rect 32263 14569 32275 14572
rect 32217 14563 32275 14569
rect 32858 14560 32864 14572
rect 32916 14560 32922 14612
rect 34238 14560 34244 14612
rect 34296 14600 34302 14612
rect 34885 14603 34943 14609
rect 34885 14600 34897 14603
rect 34296 14572 34897 14600
rect 34296 14560 34302 14572
rect 34885 14569 34897 14572
rect 34931 14569 34943 14603
rect 34885 14563 34943 14569
rect 35158 14560 35164 14612
rect 35216 14600 35222 14612
rect 35253 14603 35311 14609
rect 35253 14600 35265 14603
rect 35216 14572 35265 14600
rect 35216 14560 35222 14572
rect 35253 14569 35265 14572
rect 35299 14569 35311 14603
rect 35253 14563 35311 14569
rect 24228 14532 24256 14560
rect 24458 14535 24516 14541
rect 24458 14532 24470 14535
rect 24228 14504 24470 14532
rect 24458 14501 24470 14504
rect 24504 14501 24516 14535
rect 24458 14495 24516 14501
rect 25314 14492 25320 14544
rect 25372 14532 25378 14544
rect 25869 14535 25927 14541
rect 25869 14532 25881 14535
rect 25372 14504 25881 14532
rect 25372 14492 25378 14504
rect 25869 14501 25881 14504
rect 25915 14532 25927 14535
rect 26418 14532 26424 14544
rect 25915 14504 26424 14532
rect 25915 14501 25927 14504
rect 25869 14495 25927 14501
rect 26418 14492 26424 14504
rect 26476 14492 26482 14544
rect 28810 14492 28816 14544
rect 28868 14532 28874 14544
rect 32677 14535 32735 14541
rect 28868 14504 29776 14532
rect 28868 14492 28874 14504
rect 23106 14464 23112 14476
rect 23067 14436 23112 14464
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 23658 14424 23664 14476
rect 23716 14464 23722 14476
rect 24213 14467 24271 14473
rect 24213 14464 24225 14467
rect 23716 14436 24225 14464
rect 23716 14424 23722 14436
rect 24213 14433 24225 14436
rect 24259 14464 24271 14467
rect 24302 14464 24308 14476
rect 24259 14436 24308 14464
rect 24259 14433 24271 14436
rect 24213 14427 24271 14433
rect 24302 14424 24308 14436
rect 24360 14424 24366 14476
rect 27154 14424 27160 14476
rect 27212 14464 27218 14476
rect 27433 14467 27491 14473
rect 27433 14464 27445 14467
rect 27212 14436 27445 14464
rect 27212 14424 27218 14436
rect 27433 14433 27445 14436
rect 27479 14433 27491 14467
rect 27433 14427 27491 14433
rect 28629 14467 28687 14473
rect 28629 14433 28641 14467
rect 28675 14464 28687 14467
rect 29086 14464 29092 14476
rect 28675 14436 29092 14464
rect 28675 14433 28687 14436
rect 28629 14427 28687 14433
rect 29086 14424 29092 14436
rect 29144 14424 29150 14476
rect 29748 14473 29776 14504
rect 32677 14501 32689 14535
rect 32723 14532 32735 14535
rect 32766 14532 32772 14544
rect 32723 14504 32772 14532
rect 32723 14501 32735 14504
rect 32677 14495 32735 14501
rect 32766 14492 32772 14504
rect 32824 14492 32830 14544
rect 29733 14467 29791 14473
rect 29733 14433 29745 14467
rect 29779 14464 29791 14467
rect 31294 14464 31300 14476
rect 29779 14436 31300 14464
rect 29779 14433 29791 14436
rect 29733 14427 29791 14433
rect 31294 14424 31300 14436
rect 31352 14424 31358 14476
rect 32582 14464 32588 14476
rect 32543 14436 32588 14464
rect 32582 14424 32588 14436
rect 32640 14424 32646 14476
rect 27522 14396 27528 14408
rect 27483 14368 27528 14396
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 27706 14396 27712 14408
rect 27667 14368 27712 14396
rect 27706 14356 27712 14368
rect 27764 14356 27770 14408
rect 32861 14399 32919 14405
rect 32861 14365 32873 14399
rect 32907 14396 32919 14399
rect 32950 14396 32956 14408
rect 32907 14368 32956 14396
rect 32907 14365 32919 14368
rect 32861 14359 32919 14365
rect 32950 14356 32956 14368
rect 33008 14356 33014 14408
rect 21358 14260 21364 14272
rect 21319 14232 21364 14260
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 24394 14260 24400 14272
rect 24176 14232 24400 14260
rect 24176 14220 24182 14232
rect 24394 14220 24400 14232
rect 24452 14220 24458 14272
rect 27890 14220 27896 14272
rect 27948 14260 27954 14272
rect 28813 14263 28871 14269
rect 28813 14260 28825 14263
rect 27948 14232 28825 14260
rect 27948 14220 27954 14232
rect 28813 14229 28825 14232
rect 28859 14229 28871 14263
rect 30374 14260 30380 14272
rect 30335 14232 30380 14260
rect 28813 14223 28871 14229
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 31297 14263 31355 14269
rect 31297 14229 31309 14263
rect 31343 14260 31355 14263
rect 31478 14260 31484 14272
rect 31343 14232 31484 14260
rect 31343 14229 31355 14232
rect 31297 14223 31355 14229
rect 31478 14220 31484 14232
rect 31536 14260 31542 14272
rect 33502 14260 33508 14272
rect 31536 14232 33508 14260
rect 31536 14220 31542 14232
rect 33502 14220 33508 14232
rect 33560 14260 33566 14272
rect 33870 14260 33876 14272
rect 33560 14232 33876 14260
rect 33560 14220 33566 14232
rect 33870 14220 33876 14232
rect 33928 14260 33934 14272
rect 34425 14263 34483 14269
rect 34425 14260 34437 14263
rect 33928 14232 34437 14260
rect 33928 14220 33934 14232
rect 34425 14229 34437 14232
rect 34471 14229 34483 14263
rect 34425 14223 34483 14229
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 24302 14016 24308 14068
rect 24360 14056 24366 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 24360 14028 25053 14056
rect 24360 14016 24366 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25406 14056 25412 14068
rect 25367 14028 25412 14056
rect 25041 14019 25099 14025
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 25590 14016 25596 14068
rect 25648 14056 25654 14068
rect 25685 14059 25743 14065
rect 25685 14056 25697 14059
rect 25648 14028 25697 14056
rect 25648 14016 25654 14028
rect 25685 14025 25697 14028
rect 25731 14025 25743 14059
rect 25866 14056 25872 14068
rect 25827 14028 25872 14056
rect 25685 14019 25743 14025
rect 21358 13920 21364 13932
rect 21319 13892 21364 13920
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 23492 13920 23520 14016
rect 25700 13920 25728 14019
rect 25866 14016 25872 14028
rect 25924 14016 25930 14068
rect 27157 14059 27215 14065
rect 27157 14025 27169 14059
rect 27203 14056 27215 14059
rect 27522 14056 27528 14068
rect 27203 14028 27528 14056
rect 27203 14025 27215 14028
rect 27157 14019 27215 14025
rect 27522 14016 27528 14028
rect 27580 14056 27586 14068
rect 27617 14059 27675 14065
rect 27617 14056 27629 14059
rect 27580 14028 27629 14056
rect 27580 14016 27586 14028
rect 27617 14025 27629 14028
rect 27663 14025 27675 14059
rect 27617 14019 27675 14025
rect 27706 14016 27712 14068
rect 27764 14056 27770 14068
rect 28353 14059 28411 14065
rect 28353 14056 28365 14059
rect 27764 14028 28365 14056
rect 27764 14016 27770 14028
rect 28353 14025 28365 14028
rect 28399 14025 28411 14059
rect 29086 14056 29092 14068
rect 29047 14028 29092 14056
rect 28353 14019 28411 14025
rect 29086 14016 29092 14028
rect 29144 14016 29150 14068
rect 29178 14016 29184 14068
rect 29236 14056 29242 14068
rect 29733 14059 29791 14065
rect 29733 14056 29745 14059
rect 29236 14028 29745 14056
rect 29236 14016 29242 14028
rect 29733 14025 29745 14028
rect 29779 14025 29791 14059
rect 31294 14056 31300 14068
rect 31255 14028 31300 14056
rect 29733 14019 29791 14025
rect 27890 13988 27896 14000
rect 26436 13960 27896 13988
rect 26436 13932 26464 13960
rect 27890 13948 27896 13960
rect 27948 13948 27954 14000
rect 28534 13988 28540 14000
rect 28495 13960 28540 13988
rect 28534 13948 28540 13960
rect 28592 13948 28598 14000
rect 26329 13923 26387 13929
rect 26329 13920 26341 13923
rect 23492 13892 23796 13920
rect 25700 13892 26341 13920
rect 23106 13852 23112 13864
rect 23019 13824 23112 13852
rect 23106 13812 23112 13824
rect 23164 13852 23170 13864
rect 23658 13852 23664 13864
rect 23164 13824 23428 13852
rect 23619 13824 23664 13852
rect 23164 13812 23170 13824
rect 21266 13784 21272 13796
rect 21179 13756 21272 13784
rect 21266 13744 21272 13756
rect 21324 13784 21330 13796
rect 21634 13793 21640 13796
rect 21606 13787 21640 13793
rect 21606 13784 21618 13787
rect 21324 13756 21618 13784
rect 21324 13744 21330 13756
rect 21606 13753 21618 13756
rect 21692 13784 21698 13796
rect 23400 13784 23428 13824
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 23768 13852 23796 13892
rect 26329 13889 26341 13892
rect 26375 13889 26387 13923
rect 26329 13883 26387 13889
rect 26418 13880 26424 13932
rect 26476 13920 26482 13932
rect 26476 13892 26521 13920
rect 26476 13880 26482 13892
rect 27798 13880 27804 13932
rect 27856 13920 27862 13932
rect 28626 13920 28632 13932
rect 27856 13892 28632 13920
rect 27856 13880 27862 13892
rect 28626 13880 28632 13892
rect 28684 13920 28690 13932
rect 28684 13892 28764 13920
rect 28684 13880 28690 13892
rect 23917 13855 23975 13861
rect 23917 13852 23929 13855
rect 23768 13824 23929 13852
rect 23917 13821 23929 13824
rect 23963 13852 23975 13855
rect 27430 13852 27436 13864
rect 23963 13821 23980 13852
rect 27391 13824 27436 13852
rect 23917 13815 23980 13821
rect 23474 13784 23480 13796
rect 21692 13756 21754 13784
rect 23400 13756 23480 13784
rect 21606 13747 21640 13753
rect 21634 13744 21640 13747
rect 21692 13744 21698 13756
rect 23474 13744 23480 13756
rect 23532 13744 23538 13796
rect 23952 13784 23980 13815
rect 27430 13812 27436 13824
rect 27488 13852 27494 13864
rect 28736 13861 28764 13892
rect 27985 13855 28043 13861
rect 27985 13852 27997 13855
rect 27488 13824 27997 13852
rect 27488 13812 27494 13824
rect 27985 13821 27997 13824
rect 28031 13821 28043 13855
rect 27985 13815 28043 13821
rect 28721 13855 28779 13861
rect 28721 13821 28733 13855
rect 28767 13821 28779 13855
rect 29748 13852 29776 14019
rect 31294 14016 31300 14028
rect 31352 14016 31358 14068
rect 31478 14056 31484 14068
rect 31439 14028 31484 14056
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 32677 14059 32735 14065
rect 32677 14025 32689 14059
rect 32723 14056 32735 14059
rect 32766 14056 32772 14068
rect 32723 14028 32772 14056
rect 32723 14025 32735 14028
rect 32677 14019 32735 14025
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 32950 14056 32956 14068
rect 32911 14028 32956 14056
rect 32950 14016 32956 14028
rect 33008 14016 33014 14068
rect 31754 13988 31760 14000
rect 30392 13960 31760 13988
rect 30392 13932 30420 13960
rect 31754 13948 31760 13960
rect 31812 13948 31818 14000
rect 30374 13920 30380 13932
rect 30335 13892 30380 13920
rect 30374 13880 30380 13892
rect 30432 13880 30438 13932
rect 30561 13923 30619 13929
rect 30561 13889 30573 13923
rect 30607 13889 30619 13923
rect 30561 13883 30619 13889
rect 30282 13852 30288 13864
rect 29748 13824 30288 13852
rect 28721 13815 28779 13821
rect 30282 13812 30288 13824
rect 30340 13812 30346 13864
rect 30576 13852 30604 13883
rect 31021 13855 31079 13861
rect 31021 13852 31033 13855
rect 30576 13824 31033 13852
rect 31021 13821 31033 13824
rect 31067 13852 31079 13855
rect 31110 13852 31116 13864
rect 31067 13824 31116 13852
rect 31067 13821 31079 13824
rect 31021 13815 31079 13821
rect 31110 13812 31116 13824
rect 31168 13812 31174 13864
rect 31662 13852 31668 13864
rect 31623 13824 31668 13852
rect 31662 13812 31668 13824
rect 31720 13812 31726 13864
rect 24118 13784 24124 13796
rect 23952 13756 24124 13784
rect 24118 13744 24124 13756
rect 24176 13744 24182 13796
rect 22741 13719 22799 13725
rect 22741 13685 22753 13719
rect 22787 13716 22799 13719
rect 23014 13716 23020 13728
rect 22787 13688 23020 13716
rect 22787 13685 22799 13688
rect 22741 13679 22799 13685
rect 23014 13676 23020 13688
rect 23072 13676 23078 13728
rect 26234 13716 26240 13728
rect 26195 13688 26240 13716
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 29822 13676 29828 13728
rect 29880 13716 29886 13728
rect 29917 13719 29975 13725
rect 29917 13716 29929 13719
rect 29880 13688 29929 13716
rect 29880 13676 29886 13688
rect 29917 13685 29929 13688
rect 29963 13685 29975 13719
rect 29917 13679 29975 13685
rect 32309 13719 32367 13725
rect 32309 13685 32321 13719
rect 32355 13716 32367 13719
rect 32582 13716 32588 13728
rect 32355 13688 32588 13716
rect 32355 13685 32367 13688
rect 32309 13679 32367 13685
rect 32582 13676 32588 13688
rect 32640 13676 32646 13728
rect 34422 13676 34428 13728
rect 34480 13716 34486 13728
rect 34885 13719 34943 13725
rect 34885 13716 34897 13719
rect 34480 13688 34897 13716
rect 34480 13676 34486 13688
rect 34885 13685 34897 13688
rect 34931 13685 34943 13719
rect 34885 13679 34943 13685
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 21634 13512 21640 13524
rect 21595 13484 21640 13512
rect 21634 13472 21640 13484
rect 21692 13512 21698 13524
rect 22002 13512 22008 13524
rect 21692 13484 22008 13512
rect 21692 13472 21698 13484
rect 22002 13472 22008 13484
rect 22060 13472 22066 13524
rect 24118 13512 24124 13524
rect 24079 13484 24124 13512
rect 24118 13472 24124 13484
rect 24176 13472 24182 13524
rect 24210 13472 24216 13524
rect 24268 13512 24274 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 24268 13484 24409 13512
rect 24268 13472 24274 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 24854 13472 24860 13524
rect 24912 13512 24918 13524
rect 25041 13515 25099 13521
rect 25041 13512 25053 13515
rect 24912 13484 25053 13512
rect 24912 13472 24918 13484
rect 25041 13481 25053 13484
rect 25087 13481 25099 13515
rect 25041 13475 25099 13481
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 27154 13512 27160 13524
rect 25547 13484 27160 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 28626 13512 28632 13524
rect 28587 13484 28632 13512
rect 28626 13472 28632 13484
rect 28684 13472 28690 13524
rect 28994 13512 29000 13524
rect 28955 13484 29000 13512
rect 28994 13472 29000 13484
rect 29052 13472 29058 13524
rect 30282 13472 30288 13524
rect 30340 13512 30346 13524
rect 30469 13515 30527 13521
rect 30469 13512 30481 13515
rect 30340 13484 30481 13512
rect 30340 13472 30346 13484
rect 30469 13481 30481 13484
rect 30515 13481 30527 13515
rect 30469 13475 30527 13481
rect 30929 13515 30987 13521
rect 30929 13481 30941 13515
rect 30975 13512 30987 13515
rect 31018 13512 31024 13524
rect 30975 13484 31024 13512
rect 30975 13481 30987 13484
rect 30929 13475 30987 13481
rect 31018 13472 31024 13484
rect 31076 13472 31082 13524
rect 31754 13472 31760 13524
rect 31812 13512 31818 13524
rect 32585 13515 32643 13521
rect 32585 13512 32597 13515
rect 31812 13484 32597 13512
rect 31812 13472 31818 13484
rect 32585 13481 32597 13484
rect 32631 13512 32643 13515
rect 32950 13512 32956 13524
rect 32631 13484 32956 13512
rect 32631 13481 32643 13484
rect 32585 13475 32643 13481
rect 32950 13472 32956 13484
rect 33008 13472 33014 13524
rect 35802 13512 35808 13524
rect 35763 13484 35808 13512
rect 35802 13472 35808 13484
rect 35860 13472 35866 13524
rect 25961 13447 26019 13453
rect 25961 13413 25973 13447
rect 26007 13444 26019 13447
rect 26234 13444 26240 13456
rect 26007 13416 26240 13444
rect 26007 13413 26019 13416
rect 25961 13407 26019 13413
rect 26234 13404 26240 13416
rect 26292 13404 26298 13456
rect 20898 13336 20904 13388
rect 20956 13376 20962 13388
rect 23014 13385 23020 13388
rect 21545 13379 21603 13385
rect 21545 13376 21557 13379
rect 20956 13348 21557 13376
rect 20956 13336 20962 13348
rect 21545 13345 21557 13348
rect 21591 13376 21603 13379
rect 23008 13376 23020 13385
rect 21591 13348 23020 13376
rect 21591 13345 21603 13348
rect 21545 13339 21603 13345
rect 23008 13339 23020 13348
rect 23014 13336 23020 13339
rect 23072 13336 23078 13388
rect 25130 13336 25136 13388
rect 25188 13376 25194 13388
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 25188 13348 25237 13376
rect 25188 13336 25194 13348
rect 25225 13345 25237 13348
rect 25271 13345 25283 13379
rect 25225 13339 25283 13345
rect 25314 13336 25320 13388
rect 25372 13376 25378 13388
rect 27709 13379 27767 13385
rect 25372 13348 25417 13376
rect 25372 13336 25378 13348
rect 27709 13345 27721 13379
rect 27755 13376 27767 13379
rect 28166 13376 28172 13388
rect 27755 13348 28172 13376
rect 27755 13345 27767 13348
rect 27709 13339 27767 13345
rect 28166 13336 28172 13348
rect 28224 13336 28230 13388
rect 29012 13376 29040 13472
rect 29273 13379 29331 13385
rect 29273 13376 29285 13379
rect 29012 13348 29285 13376
rect 29273 13345 29285 13348
rect 29319 13345 29331 13379
rect 29822 13376 29828 13388
rect 29783 13348 29828 13376
rect 29273 13339 29331 13345
rect 29822 13336 29828 13348
rect 29880 13336 29886 13388
rect 33686 13336 33692 13388
rect 33744 13376 33750 13388
rect 33853 13379 33911 13385
rect 33853 13376 33865 13379
rect 33744 13348 33865 13376
rect 33744 13336 33750 13348
rect 33853 13345 33865 13348
rect 33899 13345 33911 13379
rect 33853 13339 33911 13345
rect 36173 13379 36231 13385
rect 36173 13345 36185 13379
rect 36219 13376 36231 13379
rect 36538 13376 36544 13388
rect 36219 13348 36544 13376
rect 36219 13345 36231 13348
rect 36173 13339 36231 13345
rect 36538 13336 36544 13348
rect 36596 13336 36602 13388
rect 21726 13308 21732 13320
rect 21687 13280 21732 13308
rect 21726 13268 21732 13280
rect 21784 13308 21790 13320
rect 22094 13308 22100 13320
rect 21784 13280 22100 13308
rect 21784 13268 21790 13280
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 22741 13311 22799 13317
rect 22741 13308 22753 13311
rect 22572 13280 22753 13308
rect 21174 13172 21180 13184
rect 21135 13144 21180 13172
rect 21174 13132 21180 13144
rect 21232 13132 21238 13184
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 22572 13181 22600 13280
rect 22741 13277 22753 13280
rect 22787 13277 22799 13311
rect 22741 13271 22799 13277
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13308 24915 13311
rect 25406 13308 25412 13320
rect 24903 13280 25412 13308
rect 24903 13277 24915 13280
rect 24857 13271 24915 13277
rect 25406 13268 25412 13280
rect 25464 13268 25470 13320
rect 27798 13308 27804 13320
rect 27759 13280 27804 13308
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 27890 13268 27896 13320
rect 27948 13308 27954 13320
rect 27948 13280 27993 13308
rect 27948 13268 27954 13280
rect 29178 13268 29184 13320
rect 29236 13308 29242 13320
rect 29730 13308 29736 13320
rect 29236 13280 29736 13308
rect 29236 13268 29242 13280
rect 29730 13268 29736 13280
rect 29788 13308 29794 13320
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 29788 13280 29929 13308
rect 29788 13268 29794 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 30006 13268 30012 13320
rect 30064 13308 30070 13320
rect 30064 13280 30109 13308
rect 30064 13268 30070 13280
rect 33502 13268 33508 13320
rect 33560 13308 33566 13320
rect 33597 13311 33655 13317
rect 33597 13308 33609 13311
rect 33560 13280 33609 13308
rect 33560 13268 33566 13280
rect 33597 13277 33609 13280
rect 33643 13277 33655 13311
rect 33597 13271 33655 13277
rect 35710 13268 35716 13320
rect 35768 13308 35774 13320
rect 36265 13311 36323 13317
rect 36265 13308 36277 13311
rect 35768 13280 36277 13308
rect 35768 13268 35774 13280
rect 36265 13277 36277 13280
rect 36311 13277 36323 13311
rect 36446 13308 36452 13320
rect 36407 13280 36452 13308
rect 36265 13271 36323 13277
rect 29089 13243 29147 13249
rect 29089 13209 29101 13243
rect 29135 13240 29147 13243
rect 30650 13240 30656 13252
rect 29135 13212 30656 13240
rect 29135 13209 29147 13212
rect 29089 13203 29147 13209
rect 30650 13200 30656 13212
rect 30708 13240 30714 13252
rect 31481 13243 31539 13249
rect 31481 13240 31493 13243
rect 30708 13212 31493 13240
rect 30708 13200 30714 13212
rect 31481 13209 31493 13212
rect 31527 13240 31539 13243
rect 31662 13240 31668 13252
rect 31527 13212 31668 13240
rect 31527 13209 31539 13212
rect 31481 13203 31539 13209
rect 31662 13200 31668 13212
rect 31720 13200 31726 13252
rect 36280 13240 36308 13271
rect 36446 13268 36452 13280
rect 36504 13268 36510 13320
rect 37550 13240 37556 13252
rect 36280 13212 37556 13240
rect 37550 13200 37556 13212
rect 37608 13200 37614 13252
rect 22557 13175 22615 13181
rect 22557 13172 22569 13175
rect 22244 13144 22569 13172
rect 22244 13132 22250 13144
rect 22557 13141 22569 13144
rect 22603 13141 22615 13175
rect 22557 13135 22615 13141
rect 27246 13132 27252 13184
rect 27304 13172 27310 13184
rect 27341 13175 27399 13181
rect 27341 13172 27353 13175
rect 27304 13144 27353 13172
rect 27304 13132 27310 13144
rect 27341 13141 27353 13144
rect 27387 13141 27399 13175
rect 29454 13172 29460 13184
rect 29415 13144 29460 13172
rect 27341 13135 27399 13141
rect 29454 13132 29460 13144
rect 29512 13132 29518 13184
rect 34698 13132 34704 13184
rect 34756 13172 34762 13184
rect 34977 13175 35035 13181
rect 34977 13172 34989 13175
rect 34756 13144 34989 13172
rect 34756 13132 34762 13144
rect 34977 13141 34989 13144
rect 35023 13141 35035 13175
rect 35342 13172 35348 13184
rect 35255 13144 35348 13172
rect 34977 13135 35035 13141
rect 35342 13132 35348 13144
rect 35400 13172 35406 13184
rect 36262 13172 36268 13184
rect 35400 13144 36268 13172
rect 35400 13132 35406 13144
rect 36262 13132 36268 13144
rect 36320 13132 36326 13184
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 20533 12971 20591 12977
rect 20533 12937 20545 12971
rect 20579 12968 20591 12971
rect 21726 12968 21732 12980
rect 20579 12940 21732 12968
rect 20579 12937 20591 12940
rect 20533 12931 20591 12937
rect 21726 12928 21732 12940
rect 21784 12928 21790 12980
rect 22002 12928 22008 12980
rect 22060 12968 22066 12980
rect 22741 12971 22799 12977
rect 22741 12968 22753 12971
rect 22060 12940 22753 12968
rect 22060 12928 22066 12940
rect 22741 12937 22753 12940
rect 22787 12937 22799 12971
rect 23014 12968 23020 12980
rect 22975 12940 23020 12968
rect 22741 12931 22799 12937
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 23661 12971 23719 12977
rect 23661 12968 23673 12971
rect 23532 12940 23673 12968
rect 23532 12928 23538 12940
rect 23661 12937 23673 12940
rect 23707 12937 23719 12971
rect 24762 12968 24768 12980
rect 24723 12940 24768 12968
rect 23661 12931 23719 12937
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25130 12968 25136 12980
rect 25091 12940 25136 12968
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 26789 12971 26847 12977
rect 26789 12937 26801 12971
rect 26835 12968 26847 12971
rect 27430 12968 27436 12980
rect 26835 12940 27436 12968
rect 26835 12937 26847 12940
rect 26789 12931 26847 12937
rect 27430 12928 27436 12940
rect 27488 12928 27494 12980
rect 27798 12968 27804 12980
rect 27759 12940 27804 12968
rect 27798 12928 27804 12940
rect 27856 12928 27862 12980
rect 28166 12968 28172 12980
rect 28127 12940 28172 12968
rect 28166 12928 28172 12940
rect 28224 12928 28230 12980
rect 29089 12971 29147 12977
rect 29089 12937 29101 12971
rect 29135 12968 29147 12971
rect 29362 12968 29368 12980
rect 29135 12940 29368 12968
rect 29135 12937 29147 12940
rect 29089 12931 29147 12937
rect 29362 12928 29368 12940
rect 29420 12968 29426 12980
rect 29822 12968 29828 12980
rect 29420 12940 29828 12968
rect 29420 12928 29426 12940
rect 29822 12928 29828 12940
rect 29880 12928 29886 12980
rect 29914 12928 29920 12980
rect 29972 12968 29978 12980
rect 31018 12968 31024 12980
rect 29972 12940 31024 12968
rect 29972 12928 29978 12940
rect 31018 12928 31024 12940
rect 31076 12928 31082 12980
rect 32125 12971 32183 12977
rect 32125 12937 32137 12971
rect 32171 12968 32183 12971
rect 34698 12968 34704 12980
rect 32171 12940 33180 12968
rect 34659 12940 34704 12968
rect 32171 12937 32183 12940
rect 32125 12931 32183 12937
rect 20898 12900 20904 12912
rect 20859 12872 20904 12900
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 21266 12900 21272 12912
rect 21227 12872 21272 12900
rect 21266 12860 21272 12872
rect 21324 12860 21330 12912
rect 21358 12832 21364 12844
rect 21319 12804 21364 12832
rect 21358 12792 21364 12804
rect 21416 12792 21422 12844
rect 24305 12835 24363 12841
rect 24305 12801 24317 12835
rect 24351 12832 24363 12835
rect 24670 12832 24676 12844
rect 24351 12804 24676 12832
rect 24351 12801 24363 12804
rect 24305 12795 24363 12801
rect 24670 12792 24676 12804
rect 24728 12832 24734 12844
rect 24780 12832 24808 12928
rect 26142 12860 26148 12912
rect 26200 12900 26206 12912
rect 26329 12903 26387 12909
rect 26329 12900 26341 12903
rect 26200 12872 26341 12900
rect 26200 12860 26206 12872
rect 26329 12869 26341 12872
rect 26375 12900 26387 12903
rect 26375 12872 27476 12900
rect 26375 12869 26387 12872
rect 26329 12863 26387 12869
rect 24728 12804 24808 12832
rect 24728 12792 24734 12804
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 26697 12835 26755 12841
rect 24912 12804 25452 12832
rect 24912 12792 24918 12804
rect 21376 12764 21404 12792
rect 22186 12764 22192 12776
rect 21376 12736 22192 12764
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 23658 12724 23664 12776
rect 23716 12724 23722 12776
rect 25222 12724 25228 12776
rect 25280 12764 25286 12776
rect 25424 12773 25452 12804
rect 26697 12801 26709 12835
rect 26743 12832 26755 12835
rect 27246 12832 27252 12844
rect 26743 12804 27252 12832
rect 26743 12801 26755 12804
rect 26697 12795 26755 12801
rect 27246 12792 27252 12804
rect 27304 12792 27310 12844
rect 27448 12841 27476 12872
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12832 27491 12835
rect 27522 12832 27528 12844
rect 27479 12804 27528 12832
rect 27479 12801 27491 12804
rect 27433 12795 27491 12801
rect 27522 12792 27528 12804
rect 27580 12792 27586 12844
rect 27706 12792 27712 12844
rect 27764 12832 27770 12844
rect 28184 12832 28212 12928
rect 28721 12903 28779 12909
rect 28721 12869 28733 12903
rect 28767 12900 28779 12903
rect 29454 12900 29460 12912
rect 28767 12872 29460 12900
rect 28767 12869 28779 12872
rect 28721 12863 28779 12869
rect 29454 12860 29460 12872
rect 29512 12860 29518 12912
rect 31757 12903 31815 12909
rect 31757 12869 31769 12903
rect 31803 12900 31815 12903
rect 32401 12903 32459 12909
rect 32401 12900 32413 12903
rect 31803 12872 32413 12900
rect 31803 12869 31815 12872
rect 31757 12863 31815 12869
rect 32401 12869 32413 12872
rect 32447 12869 32459 12903
rect 32401 12863 32459 12869
rect 32585 12903 32643 12909
rect 32585 12869 32597 12903
rect 32631 12900 32643 12903
rect 33042 12900 33048 12912
rect 32631 12872 33048 12900
rect 32631 12869 32643 12872
rect 32585 12863 32643 12869
rect 27764 12804 28212 12832
rect 29472 12832 29500 12860
rect 30380 12835 30438 12841
rect 30380 12832 30392 12835
rect 29472 12804 30392 12832
rect 27764 12792 27770 12804
rect 30380 12801 30392 12804
rect 30426 12801 30438 12835
rect 30380 12795 30438 12801
rect 25409 12767 25467 12773
rect 25409 12764 25421 12767
rect 25280 12736 25421 12764
rect 25280 12724 25286 12736
rect 25409 12733 25421 12736
rect 25455 12733 25467 12767
rect 29914 12764 29920 12776
rect 29875 12736 29920 12764
rect 25409 12727 25467 12733
rect 29914 12724 29920 12736
rect 29972 12724 29978 12776
rect 30282 12724 30288 12776
rect 30340 12764 30346 12776
rect 30653 12767 30711 12773
rect 30653 12764 30665 12767
rect 30340 12736 30665 12764
rect 30340 12724 30346 12736
rect 30653 12733 30665 12736
rect 30699 12733 30711 12767
rect 32416 12764 32444 12863
rect 33042 12860 33048 12872
rect 33100 12860 33106 12912
rect 33152 12841 33180 12940
rect 34698 12928 34704 12940
rect 34756 12928 34762 12980
rect 36446 12928 36452 12980
rect 36504 12968 36510 12980
rect 36814 12968 36820 12980
rect 36504 12940 36820 12968
rect 36504 12928 36510 12940
rect 36814 12928 36820 12940
rect 36872 12968 36878 12980
rect 36909 12971 36967 12977
rect 36909 12968 36921 12971
rect 36872 12940 36921 12968
rect 36872 12928 36878 12940
rect 36909 12937 36921 12940
rect 36955 12937 36967 12971
rect 37550 12968 37556 12980
rect 37511 12940 37556 12968
rect 36909 12931 36967 12937
rect 37550 12928 37556 12940
rect 37608 12928 37614 12980
rect 33137 12835 33195 12841
rect 33137 12801 33149 12835
rect 33183 12832 33195 12835
rect 33597 12835 33655 12841
rect 33597 12832 33609 12835
rect 33183 12804 33609 12832
rect 33183 12801 33195 12804
rect 33137 12795 33195 12801
rect 33597 12801 33609 12804
rect 33643 12832 33655 12835
rect 33686 12832 33692 12844
rect 33643 12804 33692 12832
rect 33643 12801 33655 12804
rect 33597 12795 33655 12801
rect 33686 12792 33692 12804
rect 33744 12792 33750 12844
rect 34716 12832 34744 12928
rect 36538 12900 36544 12912
rect 36499 12872 36544 12900
rect 36538 12860 36544 12872
rect 36596 12860 36602 12912
rect 36556 12832 36584 12860
rect 37093 12835 37151 12841
rect 37093 12832 37105 12835
rect 34716 12804 35020 12832
rect 36556 12804 37105 12832
rect 33045 12767 33103 12773
rect 33045 12764 33057 12767
rect 32416 12736 33057 12764
rect 30653 12727 30711 12733
rect 33045 12733 33057 12736
rect 33091 12764 33103 12767
rect 33410 12764 33416 12776
rect 33091 12736 33416 12764
rect 33091 12733 33103 12736
rect 33045 12727 33103 12733
rect 33410 12724 33416 12736
rect 33468 12724 33474 12776
rect 33502 12724 33508 12776
rect 33560 12764 33566 12776
rect 34057 12767 34115 12773
rect 34057 12764 34069 12767
rect 33560 12736 34069 12764
rect 33560 12724 33566 12736
rect 34057 12733 34069 12736
rect 34103 12764 34115 12767
rect 34885 12767 34943 12773
rect 34885 12764 34897 12767
rect 34103 12736 34897 12764
rect 34103 12733 34115 12736
rect 34057 12727 34115 12733
rect 34885 12733 34897 12736
rect 34931 12733 34943 12767
rect 34992 12764 35020 12804
rect 37093 12801 37105 12804
rect 37139 12801 37151 12835
rect 37093 12795 37151 12801
rect 35141 12767 35199 12773
rect 35141 12764 35153 12767
rect 34992 12736 35153 12764
rect 34885 12727 34943 12733
rect 35141 12733 35153 12736
rect 35187 12733 35199 12767
rect 35141 12727 35199 12733
rect 21450 12656 21456 12708
rect 21508 12696 21514 12708
rect 21606 12699 21664 12705
rect 21606 12696 21618 12699
rect 21508 12668 21618 12696
rect 21508 12656 21514 12668
rect 21606 12665 21618 12668
rect 21652 12665 21664 12699
rect 21606 12659 21664 12665
rect 23477 12699 23535 12705
rect 23477 12665 23489 12699
rect 23523 12696 23535 12699
rect 23676 12696 23704 12724
rect 24121 12699 24179 12705
rect 24121 12696 24133 12699
rect 23523 12668 24133 12696
rect 23523 12665 23535 12668
rect 23477 12659 23535 12665
rect 24121 12665 24133 12668
rect 24167 12665 24179 12699
rect 24121 12659 24179 12665
rect 24210 12656 24216 12708
rect 24268 12696 24274 12708
rect 25314 12696 25320 12708
rect 24268 12668 25320 12696
rect 24268 12656 24274 12668
rect 25314 12656 25320 12668
rect 25372 12696 25378 12708
rect 25685 12699 25743 12705
rect 25685 12696 25697 12699
rect 25372 12668 25697 12696
rect 25372 12656 25378 12668
rect 25685 12665 25697 12668
rect 25731 12665 25743 12699
rect 32950 12696 32956 12708
rect 32911 12668 32956 12696
rect 25685 12659 25743 12665
rect 32950 12656 32956 12668
rect 33008 12656 33014 12708
rect 34900 12696 34928 12727
rect 35342 12696 35348 12708
rect 34900 12668 35348 12696
rect 35342 12656 35348 12668
rect 35400 12656 35406 12708
rect 24026 12628 24032 12640
rect 23987 12600 24032 12628
rect 24026 12588 24032 12600
rect 24084 12588 24090 12640
rect 25225 12631 25283 12637
rect 25225 12597 25237 12631
rect 25271 12628 25283 12631
rect 25866 12628 25872 12640
rect 25271 12600 25872 12628
rect 25271 12597 25283 12600
rect 25225 12591 25283 12597
rect 25866 12588 25872 12600
rect 25924 12588 25930 12640
rect 26970 12588 26976 12640
rect 27028 12628 27034 12640
rect 27157 12631 27215 12637
rect 27157 12628 27169 12631
rect 27028 12600 27169 12628
rect 27028 12588 27034 12600
rect 27157 12597 27169 12600
rect 27203 12597 27215 12631
rect 27157 12591 27215 12597
rect 29825 12631 29883 12637
rect 29825 12597 29837 12631
rect 29871 12628 29883 12631
rect 30383 12631 30441 12637
rect 30383 12628 30395 12631
rect 29871 12600 30395 12628
rect 29871 12597 29883 12600
rect 29825 12591 29883 12597
rect 30383 12597 30395 12600
rect 30429 12628 30441 12631
rect 31294 12628 31300 12640
rect 30429 12600 31300 12628
rect 30429 12597 30441 12600
rect 30383 12591 30441 12597
rect 31294 12588 31300 12600
rect 31352 12588 31358 12640
rect 35986 12588 35992 12640
rect 36044 12628 36050 12640
rect 36265 12631 36323 12637
rect 36265 12628 36277 12631
rect 36044 12600 36277 12628
rect 36044 12588 36050 12600
rect 36265 12597 36277 12600
rect 36311 12597 36323 12631
rect 36265 12591 36323 12597
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 21450 12424 21456 12436
rect 21411 12396 21456 12424
rect 21450 12384 21456 12396
rect 21508 12424 21514 12436
rect 23385 12427 23443 12433
rect 23385 12424 23397 12427
rect 21508 12396 23397 12424
rect 21508 12384 21514 12396
rect 23385 12393 23397 12396
rect 23431 12424 23443 12427
rect 23661 12427 23719 12433
rect 23661 12424 23673 12427
rect 23431 12396 23673 12424
rect 23431 12393 23443 12396
rect 23385 12387 23443 12393
rect 23661 12393 23673 12396
rect 23707 12424 23719 12427
rect 23842 12424 23848 12436
rect 23707 12396 23848 12424
rect 23707 12393 23719 12396
rect 23661 12387 23719 12393
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 24026 12424 24032 12436
rect 23987 12396 24032 12424
rect 24026 12384 24032 12396
rect 24084 12384 24090 12436
rect 24210 12424 24216 12436
rect 24171 12396 24216 12424
rect 24210 12384 24216 12396
rect 24268 12384 24274 12436
rect 25222 12424 25228 12436
rect 25183 12396 25228 12424
rect 25222 12384 25228 12396
rect 25280 12384 25286 12436
rect 27706 12384 27712 12436
rect 27764 12424 27770 12436
rect 28721 12427 28779 12433
rect 28721 12424 28733 12427
rect 27764 12396 28733 12424
rect 27764 12384 27770 12396
rect 28721 12393 28733 12396
rect 28767 12393 28779 12427
rect 29178 12424 29184 12436
rect 29139 12396 29184 12424
rect 28721 12387 28779 12393
rect 29178 12384 29184 12396
rect 29236 12384 29242 12436
rect 29546 12424 29552 12436
rect 29459 12396 29552 12424
rect 29546 12384 29552 12396
rect 29604 12424 29610 12436
rect 30006 12424 30012 12436
rect 29604 12396 30012 12424
rect 29604 12384 29610 12396
rect 30006 12384 30012 12396
rect 30064 12384 30070 12436
rect 31110 12424 31116 12436
rect 31071 12396 31116 12424
rect 31110 12384 31116 12396
rect 31168 12384 31174 12436
rect 34238 12384 34244 12436
rect 34296 12424 34302 12436
rect 34698 12424 34704 12436
rect 34296 12396 34704 12424
rect 34296 12384 34302 12396
rect 34698 12384 34704 12396
rect 34756 12384 34762 12436
rect 36814 12424 36820 12436
rect 36775 12396 36820 12424
rect 36814 12384 36820 12396
rect 36872 12384 36878 12436
rect 27249 12359 27307 12365
rect 27249 12325 27261 12359
rect 27295 12356 27307 12359
rect 27338 12356 27344 12368
rect 27295 12328 27344 12356
rect 27295 12325 27307 12328
rect 27249 12319 27307 12325
rect 27338 12316 27344 12328
rect 27396 12356 27402 12368
rect 27890 12356 27896 12368
rect 27396 12328 27896 12356
rect 27396 12316 27402 12328
rect 27890 12316 27896 12328
rect 27948 12316 27954 12368
rect 35345 12359 35403 12365
rect 35345 12325 35357 12359
rect 35391 12356 35403 12359
rect 35704 12359 35762 12365
rect 35704 12356 35716 12359
rect 35391 12328 35716 12356
rect 35391 12325 35403 12328
rect 35345 12319 35403 12325
rect 35704 12325 35716 12328
rect 35750 12356 35762 12359
rect 35986 12356 35992 12368
rect 35750 12328 35992 12356
rect 35750 12325 35762 12328
rect 35704 12319 35762 12325
rect 35986 12316 35992 12328
rect 36044 12316 36050 12368
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22261 12291 22319 12297
rect 22261 12288 22273 12291
rect 22152 12260 22273 12288
rect 22152 12248 22158 12260
rect 22261 12257 22273 12260
rect 22307 12257 22319 12291
rect 24578 12288 24584 12300
rect 24539 12260 24584 12288
rect 22261 12251 22319 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 27614 12297 27620 12300
rect 27608 12288 27620 12297
rect 27575 12260 27620 12288
rect 27608 12251 27620 12260
rect 27614 12248 27620 12251
rect 27672 12248 27678 12300
rect 30006 12297 30012 12300
rect 30000 12288 30012 12297
rect 29967 12260 30012 12288
rect 30000 12251 30012 12260
rect 30006 12248 30012 12251
rect 30064 12248 30070 12300
rect 32398 12248 32404 12300
rect 32456 12288 32462 12300
rect 33092 12291 33150 12297
rect 33092 12288 33104 12291
rect 32456 12260 33104 12288
rect 32456 12248 32462 12260
rect 33092 12257 33104 12260
rect 33138 12257 33150 12291
rect 34238 12288 34244 12300
rect 33092 12251 33150 12257
rect 33336 12260 34244 12288
rect 22005 12223 22063 12229
rect 22005 12189 22017 12223
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 21821 12087 21879 12093
rect 21821 12053 21833 12087
rect 21867 12084 21879 12087
rect 22020 12084 22048 12183
rect 24486 12180 24492 12232
rect 24544 12220 24550 12232
rect 24673 12223 24731 12229
rect 24673 12220 24685 12223
rect 24544 12192 24685 12220
rect 24544 12180 24550 12192
rect 24673 12189 24685 12192
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 24762 12180 24768 12232
rect 24820 12220 24826 12232
rect 24820 12192 24913 12220
rect 24820 12180 24826 12192
rect 26694 12180 26700 12232
rect 26752 12220 26758 12232
rect 27341 12223 27399 12229
rect 27341 12220 27353 12223
rect 26752 12192 27353 12220
rect 26752 12180 26758 12192
rect 27341 12189 27353 12192
rect 27387 12189 27399 12223
rect 27341 12183 27399 12189
rect 29733 12223 29791 12229
rect 29733 12189 29745 12223
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 24302 12112 24308 12164
rect 24360 12152 24366 12164
rect 24780 12152 24808 12180
rect 24360 12124 24808 12152
rect 24360 12112 24366 12124
rect 22186 12084 22192 12096
rect 21867 12056 22192 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 26881 12087 26939 12093
rect 26881 12053 26893 12087
rect 26927 12084 26939 12087
rect 26970 12084 26976 12096
rect 26927 12056 26976 12084
rect 26927 12053 26939 12056
rect 26881 12047 26939 12053
rect 26970 12044 26976 12056
rect 27028 12044 27034 12096
rect 29748 12084 29776 12183
rect 31018 12180 31024 12232
rect 31076 12220 31082 12232
rect 31938 12220 31944 12232
rect 31076 12192 31944 12220
rect 31076 12180 31082 12192
rect 31938 12180 31944 12192
rect 31996 12220 32002 12232
rect 32769 12223 32827 12229
rect 32769 12220 32781 12223
rect 31996 12192 32781 12220
rect 31996 12180 32002 12192
rect 32769 12189 32781 12192
rect 32815 12189 32827 12223
rect 32769 12183 32827 12189
rect 33226 12180 33232 12232
rect 33284 12220 33290 12232
rect 33336 12220 33364 12260
rect 34238 12248 34244 12260
rect 34296 12288 34302 12300
rect 34885 12291 34943 12297
rect 34885 12288 34897 12291
rect 34296 12260 34897 12288
rect 34296 12248 34302 12260
rect 34885 12257 34897 12260
rect 34931 12257 34943 12291
rect 34885 12251 34943 12257
rect 35437 12291 35495 12297
rect 35437 12257 35449 12291
rect 35483 12288 35495 12291
rect 36262 12288 36268 12300
rect 35483 12260 36268 12288
rect 35483 12257 35495 12260
rect 35437 12251 35495 12257
rect 33284 12192 33364 12220
rect 33284 12180 33290 12192
rect 33410 12180 33416 12232
rect 33468 12220 33474 12232
rect 33505 12223 33563 12229
rect 33505 12220 33517 12223
rect 33468 12192 33517 12220
rect 33468 12180 33474 12192
rect 33505 12189 33517 12192
rect 33551 12220 33563 12223
rect 34146 12220 34152 12232
rect 33551 12192 34152 12220
rect 33551 12189 33563 12192
rect 33505 12183 33563 12189
rect 34146 12180 34152 12192
rect 34204 12180 34210 12232
rect 34900 12220 34928 12251
rect 36262 12248 36268 12260
rect 36320 12248 36326 12300
rect 35250 12220 35256 12232
rect 34900 12192 35256 12220
rect 35250 12180 35256 12192
rect 35308 12180 35314 12232
rect 31941 12087 31999 12093
rect 31941 12084 31953 12087
rect 29748 12056 31953 12084
rect 31941 12053 31953 12056
rect 31987 12084 31999 12087
rect 32030 12084 32036 12096
rect 31987 12056 32036 12084
rect 31987 12053 31999 12056
rect 31941 12047 31999 12053
rect 32030 12044 32036 12056
rect 32088 12044 32094 12096
rect 32490 12084 32496 12096
rect 32451 12056 32496 12084
rect 32490 12044 32496 12056
rect 32548 12044 32554 12096
rect 32582 12044 32588 12096
rect 32640 12084 32646 12096
rect 34609 12087 34667 12093
rect 34609 12084 34621 12087
rect 32640 12056 34621 12084
rect 32640 12044 32646 12056
rect 34609 12053 34621 12056
rect 34655 12084 34667 12087
rect 34790 12084 34796 12096
rect 34655 12056 34796 12084
rect 34655 12053 34667 12056
rect 34609 12047 34667 12053
rect 34790 12044 34796 12056
rect 34848 12044 34854 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 23382 11880 23388 11892
rect 22152 11852 23388 11880
rect 22152 11840 22158 11852
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 23658 11880 23664 11892
rect 23619 11852 23664 11880
rect 23658 11840 23664 11852
rect 23716 11840 23722 11892
rect 24578 11840 24584 11892
rect 24636 11880 24642 11892
rect 25041 11883 25099 11889
rect 25041 11880 25053 11883
rect 24636 11852 25053 11880
rect 24636 11840 24642 11852
rect 25041 11849 25053 11852
rect 25087 11849 25099 11883
rect 25041 11843 25099 11849
rect 26605 11883 26663 11889
rect 26605 11849 26617 11883
rect 26651 11880 26663 11883
rect 27614 11880 27620 11892
rect 26651 11852 27620 11880
rect 26651 11849 26663 11852
rect 26605 11843 26663 11849
rect 27614 11840 27620 11852
rect 27672 11840 27678 11892
rect 29546 11840 29552 11892
rect 29604 11880 29610 11892
rect 30653 11883 30711 11889
rect 30653 11880 30665 11883
rect 29604 11852 30665 11880
rect 29604 11840 29610 11852
rect 30653 11849 30665 11852
rect 30699 11849 30711 11883
rect 32398 11880 32404 11892
rect 32359 11852 32404 11880
rect 30653 11843 30711 11849
rect 32398 11840 32404 11852
rect 32456 11840 32462 11892
rect 33502 11880 33508 11892
rect 32511 11852 33508 11880
rect 31389 11815 31447 11821
rect 31389 11781 31401 11815
rect 31435 11812 31447 11815
rect 32030 11812 32036 11824
rect 31435 11784 32036 11812
rect 31435 11781 31447 11784
rect 31389 11775 31447 11781
rect 32030 11772 32036 11784
rect 32088 11812 32094 11824
rect 32511 11812 32539 11852
rect 33502 11840 33508 11852
rect 33560 11840 33566 11892
rect 33686 11840 33692 11892
rect 33744 11880 33750 11892
rect 33873 11883 33931 11889
rect 33873 11880 33885 11883
rect 33744 11852 33885 11880
rect 33744 11840 33750 11852
rect 33873 11849 33885 11852
rect 33919 11849 33931 11883
rect 34146 11880 34152 11892
rect 34107 11852 34152 11880
rect 33873 11843 33931 11849
rect 34146 11840 34152 11852
rect 34204 11840 34210 11892
rect 35986 11880 35992 11892
rect 35947 11852 35992 11880
rect 35986 11840 35992 11852
rect 36044 11840 36050 11892
rect 36262 11880 36268 11892
rect 36223 11852 36268 11880
rect 36262 11840 36268 11852
rect 36320 11840 36326 11892
rect 32088 11784 32539 11812
rect 32088 11772 32094 11784
rect 23109 11747 23167 11753
rect 23109 11713 23121 11747
rect 23155 11744 23167 11747
rect 24210 11744 24216 11756
rect 23155 11716 24216 11744
rect 23155 11713 23167 11716
rect 23109 11707 23167 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 32511 11753 32539 11784
rect 34609 11815 34667 11821
rect 34609 11781 34621 11815
rect 34655 11812 34667 11815
rect 34790 11812 34796 11824
rect 34655 11784 34796 11812
rect 34655 11781 34667 11784
rect 34609 11775 34667 11781
rect 34790 11772 34796 11784
rect 34848 11812 34854 11824
rect 34848 11784 35388 11812
rect 34848 11772 34854 11784
rect 28721 11747 28779 11753
rect 28721 11713 28733 11747
rect 28767 11744 28779 11747
rect 32493 11747 32551 11753
rect 28767 11716 29408 11744
rect 28767 11713 28779 11716
rect 28721 11707 28779 11713
rect 23842 11636 23848 11688
rect 23900 11676 23906 11688
rect 24029 11679 24087 11685
rect 24029 11676 24041 11679
rect 23900 11648 24041 11676
rect 23900 11636 23906 11648
rect 24029 11645 24041 11648
rect 24075 11645 24087 11679
rect 24029 11639 24087 11645
rect 25869 11679 25927 11685
rect 25869 11645 25881 11679
rect 25915 11676 25927 11679
rect 26237 11679 26295 11685
rect 26237 11676 26249 11679
rect 25915 11648 26249 11676
rect 25915 11645 25927 11648
rect 25869 11639 25927 11645
rect 26237 11645 26249 11648
rect 26283 11676 26295 11679
rect 26694 11676 26700 11688
rect 26283 11648 26700 11676
rect 26283 11645 26295 11648
rect 26237 11639 26295 11645
rect 26694 11636 26700 11648
rect 26752 11636 26758 11688
rect 29270 11676 29276 11688
rect 29231 11648 29276 11676
rect 29270 11636 29276 11648
rect 29328 11636 29334 11688
rect 29380 11676 29408 11716
rect 32493 11713 32505 11747
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 33962 11704 33968 11756
rect 34020 11744 34026 11756
rect 34146 11744 34152 11756
rect 34020 11716 34152 11744
rect 34020 11704 34026 11716
rect 34146 11704 34152 11716
rect 34204 11704 34210 11756
rect 35360 11753 35388 11784
rect 35345 11747 35403 11753
rect 35345 11713 35357 11747
rect 35391 11713 35403 11747
rect 35345 11707 35403 11713
rect 35529 11747 35587 11753
rect 35529 11713 35541 11747
rect 35575 11744 35587 11747
rect 36004 11744 36032 11840
rect 35575 11716 36032 11744
rect 35575 11713 35587 11716
rect 35529 11707 35587 11713
rect 29540 11679 29598 11685
rect 29540 11676 29552 11679
rect 29380 11648 29552 11676
rect 29540 11645 29552 11648
rect 29586 11676 29598 11679
rect 31110 11676 31116 11688
rect 29586 11648 31116 11676
rect 29586 11645 29598 11648
rect 29540 11639 29598 11645
rect 31110 11636 31116 11648
rect 31168 11636 31174 11688
rect 32033 11679 32091 11685
rect 32033 11645 32045 11679
rect 32079 11676 32091 11679
rect 33226 11676 33232 11688
rect 32079 11648 33232 11676
rect 32079 11645 32091 11648
rect 32033 11639 32091 11645
rect 33226 11636 33232 11648
rect 33284 11636 33290 11688
rect 35250 11676 35256 11688
rect 35211 11648 35256 11676
rect 35250 11636 35256 11648
rect 35308 11636 35314 11688
rect 36446 11676 36452 11688
rect 36359 11648 36452 11676
rect 36446 11636 36452 11648
rect 36504 11676 36510 11688
rect 37001 11679 37059 11685
rect 37001 11676 37013 11679
rect 36504 11648 37013 11676
rect 36504 11636 36510 11648
rect 37001 11645 37013 11648
rect 37047 11645 37059 11679
rect 37001 11639 37059 11645
rect 23382 11568 23388 11620
rect 23440 11608 23446 11620
rect 24121 11611 24179 11617
rect 24121 11608 24133 11611
rect 23440 11580 24133 11608
rect 23440 11568 23446 11580
rect 24121 11577 24133 11580
rect 24167 11577 24179 11611
rect 24121 11571 24179 11577
rect 26878 11568 26884 11620
rect 26936 11617 26942 11620
rect 26936 11611 27000 11617
rect 26936 11577 26954 11611
rect 26988 11577 27000 11611
rect 29288 11608 29316 11636
rect 30929 11611 30987 11617
rect 30929 11608 30941 11611
rect 29288 11580 30941 11608
rect 26936 11571 27000 11577
rect 30929 11577 30941 11580
rect 30975 11577 30987 11611
rect 30929 11571 30987 11577
rect 26936 11568 26942 11571
rect 31662 11568 31668 11620
rect 31720 11608 31726 11620
rect 32398 11608 32404 11620
rect 31720 11580 32404 11608
rect 31720 11568 31726 11580
rect 32398 11568 32404 11580
rect 32456 11568 32462 11620
rect 32490 11568 32496 11620
rect 32548 11608 32554 11620
rect 32738 11611 32796 11617
rect 32738 11608 32750 11611
rect 32548 11580 32750 11608
rect 32548 11568 32554 11580
rect 32738 11577 32750 11580
rect 32784 11577 32796 11611
rect 35710 11608 35716 11620
rect 32738 11571 32796 11577
rect 34900 11580 35716 11608
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 22373 11543 22431 11549
rect 22373 11540 22385 11543
rect 22244 11512 22385 11540
rect 22244 11500 22250 11512
rect 22373 11509 22385 11512
rect 22419 11509 22431 11543
rect 22373 11503 22431 11509
rect 24486 11500 24492 11552
rect 24544 11540 24550 11552
rect 24670 11540 24676 11552
rect 24544 11512 24676 11540
rect 24544 11500 24550 11512
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 27614 11500 27620 11552
rect 27672 11540 27678 11552
rect 28077 11543 28135 11549
rect 28077 11540 28089 11543
rect 27672 11512 28089 11540
rect 27672 11500 27678 11512
rect 28077 11509 28089 11512
rect 28123 11509 28135 11543
rect 28077 11503 28135 11509
rect 29089 11543 29147 11549
rect 29089 11509 29101 11543
rect 29135 11540 29147 11543
rect 30006 11540 30012 11552
rect 29135 11512 30012 11540
rect 29135 11509 29147 11512
rect 29089 11503 29147 11509
rect 30006 11500 30012 11512
rect 30064 11500 30070 11552
rect 31481 11543 31539 11549
rect 31481 11509 31493 11543
rect 31527 11540 31539 11543
rect 31754 11540 31760 11552
rect 31527 11512 31760 11540
rect 31527 11509 31539 11512
rect 31481 11503 31539 11509
rect 31754 11500 31760 11512
rect 31812 11500 31818 11552
rect 34900 11549 34928 11580
rect 35710 11568 35716 11580
rect 35768 11568 35774 11620
rect 34885 11543 34943 11549
rect 34885 11509 34897 11543
rect 34931 11509 34943 11543
rect 36630 11540 36636 11552
rect 36591 11512 36636 11540
rect 34885 11503 34943 11509
rect 36630 11500 36636 11512
rect 36688 11500 36694 11552
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 23382 11296 23388 11348
rect 23440 11336 23446 11348
rect 23569 11339 23627 11345
rect 23569 11336 23581 11339
rect 23440 11308 23581 11336
rect 23440 11296 23446 11308
rect 23569 11305 23581 11308
rect 23615 11305 23627 11339
rect 24302 11336 24308 11348
rect 24263 11308 24308 11336
rect 23569 11299 23627 11305
rect 24302 11296 24308 11308
rect 24360 11296 24366 11348
rect 24397 11339 24455 11345
rect 24397 11305 24409 11339
rect 24443 11336 24455 11339
rect 24578 11336 24584 11348
rect 24443 11308 24584 11336
rect 24443 11305 24455 11308
rect 24397 11299 24455 11305
rect 24578 11296 24584 11308
rect 24636 11296 24642 11348
rect 30374 11296 30380 11348
rect 30432 11336 30438 11348
rect 30653 11339 30711 11345
rect 30653 11336 30665 11339
rect 30432 11308 30665 11336
rect 30432 11296 30438 11308
rect 30653 11305 30665 11308
rect 30699 11305 30711 11339
rect 31938 11336 31944 11348
rect 31899 11308 31944 11336
rect 30653 11299 30711 11305
rect 31938 11296 31944 11308
rect 31996 11296 32002 11348
rect 32490 11296 32496 11348
rect 32548 11336 32554 11348
rect 33505 11339 33563 11345
rect 33505 11336 33517 11339
rect 32548 11308 33517 11336
rect 32548 11296 32554 11308
rect 33505 11305 33517 11308
rect 33551 11305 33563 11339
rect 33505 11299 33563 11305
rect 34422 11296 34428 11348
rect 34480 11336 34486 11348
rect 34885 11339 34943 11345
rect 34885 11336 34897 11339
rect 34480 11308 34897 11336
rect 34480 11296 34486 11308
rect 34885 11305 34897 11308
rect 34931 11305 34943 11339
rect 36446 11336 36452 11348
rect 36407 11308 36452 11336
rect 34885 11299 34943 11305
rect 36446 11296 36452 11308
rect 36504 11296 36510 11348
rect 24210 11228 24216 11280
rect 24268 11268 24274 11280
rect 27332 11271 27390 11277
rect 24268 11240 25084 11268
rect 24268 11228 24274 11240
rect 22278 11160 22284 11212
rect 22336 11200 22342 11212
rect 22445 11203 22503 11209
rect 22445 11200 22457 11203
rect 22336 11172 22457 11200
rect 22336 11160 22342 11172
rect 22445 11169 22457 11172
rect 22491 11169 22503 11203
rect 24762 11200 24768 11212
rect 24723 11172 24768 11200
rect 22445 11163 22503 11169
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 22186 11132 22192 11144
rect 22147 11104 22192 11132
rect 22186 11092 22192 11104
rect 22244 11092 22250 11144
rect 25056 11141 25084 11240
rect 27332 11237 27344 11271
rect 27378 11268 27390 11271
rect 27706 11268 27712 11280
rect 27378 11240 27712 11268
rect 27378 11237 27390 11240
rect 27332 11231 27390 11237
rect 27706 11228 27712 11240
rect 27764 11228 27770 11280
rect 29546 11277 29552 11280
rect 29540 11268 29552 11277
rect 29507 11240 29552 11268
rect 29540 11231 29552 11240
rect 29546 11228 29552 11231
rect 29604 11228 29610 11280
rect 33134 11228 33140 11280
rect 33192 11268 33198 11280
rect 34333 11271 34391 11277
rect 34333 11268 34345 11271
rect 33192 11240 34345 11268
rect 33192 11228 33198 11240
rect 34333 11237 34345 11240
rect 34379 11268 34391 11271
rect 34977 11271 35035 11277
rect 34977 11268 34989 11271
rect 34379 11240 34989 11268
rect 34379 11237 34391 11240
rect 34333 11231 34391 11237
rect 34977 11237 34989 11240
rect 35023 11237 35035 11271
rect 36078 11268 36084 11280
rect 36039 11240 36084 11268
rect 34977 11231 35035 11237
rect 36078 11228 36084 11240
rect 36136 11228 36142 11280
rect 26694 11160 26700 11212
rect 26752 11200 26758 11212
rect 27065 11203 27123 11209
rect 27065 11200 27077 11203
rect 26752 11172 27077 11200
rect 26752 11160 26758 11172
rect 27065 11169 27077 11172
rect 27111 11200 27123 11203
rect 32392 11203 32450 11209
rect 27111 11172 28764 11200
rect 27111 11169 27123 11172
rect 27065 11163 27123 11169
rect 28736 11144 28764 11172
rect 32392 11169 32404 11203
rect 32438 11200 32450 11203
rect 32674 11200 32680 11212
rect 32438 11172 32680 11200
rect 32438 11169 32450 11172
rect 32392 11163 32450 11169
rect 32674 11160 32680 11172
rect 32732 11160 32738 11212
rect 34606 11160 34612 11212
rect 34664 11200 34670 11212
rect 34664 11172 35112 11200
rect 34664 11160 34670 11172
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 25041 11135 25099 11141
rect 25041 11101 25053 11135
rect 25087 11132 25099 11135
rect 25087 11104 25176 11132
rect 25087 11101 25099 11104
rect 25041 11095 25099 11101
rect 24872 10996 24900 11095
rect 25038 10996 25044 11008
rect 24872 10968 25044 10996
rect 25038 10956 25044 10968
rect 25096 10956 25102 11008
rect 25148 10996 25176 11104
rect 28718 11092 28724 11144
rect 28776 11132 28782 11144
rect 29270 11132 29276 11144
rect 28776 11104 29276 11132
rect 28776 11092 28782 11104
rect 29270 11092 29276 11104
rect 29328 11092 29334 11144
rect 31478 11092 31484 11144
rect 31536 11132 31542 11144
rect 35084 11141 35112 11172
rect 36170 11160 36176 11212
rect 36228 11200 36234 11212
rect 36265 11203 36323 11209
rect 36265 11200 36277 11203
rect 36228 11172 36277 11200
rect 36228 11160 36234 11172
rect 36265 11169 36277 11172
rect 36311 11169 36323 11203
rect 36265 11163 36323 11169
rect 32125 11135 32183 11141
rect 32125 11132 32137 11135
rect 31536 11104 32137 11132
rect 31536 11092 31542 11104
rect 32125 11101 32137 11104
rect 32171 11101 32183 11135
rect 32125 11095 32183 11101
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11101 35127 11135
rect 35069 11095 35127 11101
rect 28445 11067 28503 11073
rect 28445 11064 28457 11067
rect 28000 11036 28457 11064
rect 25406 10996 25412 11008
rect 25148 10968 25412 10996
rect 25406 10956 25412 10968
rect 25464 10956 25470 11008
rect 26789 10999 26847 11005
rect 26789 10965 26801 10999
rect 26835 10996 26847 10999
rect 26878 10996 26884 11008
rect 26835 10968 26884 10996
rect 26835 10965 26847 10968
rect 26789 10959 26847 10965
rect 26878 10956 26884 10968
rect 26936 10996 26942 11008
rect 27430 10996 27436 11008
rect 26936 10968 27436 10996
rect 26936 10956 26942 10968
rect 27430 10956 27436 10968
rect 27488 10996 27494 11008
rect 28000 10996 28028 11036
rect 28445 11033 28457 11036
rect 28491 11033 28503 11067
rect 34514 11064 34520 11076
rect 34475 11036 34520 11064
rect 28445 11027 28503 11033
rect 34514 11024 34520 11036
rect 34572 11024 34578 11076
rect 27488 10968 28028 10996
rect 35621 10999 35679 11005
rect 27488 10956 27494 10968
rect 35621 10965 35633 10999
rect 35667 10996 35679 10999
rect 35986 10996 35992 11008
rect 35667 10968 35992 10996
rect 35667 10965 35679 10968
rect 35621 10959 35679 10965
rect 35986 10956 35992 10968
rect 36044 10956 36050 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 22278 10792 22284 10804
rect 22239 10764 22284 10792
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 25406 10792 25412 10804
rect 25319 10764 25412 10792
rect 25406 10752 25412 10764
rect 25464 10792 25470 10804
rect 27338 10792 27344 10804
rect 25464 10764 27344 10792
rect 25464 10752 25470 10764
rect 27338 10752 27344 10764
rect 27396 10752 27402 10804
rect 27617 10795 27675 10801
rect 27617 10761 27629 10795
rect 27663 10792 27675 10795
rect 27706 10792 27712 10804
rect 27663 10764 27712 10792
rect 27663 10761 27675 10764
rect 27617 10755 27675 10761
rect 27706 10752 27712 10764
rect 27764 10752 27770 10804
rect 29546 10752 29552 10804
rect 29604 10792 29610 10804
rect 29917 10795 29975 10801
rect 29917 10792 29929 10795
rect 29604 10764 29929 10792
rect 29604 10752 29610 10764
rect 29917 10761 29929 10764
rect 29963 10761 29975 10795
rect 29917 10755 29975 10761
rect 31754 10752 31760 10804
rect 31812 10792 31818 10804
rect 31941 10795 31999 10801
rect 31812 10764 31857 10792
rect 31812 10752 31818 10764
rect 31941 10761 31953 10795
rect 31987 10792 31999 10795
rect 32950 10792 32956 10804
rect 31987 10764 32956 10792
rect 31987 10761 31999 10764
rect 31941 10755 31999 10761
rect 32950 10752 32956 10764
rect 33008 10752 33014 10804
rect 34422 10752 34428 10804
rect 34480 10792 34486 10804
rect 34517 10795 34575 10801
rect 34517 10792 34529 10795
rect 34480 10764 34529 10792
rect 34480 10752 34486 10764
rect 34517 10761 34529 10764
rect 34563 10761 34575 10795
rect 34517 10755 34575 10761
rect 29362 10616 29368 10668
rect 29420 10656 29426 10668
rect 29457 10659 29515 10665
rect 29457 10656 29469 10659
rect 29420 10628 29469 10656
rect 29420 10616 29426 10628
rect 29457 10625 29469 10628
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 31481 10659 31539 10665
rect 31481 10625 31493 10659
rect 31527 10656 31539 10659
rect 32490 10656 32496 10668
rect 31527 10628 32496 10656
rect 31527 10625 31539 10628
rect 31481 10619 31539 10625
rect 32490 10616 32496 10628
rect 32548 10616 32554 10668
rect 33042 10656 33048 10668
rect 33003 10628 33048 10656
rect 33042 10616 33048 10628
rect 33100 10616 33106 10668
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22649 10591 22707 10597
rect 22649 10588 22661 10591
rect 22244 10560 22661 10588
rect 22244 10548 22250 10560
rect 22649 10557 22661 10560
rect 22695 10588 22707 10591
rect 22738 10588 22744 10600
rect 22695 10560 22744 10588
rect 22695 10557 22707 10560
rect 22649 10551 22707 10557
rect 22738 10548 22744 10560
rect 22796 10588 22802 10600
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22796 10560 23121 10588
rect 22796 10548 22802 10560
rect 23109 10557 23121 10560
rect 23155 10588 23167 10591
rect 23661 10591 23719 10597
rect 23661 10588 23673 10591
rect 23155 10560 23673 10588
rect 23155 10557 23167 10560
rect 23109 10551 23167 10557
rect 23661 10557 23673 10560
rect 23707 10588 23719 10591
rect 23750 10588 23756 10600
rect 23707 10560 23756 10588
rect 23707 10557 23719 10560
rect 23661 10551 23719 10557
rect 23750 10548 23756 10560
rect 23808 10548 23814 10600
rect 25866 10588 25872 10600
rect 25827 10560 25872 10588
rect 25866 10548 25872 10560
rect 25924 10548 25930 10600
rect 30650 10588 30656 10600
rect 30611 10560 30656 10588
rect 30650 10548 30656 10560
rect 30708 10548 30714 10600
rect 30837 10591 30895 10597
rect 30837 10557 30849 10591
rect 30883 10588 30895 10591
rect 31202 10588 31208 10600
rect 30883 10560 31208 10588
rect 30883 10557 30895 10560
rect 30837 10551 30895 10557
rect 23477 10523 23535 10529
rect 23477 10489 23489 10523
rect 23523 10520 23535 10523
rect 23906 10523 23964 10529
rect 23906 10520 23918 10523
rect 23523 10492 23918 10520
rect 23523 10489 23535 10492
rect 23477 10483 23535 10489
rect 23906 10489 23918 10492
rect 23952 10520 23964 10523
rect 24486 10520 24492 10532
rect 23952 10492 24492 10520
rect 23952 10489 23964 10492
rect 23906 10483 23964 10489
rect 24486 10480 24492 10492
rect 24544 10480 24550 10532
rect 26142 10529 26148 10532
rect 25777 10523 25835 10529
rect 25777 10489 25789 10523
rect 25823 10520 25835 10523
rect 26136 10520 26148 10529
rect 25823 10492 26148 10520
rect 25823 10489 25835 10492
rect 25777 10483 25835 10489
rect 26136 10483 26148 10492
rect 26200 10520 26206 10532
rect 27522 10520 27528 10532
rect 26200 10492 27528 10520
rect 26142 10480 26148 10483
rect 26200 10480 26206 10492
rect 27522 10480 27528 10492
rect 27580 10480 27586 10532
rect 30377 10523 30435 10529
rect 30377 10489 30389 10523
rect 30423 10520 30435 10523
rect 30852 10520 30880 10551
rect 31202 10548 31208 10560
rect 31260 10548 31266 10600
rect 31754 10548 31760 10600
rect 31812 10588 31818 10600
rect 32309 10591 32367 10597
rect 32309 10588 32321 10591
rect 31812 10560 32321 10588
rect 31812 10548 31818 10560
rect 32309 10557 32321 10560
rect 32355 10557 32367 10591
rect 32309 10551 32367 10557
rect 33134 10548 33140 10600
rect 33192 10588 33198 10600
rect 33505 10591 33563 10597
rect 33505 10588 33517 10591
rect 33192 10560 33517 10588
rect 33192 10548 33198 10560
rect 33505 10557 33517 10560
rect 33551 10588 33563 10591
rect 34057 10591 34115 10597
rect 34057 10588 34069 10591
rect 33551 10560 34069 10588
rect 33551 10557 33563 10560
rect 33505 10551 33563 10557
rect 34057 10557 34069 10560
rect 34103 10557 34115 10591
rect 34057 10551 34115 10557
rect 35437 10591 35495 10597
rect 35437 10557 35449 10591
rect 35483 10588 35495 10591
rect 35986 10588 35992 10600
rect 35483 10560 35992 10588
rect 35483 10557 35495 10560
rect 35437 10551 35495 10557
rect 35986 10548 35992 10560
rect 36044 10548 36050 10600
rect 30423 10492 30880 10520
rect 30423 10489 30435 10492
rect 30377 10483 30435 10489
rect 32674 10480 32680 10532
rect 32732 10520 32738 10532
rect 33410 10520 33416 10532
rect 32732 10492 33416 10520
rect 32732 10480 32738 10492
rect 33410 10480 33416 10492
rect 33468 10520 33474 10532
rect 35345 10523 35403 10529
rect 33468 10492 33824 10520
rect 33468 10480 33474 10492
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 27246 10452 27252 10464
rect 27207 10424 27252 10452
rect 27246 10412 27252 10424
rect 27304 10412 27310 10464
rect 27985 10455 28043 10461
rect 27985 10421 27997 10455
rect 28031 10452 28043 10455
rect 28718 10452 28724 10464
rect 28031 10424 28724 10452
rect 28031 10421 28043 10424
rect 27985 10415 28043 10421
rect 28718 10412 28724 10424
rect 28776 10452 28782 10464
rect 28997 10455 29055 10461
rect 28997 10452 29009 10455
rect 28776 10424 29009 10452
rect 28776 10412 28782 10424
rect 28997 10421 29009 10424
rect 29043 10452 29055 10455
rect 30469 10455 30527 10461
rect 30469 10452 30481 10455
rect 29043 10424 30481 10452
rect 29043 10421 29055 10424
rect 28997 10415 29055 10421
rect 30469 10421 30481 10424
rect 30515 10452 30527 10455
rect 30834 10452 30840 10464
rect 30515 10424 30840 10452
rect 30515 10421 30527 10424
rect 30469 10415 30527 10421
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 31018 10452 31024 10464
rect 30979 10424 31024 10452
rect 31018 10412 31024 10424
rect 31076 10412 31082 10464
rect 32398 10412 32404 10464
rect 32456 10452 32462 10464
rect 33686 10452 33692 10464
rect 32456 10424 32501 10452
rect 33647 10424 33692 10452
rect 32456 10412 32462 10424
rect 33686 10412 33692 10424
rect 33744 10412 33750 10464
rect 33796 10452 33824 10492
rect 35345 10489 35357 10523
rect 35391 10520 35403 10523
rect 35704 10523 35762 10529
rect 35704 10520 35716 10523
rect 35391 10492 35716 10520
rect 35391 10489 35403 10492
rect 35345 10483 35403 10489
rect 35704 10489 35716 10492
rect 35750 10520 35762 10523
rect 36170 10520 36176 10532
rect 35750 10492 36176 10520
rect 35750 10489 35762 10492
rect 35704 10483 35762 10489
rect 36170 10480 36176 10492
rect 36228 10520 36234 10532
rect 36228 10492 37136 10520
rect 36228 10480 36234 10492
rect 37108 10464 37136 10492
rect 36817 10455 36875 10461
rect 36817 10452 36829 10455
rect 33796 10424 36829 10452
rect 36817 10421 36829 10424
rect 36863 10421 36875 10455
rect 37090 10452 37096 10464
rect 37051 10424 37096 10452
rect 36817 10415 36875 10421
rect 37090 10412 37096 10424
rect 37148 10412 37154 10464
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 22278 10208 22284 10260
rect 22336 10248 22342 10260
rect 24121 10251 24179 10257
rect 24121 10248 24133 10251
rect 22336 10220 24133 10248
rect 22336 10208 22342 10220
rect 24121 10217 24133 10220
rect 24167 10248 24179 10251
rect 24762 10248 24768 10260
rect 24167 10220 24768 10248
rect 24167 10217 24179 10220
rect 24121 10211 24179 10217
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 26970 10248 26976 10260
rect 26931 10220 26976 10248
rect 26970 10208 26976 10220
rect 27028 10208 27034 10260
rect 27341 10251 27399 10257
rect 27341 10217 27353 10251
rect 27387 10248 27399 10251
rect 27522 10248 27528 10260
rect 27387 10220 27528 10248
rect 27387 10217 27399 10220
rect 27341 10211 27399 10217
rect 27522 10208 27528 10220
rect 27580 10208 27586 10260
rect 30561 10251 30619 10257
rect 30561 10217 30573 10251
rect 30607 10248 30619 10251
rect 30650 10248 30656 10260
rect 30607 10220 30656 10248
rect 30607 10217 30619 10220
rect 30561 10211 30619 10217
rect 30650 10208 30656 10220
rect 30708 10208 30714 10260
rect 30834 10208 30840 10260
rect 30892 10248 30898 10260
rect 31478 10248 31484 10260
rect 30892 10220 31484 10248
rect 30892 10208 30898 10220
rect 31478 10208 31484 10220
rect 31536 10208 31542 10260
rect 31941 10251 31999 10257
rect 31941 10217 31953 10251
rect 31987 10248 31999 10251
rect 32398 10248 32404 10260
rect 31987 10220 32404 10248
rect 31987 10217 31999 10220
rect 31941 10211 31999 10217
rect 32398 10208 32404 10220
rect 32456 10208 32462 10260
rect 32582 10208 32588 10260
rect 32640 10248 32646 10260
rect 32861 10251 32919 10257
rect 32861 10248 32873 10251
rect 32640 10220 32873 10248
rect 32640 10208 32646 10220
rect 32861 10217 32873 10220
rect 32907 10248 32919 10251
rect 33686 10248 33692 10260
rect 32907 10220 33692 10248
rect 32907 10217 32919 10220
rect 32861 10211 32919 10217
rect 33686 10208 33692 10220
rect 33744 10208 33750 10260
rect 34149 10251 34207 10257
rect 34149 10217 34161 10251
rect 34195 10248 34207 10251
rect 34238 10248 34244 10260
rect 34195 10220 34244 10248
rect 34195 10217 34207 10220
rect 34149 10211 34207 10217
rect 34238 10208 34244 10220
rect 34296 10208 34302 10260
rect 34606 10248 34612 10260
rect 34567 10220 34612 10248
rect 34606 10208 34612 10220
rect 34664 10208 34670 10260
rect 35526 10208 35532 10260
rect 35584 10248 35590 10260
rect 35710 10248 35716 10260
rect 35584 10220 35716 10248
rect 35584 10208 35590 10220
rect 35710 10208 35716 10220
rect 35768 10208 35774 10260
rect 36078 10248 36084 10260
rect 36039 10220 36084 10248
rect 36078 10208 36084 10220
rect 36136 10208 36142 10260
rect 31018 10140 31024 10192
rect 31076 10180 31082 10192
rect 32490 10180 32496 10192
rect 31076 10152 32496 10180
rect 31076 10140 31082 10152
rect 32490 10140 32496 10152
rect 32548 10180 32554 10192
rect 32769 10183 32827 10189
rect 32769 10180 32781 10183
rect 32548 10152 32781 10180
rect 32548 10140 32554 10152
rect 32769 10149 32781 10152
rect 32815 10149 32827 10183
rect 35618 10180 35624 10192
rect 32769 10143 32827 10149
rect 34624 10152 35624 10180
rect 34624 10124 34652 10152
rect 35618 10140 35624 10152
rect 35676 10140 35682 10192
rect 22738 10112 22744 10124
rect 22699 10084 22744 10112
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 22830 10072 22836 10124
rect 22888 10112 22894 10124
rect 22997 10115 23055 10121
rect 22997 10112 23009 10115
rect 22888 10084 23009 10112
rect 22888 10072 22894 10084
rect 22997 10081 23009 10084
rect 23043 10112 23055 10115
rect 24397 10115 24455 10121
rect 24397 10112 24409 10115
rect 23043 10084 24409 10112
rect 23043 10081 23055 10084
rect 22997 10075 23055 10081
rect 24397 10081 24409 10084
rect 24443 10112 24455 10115
rect 25038 10112 25044 10124
rect 24443 10084 25044 10112
rect 24443 10081 24455 10084
rect 24397 10075 24455 10081
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 27338 10072 27344 10124
rect 27396 10112 27402 10124
rect 33505 10115 33563 10121
rect 27396 10084 27568 10112
rect 27396 10072 27402 10084
rect 27430 10044 27436 10056
rect 27391 10016 27436 10044
rect 27430 10004 27436 10016
rect 27488 10004 27494 10056
rect 27540 10053 27568 10084
rect 33505 10081 33517 10115
rect 33551 10112 33563 10115
rect 33962 10112 33968 10124
rect 33551 10084 33968 10112
rect 33551 10081 33563 10084
rect 33505 10075 33563 10081
rect 33962 10072 33968 10084
rect 34020 10072 34026 10124
rect 34606 10072 34612 10124
rect 34664 10072 34670 10124
rect 35437 10115 35495 10121
rect 35437 10081 35449 10115
rect 35483 10112 35495 10115
rect 36262 10112 36268 10124
rect 35483 10084 36268 10112
rect 35483 10081 35495 10084
rect 35437 10075 35495 10081
rect 36262 10072 36268 10084
rect 36320 10072 36326 10124
rect 36538 10112 36544 10124
rect 36499 10084 36544 10112
rect 36538 10072 36544 10084
rect 36596 10072 36602 10124
rect 27525 10047 27583 10053
rect 27525 10013 27537 10047
rect 27571 10044 27583 10047
rect 27614 10044 27620 10056
rect 27571 10016 27620 10044
rect 27571 10013 27583 10016
rect 27525 10007 27583 10013
rect 27614 10004 27620 10016
rect 27672 10004 27678 10056
rect 33045 10047 33103 10053
rect 33045 10013 33057 10047
rect 33091 10044 33103 10047
rect 33410 10044 33416 10056
rect 33091 10016 33416 10044
rect 33091 10013 33103 10016
rect 33045 10007 33103 10013
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 35253 9979 35311 9985
rect 35253 9945 35265 9979
rect 35299 9976 35311 9979
rect 35526 9976 35532 9988
rect 35299 9948 35532 9976
rect 35299 9945 35311 9948
rect 35253 9939 35311 9945
rect 35526 9936 35532 9948
rect 35584 9936 35590 9988
rect 25314 9868 25320 9920
rect 25372 9908 25378 9920
rect 25866 9908 25872 9920
rect 25372 9880 25872 9908
rect 25372 9868 25378 9880
rect 25866 9868 25872 9880
rect 25924 9868 25930 9920
rect 31110 9908 31116 9920
rect 31071 9880 31116 9908
rect 31110 9868 31116 9880
rect 31168 9868 31174 9920
rect 35621 9911 35679 9917
rect 35621 9877 35633 9911
rect 35667 9908 35679 9911
rect 35894 9908 35900 9920
rect 35667 9880 35900 9908
rect 35667 9877 35679 9880
rect 35621 9871 35679 9877
rect 35894 9868 35900 9880
rect 35952 9868 35958 9920
rect 36722 9908 36728 9920
rect 36683 9880 36728 9908
rect 36722 9868 36728 9880
rect 36780 9868 36786 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 22830 9704 22836 9716
rect 22791 9676 22836 9704
rect 22830 9664 22836 9676
rect 22888 9664 22894 9716
rect 26142 9704 26148 9716
rect 26103 9676 26148 9704
rect 26142 9664 26148 9676
rect 26200 9664 26206 9716
rect 26513 9707 26571 9713
rect 26513 9673 26525 9707
rect 26559 9704 26571 9707
rect 27430 9704 27436 9716
rect 26559 9676 27436 9704
rect 26559 9673 26571 9676
rect 26513 9667 26571 9673
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 32490 9704 32496 9716
rect 32451 9676 32496 9704
rect 32490 9664 32496 9676
rect 32548 9664 32554 9716
rect 33962 9704 33968 9716
rect 33923 9676 33968 9704
rect 33962 9664 33968 9676
rect 34020 9664 34026 9716
rect 34146 9704 34152 9716
rect 34072 9676 34152 9704
rect 22465 9639 22523 9645
rect 22465 9605 22477 9639
rect 22511 9636 22523 9639
rect 22738 9636 22744 9648
rect 22511 9608 22744 9636
rect 22511 9605 22523 9608
rect 22465 9599 22523 9605
rect 22738 9596 22744 9608
rect 22796 9596 22802 9648
rect 27614 9596 27620 9648
rect 27672 9636 27678 9648
rect 28353 9639 28411 9645
rect 28353 9636 28365 9639
rect 27672 9608 28365 9636
rect 27672 9596 27678 9608
rect 28353 9605 28365 9608
rect 28399 9605 28411 9639
rect 28353 9599 28411 9605
rect 29641 9639 29699 9645
rect 29641 9605 29653 9639
rect 29687 9636 29699 9639
rect 30837 9639 30895 9645
rect 30837 9636 30849 9639
rect 29687 9608 30849 9636
rect 29687 9605 29699 9608
rect 29641 9599 29699 9605
rect 30837 9605 30849 9608
rect 30883 9636 30895 9639
rect 32125 9639 32183 9645
rect 30883 9608 31524 9636
rect 30883 9605 30895 9608
rect 30837 9599 30895 9605
rect 26881 9571 26939 9577
rect 26881 9537 26893 9571
rect 26927 9568 26939 9571
rect 27893 9571 27951 9577
rect 27893 9568 27905 9571
rect 26927 9540 27905 9568
rect 26927 9537 26939 9540
rect 26881 9531 26939 9537
rect 27893 9537 27905 9540
rect 27939 9568 27951 9571
rect 28258 9568 28264 9580
rect 27939 9540 28264 9568
rect 27939 9537 27951 9540
rect 27893 9531 27951 9537
rect 28258 9528 28264 9540
rect 28316 9528 28322 9580
rect 31496 9577 31524 9608
rect 32125 9605 32137 9639
rect 32171 9636 32183 9639
rect 32582 9636 32588 9648
rect 32171 9608 32588 9636
rect 32171 9605 32183 9608
rect 32125 9599 32183 9605
rect 32582 9596 32588 9608
rect 32640 9596 32646 9648
rect 32861 9639 32919 9645
rect 32861 9605 32873 9639
rect 32907 9636 32919 9639
rect 33042 9636 33048 9648
rect 32907 9608 33048 9636
rect 32907 9605 32919 9608
rect 32861 9599 32919 9605
rect 33042 9596 33048 9608
rect 33100 9596 33106 9648
rect 33870 9596 33876 9648
rect 33928 9636 33934 9648
rect 34072 9636 34100 9676
rect 34146 9664 34152 9676
rect 34204 9664 34210 9716
rect 34606 9664 34612 9716
rect 34664 9704 34670 9716
rect 35250 9704 35256 9716
rect 34664 9676 35256 9704
rect 34664 9664 34670 9676
rect 35250 9664 35256 9676
rect 35308 9664 35314 9716
rect 35894 9704 35900 9716
rect 35636 9676 35900 9704
rect 33928 9608 34100 9636
rect 33928 9596 33934 9608
rect 34514 9596 34520 9648
rect 34572 9636 34578 9648
rect 35161 9639 35219 9645
rect 35161 9636 35173 9639
rect 34572 9608 35173 9636
rect 34572 9596 34578 9608
rect 35161 9605 35173 9608
rect 35207 9605 35219 9639
rect 35161 9599 35219 9605
rect 31481 9571 31539 9577
rect 31481 9537 31493 9571
rect 31527 9537 31539 9571
rect 31481 9531 31539 9537
rect 31573 9571 31631 9577
rect 31573 9537 31585 9571
rect 31619 9537 31631 9571
rect 31573 9531 31631 9537
rect 23750 9500 23756 9512
rect 23711 9472 23756 9500
rect 23750 9460 23756 9472
rect 23808 9460 23814 9512
rect 27614 9460 27620 9512
rect 27672 9500 27678 9512
rect 29457 9503 29515 9509
rect 29457 9500 29469 9503
rect 27672 9472 29469 9500
rect 27672 9460 27678 9472
rect 29457 9469 29469 9472
rect 29503 9500 29515 9503
rect 30009 9503 30067 9509
rect 30009 9500 30021 9503
rect 29503 9472 30021 9500
rect 29503 9469 29515 9472
rect 29457 9463 29515 9469
rect 30009 9469 30021 9472
rect 30055 9469 30067 9503
rect 30009 9463 30067 9469
rect 31110 9460 31116 9512
rect 31168 9500 31174 9512
rect 31389 9503 31447 9509
rect 31389 9500 31401 9503
rect 31168 9472 31401 9500
rect 31168 9460 31174 9472
rect 31389 9469 31401 9472
rect 31435 9469 31447 9503
rect 31389 9463 31447 9469
rect 31588 9444 31616 9531
rect 32950 9528 32956 9580
rect 33008 9568 33014 9580
rect 33413 9571 33471 9577
rect 33413 9568 33425 9571
rect 33008 9540 33425 9568
rect 33008 9528 33014 9540
rect 33413 9537 33425 9540
rect 33459 9537 33471 9571
rect 33413 9531 33471 9537
rect 34606 9528 34612 9580
rect 34664 9568 34670 9580
rect 35636 9568 35664 9676
rect 35894 9664 35900 9676
rect 35952 9664 35958 9716
rect 36538 9704 36544 9716
rect 36499 9676 36544 9704
rect 36538 9664 36544 9676
rect 36596 9664 36602 9716
rect 36262 9636 36268 9648
rect 36223 9608 36268 9636
rect 36262 9596 36268 9608
rect 36320 9596 36326 9648
rect 37182 9596 37188 9648
rect 37240 9636 37246 9648
rect 37277 9639 37335 9645
rect 37277 9636 37289 9639
rect 37240 9608 37289 9636
rect 37240 9596 37246 9608
rect 37277 9605 37289 9608
rect 37323 9605 37335 9639
rect 37277 9599 37335 9605
rect 35713 9571 35771 9577
rect 35713 9568 35725 9571
rect 34664 9540 35725 9568
rect 34664 9528 34670 9540
rect 35713 9537 35725 9540
rect 35759 9537 35771 9571
rect 35713 9531 35771 9537
rect 33226 9500 33232 9512
rect 33139 9472 33232 9500
rect 33226 9460 33232 9472
rect 33284 9500 33290 9512
rect 33962 9500 33968 9512
rect 33284 9472 33968 9500
rect 33284 9460 33290 9472
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 36725 9503 36783 9509
rect 36725 9469 36737 9503
rect 36771 9500 36783 9503
rect 37200 9500 37228 9596
rect 36771 9472 37228 9500
rect 36771 9469 36783 9472
rect 36725 9463 36783 9469
rect 23477 9435 23535 9441
rect 23477 9401 23489 9435
rect 23523 9432 23535 9435
rect 24020 9435 24078 9441
rect 24020 9432 24032 9435
rect 23523 9404 24032 9432
rect 23523 9401 23535 9404
rect 23477 9395 23535 9401
rect 24020 9401 24032 9404
rect 24066 9432 24078 9435
rect 24578 9432 24584 9444
rect 24066 9404 24584 9432
rect 24066 9401 24078 9404
rect 24020 9395 24078 9401
rect 24578 9392 24584 9404
rect 24636 9392 24642 9444
rect 26694 9392 26700 9444
rect 26752 9432 26758 9444
rect 27249 9435 27307 9441
rect 27249 9432 27261 9435
rect 26752 9404 27261 9432
rect 26752 9392 26758 9404
rect 27249 9401 27261 9404
rect 27295 9432 27307 9435
rect 27801 9435 27859 9441
rect 27801 9432 27813 9435
rect 27295 9404 27813 9432
rect 27295 9401 27307 9404
rect 27249 9395 27307 9401
rect 27801 9401 27813 9404
rect 27847 9401 27859 9435
rect 27801 9395 27859 9401
rect 30561 9435 30619 9441
rect 30561 9401 30573 9435
rect 30607 9432 30619 9435
rect 31570 9432 31576 9444
rect 30607 9404 31576 9432
rect 30607 9401 30619 9404
rect 30561 9395 30619 9401
rect 31570 9392 31576 9404
rect 31628 9392 31634 9444
rect 35250 9392 35256 9444
rect 35308 9432 35314 9444
rect 35621 9435 35679 9441
rect 35621 9432 35633 9435
rect 35308 9404 35633 9432
rect 35308 9392 35314 9404
rect 35621 9401 35633 9404
rect 35667 9401 35679 9435
rect 35621 9395 35679 9401
rect 24486 9324 24492 9376
rect 24544 9364 24550 9376
rect 25133 9367 25191 9373
rect 25133 9364 25145 9367
rect 24544 9336 25145 9364
rect 24544 9324 24550 9336
rect 25133 9333 25145 9336
rect 25179 9333 25191 9367
rect 27338 9364 27344 9376
rect 27299 9336 27344 9364
rect 25133 9327 25191 9333
rect 27338 9324 27344 9336
rect 27396 9324 27402 9376
rect 27430 9324 27436 9376
rect 27488 9364 27494 9376
rect 27709 9367 27767 9373
rect 27709 9364 27721 9367
rect 27488 9336 27721 9364
rect 27488 9324 27494 9336
rect 27709 9333 27721 9336
rect 27755 9333 27767 9367
rect 27709 9327 27767 9333
rect 31021 9367 31079 9373
rect 31021 9333 31033 9367
rect 31067 9364 31079 9367
rect 31202 9364 31208 9376
rect 31067 9336 31208 9364
rect 31067 9333 31079 9336
rect 31021 9327 31079 9333
rect 31202 9324 31208 9336
rect 31260 9324 31266 9376
rect 32950 9324 32956 9376
rect 33008 9364 33014 9376
rect 33321 9367 33379 9373
rect 33321 9364 33333 9367
rect 33008 9336 33333 9364
rect 33008 9324 33014 9336
rect 33321 9333 33333 9336
rect 33367 9333 33379 9367
rect 34606 9364 34612 9376
rect 34567 9336 34612 9364
rect 33321 9327 33379 9333
rect 34606 9324 34612 9336
rect 34664 9324 34670 9376
rect 35526 9364 35532 9376
rect 35487 9336 35532 9364
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 36906 9364 36912 9376
rect 36867 9336 36912 9364
rect 36906 9324 36912 9336
rect 36964 9324 36970 9376
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 24121 9163 24179 9169
rect 24121 9129 24133 9163
rect 24167 9160 24179 9163
rect 24670 9160 24676 9172
rect 24167 9132 24676 9160
rect 24167 9129 24179 9132
rect 24121 9123 24179 9129
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 27430 9160 27436 9172
rect 27391 9132 27436 9160
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 31021 9163 31079 9169
rect 31021 9129 31033 9163
rect 31067 9160 31079 9163
rect 31110 9160 31116 9172
rect 31067 9132 31116 9160
rect 31067 9129 31079 9132
rect 31021 9123 31079 9129
rect 31110 9120 31116 9132
rect 31168 9120 31174 9172
rect 31202 9120 31208 9172
rect 31260 9160 31266 9172
rect 33226 9160 33232 9172
rect 31260 9132 32996 9160
rect 33187 9132 33232 9160
rect 31260 9120 31266 9132
rect 32968 9104 32996 9132
rect 33226 9120 33232 9132
rect 33284 9120 33290 9172
rect 34330 9160 34336 9172
rect 34291 9132 34336 9160
rect 34330 9120 34336 9132
rect 34388 9120 34394 9172
rect 36817 9163 36875 9169
rect 36817 9129 36829 9163
rect 36863 9160 36875 9163
rect 37090 9160 37096 9172
rect 36863 9132 37096 9160
rect 36863 9129 36875 9132
rect 36817 9123 36875 9129
rect 37090 9120 37096 9132
rect 37148 9120 37154 9172
rect 24486 9092 24492 9104
rect 24447 9064 24492 9092
rect 24486 9052 24492 9064
rect 24544 9052 24550 9104
rect 24578 9052 24584 9104
rect 24636 9092 24642 9104
rect 31941 9095 31999 9101
rect 24636 9064 24681 9092
rect 24636 9052 24642 9064
rect 31941 9061 31953 9095
rect 31987 9092 31999 9095
rect 32674 9092 32680 9104
rect 31987 9064 32680 9092
rect 31987 9061 31999 9064
rect 31941 9055 31999 9061
rect 32674 9052 32680 9064
rect 32732 9052 32738 9104
rect 32950 9092 32956 9104
rect 32911 9064 32956 9092
rect 32950 9052 32956 9064
rect 33008 9052 33014 9104
rect 34885 9095 34943 9101
rect 34885 9061 34897 9095
rect 34931 9092 34943 9095
rect 35986 9092 35992 9104
rect 34931 9064 35992 9092
rect 34931 9061 34943 9064
rect 34885 9055 34943 9061
rect 23750 8984 23756 9036
rect 23808 9024 23814 9036
rect 23845 9027 23903 9033
rect 23845 9024 23857 9027
rect 23808 8996 23857 9024
rect 23808 8984 23814 8996
rect 23845 8993 23857 8996
rect 23891 9024 23903 9027
rect 25314 9024 25320 9036
rect 23891 8996 25320 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 27154 8984 27160 9036
rect 27212 9024 27218 9036
rect 28077 9027 28135 9033
rect 28077 9024 28089 9027
rect 27212 8996 28089 9024
rect 27212 8984 27218 8996
rect 28077 8993 28089 8996
rect 28123 9024 28135 9027
rect 28810 9024 28816 9036
rect 28123 8996 28816 9024
rect 28123 8993 28135 8996
rect 28077 8987 28135 8993
rect 28810 8984 28816 8996
rect 28868 8984 28874 9036
rect 29181 9027 29239 9033
rect 29181 8993 29193 9027
rect 29227 9024 29239 9027
rect 29638 9024 29644 9036
rect 29227 8996 29644 9024
rect 29227 8993 29239 8996
rect 29181 8987 29239 8993
rect 29638 8984 29644 8996
rect 29696 8984 29702 9036
rect 30837 9027 30895 9033
rect 30837 8993 30849 9027
rect 30883 8993 30895 9027
rect 30837 8987 30895 8993
rect 24210 8916 24216 8968
rect 24268 8956 24274 8968
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 24268 8928 24685 8956
rect 24268 8916 24274 8928
rect 24673 8925 24685 8928
rect 24719 8925 24731 8959
rect 28166 8956 28172 8968
rect 28127 8928 28172 8956
rect 24673 8919 24731 8925
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 28258 8916 28264 8968
rect 28316 8956 28322 8968
rect 28316 8928 28361 8956
rect 28316 8916 28322 8928
rect 28994 8916 29000 8968
rect 29052 8956 29058 8968
rect 29730 8956 29736 8968
rect 29052 8928 29736 8956
rect 29052 8916 29058 8928
rect 29730 8916 29736 8928
rect 29788 8916 29794 8968
rect 29914 8956 29920 8968
rect 29875 8928 29920 8956
rect 29914 8916 29920 8928
rect 29972 8916 29978 8968
rect 30852 8900 30880 8987
rect 32030 8984 32036 9036
rect 32088 9024 32094 9036
rect 32125 9027 32183 9033
rect 32125 9024 32137 9027
rect 32088 8996 32137 9024
rect 32088 8984 32094 8996
rect 32125 8993 32137 8996
rect 32171 8993 32183 9027
rect 32125 8987 32183 8993
rect 33318 8984 33324 9036
rect 33376 9024 33382 9036
rect 35452 9033 35480 9064
rect 35986 9052 35992 9064
rect 36044 9052 36050 9104
rect 33597 9027 33655 9033
rect 33597 9024 33609 9027
rect 33376 8996 33609 9024
rect 33376 8984 33382 8996
rect 33597 8993 33609 8996
rect 33643 8993 33655 9027
rect 33597 8987 33655 8993
rect 35437 9027 35495 9033
rect 35437 8993 35449 9027
rect 35483 8993 35495 9027
rect 35437 8987 35495 8993
rect 35526 8984 35532 9036
rect 35584 9024 35590 9036
rect 35704 9027 35762 9033
rect 35704 9024 35716 9027
rect 35584 8996 35716 9024
rect 35584 8984 35590 8996
rect 35704 8993 35716 8996
rect 35750 9024 35762 9027
rect 36814 9024 36820 9036
rect 35750 8996 36820 9024
rect 35750 8993 35762 8996
rect 35704 8987 35762 8993
rect 36814 8984 36820 8996
rect 36872 8984 36878 9036
rect 33686 8956 33692 8968
rect 33647 8928 33692 8956
rect 33686 8916 33692 8928
rect 33744 8916 33750 8968
rect 33873 8959 33931 8965
rect 33873 8925 33885 8959
rect 33919 8956 33931 8959
rect 34330 8956 34336 8968
rect 33919 8928 34336 8956
rect 33919 8925 33931 8928
rect 33873 8919 33931 8925
rect 34330 8916 34336 8928
rect 34388 8916 34394 8968
rect 27065 8891 27123 8897
rect 27065 8857 27077 8891
rect 27111 8888 27123 8891
rect 29273 8891 29331 8897
rect 27111 8860 28304 8888
rect 27111 8857 27123 8860
rect 27065 8851 27123 8857
rect 28276 8832 28304 8860
rect 29273 8857 29285 8891
rect 29319 8888 29331 8891
rect 30834 8888 30840 8900
rect 29319 8860 30840 8888
rect 29319 8857 29331 8860
rect 29273 8851 29331 8857
rect 30834 8848 30840 8860
rect 30892 8848 30898 8900
rect 27706 8820 27712 8832
rect 27667 8792 27712 8820
rect 27706 8780 27712 8792
rect 27764 8780 27770 8832
rect 28258 8780 28264 8832
rect 28316 8820 28322 8832
rect 28813 8823 28871 8829
rect 28813 8820 28825 8823
rect 28316 8792 28825 8820
rect 28316 8780 28322 8792
rect 28813 8789 28825 8792
rect 28859 8820 28871 8823
rect 29914 8820 29920 8832
rect 28859 8792 29920 8820
rect 28859 8789 28871 8792
rect 28813 8783 28871 8789
rect 29914 8780 29920 8792
rect 29972 8780 29978 8832
rect 30282 8820 30288 8832
rect 30243 8792 30288 8820
rect 30282 8780 30288 8792
rect 30340 8780 30346 8832
rect 32306 8820 32312 8832
rect 32267 8792 32312 8820
rect 32306 8780 32312 8792
rect 32364 8780 32370 8832
rect 35250 8820 35256 8832
rect 35211 8792 35256 8820
rect 35250 8780 35256 8792
rect 35308 8780 35314 8832
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 24486 8616 24492 8628
rect 24447 8588 24492 8616
rect 24486 8576 24492 8588
rect 24544 8576 24550 8628
rect 26694 8616 26700 8628
rect 26655 8588 26700 8616
rect 26694 8576 26700 8588
rect 26752 8576 26758 8628
rect 27154 8616 27160 8628
rect 27115 8588 27160 8616
rect 27154 8576 27160 8588
rect 27212 8576 27218 8628
rect 27525 8619 27583 8625
rect 27525 8585 27537 8619
rect 27571 8616 27583 8619
rect 28166 8616 28172 8628
rect 27571 8588 28172 8616
rect 27571 8585 27583 8588
rect 27525 8579 27583 8585
rect 28166 8576 28172 8588
rect 28224 8576 28230 8628
rect 29638 8616 29644 8628
rect 29599 8588 29644 8616
rect 29638 8576 29644 8588
rect 29696 8576 29702 8628
rect 29730 8576 29736 8628
rect 29788 8616 29794 8628
rect 30653 8619 30711 8625
rect 30653 8616 30665 8619
rect 29788 8588 30665 8616
rect 29788 8576 29794 8588
rect 30653 8585 30665 8588
rect 30699 8585 30711 8619
rect 30653 8579 30711 8585
rect 32306 8576 32312 8628
rect 32364 8616 32370 8628
rect 33229 8619 33287 8625
rect 33229 8616 33241 8619
rect 32364 8588 33241 8616
rect 32364 8576 32370 8588
rect 33229 8585 33241 8588
rect 33275 8616 33287 8619
rect 33686 8616 33692 8628
rect 33275 8588 33692 8616
rect 33275 8585 33287 8588
rect 33229 8579 33287 8585
rect 33686 8576 33692 8588
rect 33744 8576 33750 8628
rect 34701 8619 34759 8625
rect 34701 8585 34713 8619
rect 34747 8616 34759 8619
rect 35434 8616 35440 8628
rect 34747 8588 35440 8616
rect 34747 8585 34759 8588
rect 34701 8579 34759 8585
rect 35434 8576 35440 8588
rect 35492 8576 35498 8628
rect 36814 8616 36820 8628
rect 36775 8588 36820 8616
rect 36814 8576 36820 8588
rect 36872 8576 36878 8628
rect 24394 8508 24400 8560
rect 24452 8548 24458 8560
rect 25133 8551 25191 8557
rect 25133 8548 25145 8551
rect 24452 8520 25145 8548
rect 24452 8508 24458 8520
rect 25133 8517 25145 8520
rect 25179 8517 25191 8551
rect 27614 8548 27620 8560
rect 27575 8520 27620 8548
rect 25133 8511 25191 8517
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8480 24271 8483
rect 24578 8480 24584 8492
rect 24259 8452 24584 8480
rect 24259 8449 24271 8452
rect 24213 8443 24271 8449
rect 24578 8440 24584 8452
rect 24636 8440 24642 8492
rect 25148 8480 25176 8511
rect 27614 8508 27620 8520
rect 27672 8508 27678 8560
rect 28629 8551 28687 8557
rect 28629 8548 28641 8551
rect 28092 8520 28641 8548
rect 25148 8452 25452 8480
rect 25314 8412 25320 8424
rect 25275 8384 25320 8412
rect 25314 8372 25320 8384
rect 25372 8372 25378 8424
rect 25424 8412 25452 8452
rect 27338 8440 27344 8492
rect 27396 8480 27402 8492
rect 28092 8489 28120 8520
rect 28629 8517 28641 8520
rect 28675 8517 28687 8551
rect 33778 8548 33784 8560
rect 28629 8511 28687 8517
rect 31864 8520 33784 8548
rect 31864 8492 31892 8520
rect 28077 8483 28135 8489
rect 28077 8480 28089 8483
rect 27396 8452 28089 8480
rect 27396 8440 27402 8452
rect 28077 8449 28089 8452
rect 28123 8449 28135 8483
rect 28258 8480 28264 8492
rect 28219 8452 28264 8480
rect 28077 8443 28135 8449
rect 28258 8440 28264 8452
rect 28316 8440 28322 8492
rect 28350 8440 28356 8492
rect 28408 8480 28414 8492
rect 30193 8483 30251 8489
rect 30193 8480 30205 8483
rect 28408 8452 30205 8480
rect 28408 8440 28414 8452
rect 30193 8449 30205 8452
rect 30239 8480 30251 8483
rect 30282 8480 30288 8492
rect 30239 8452 30288 8480
rect 30239 8449 30251 8452
rect 30193 8443 30251 8449
rect 30282 8440 30288 8452
rect 30340 8480 30346 8492
rect 31846 8480 31852 8492
rect 30340 8452 31852 8480
rect 30340 8440 30346 8452
rect 31846 8440 31852 8452
rect 31904 8440 31910 8492
rect 32033 8483 32091 8489
rect 32033 8449 32045 8483
rect 32079 8480 32091 8483
rect 32582 8480 32588 8492
rect 32079 8452 32588 8480
rect 32079 8449 32091 8452
rect 32033 8443 32091 8449
rect 32582 8440 32588 8452
rect 32640 8440 32646 8492
rect 32692 8489 32720 8520
rect 33778 8508 33784 8520
rect 33836 8548 33842 8560
rect 34606 8548 34612 8560
rect 33836 8520 34612 8548
rect 33836 8508 33842 8520
rect 34606 8508 34612 8520
rect 34664 8508 34670 8560
rect 32677 8483 32735 8489
rect 32677 8449 32689 8483
rect 32723 8449 32735 8483
rect 32677 8443 32735 8449
rect 25573 8415 25631 8421
rect 25573 8412 25585 8415
rect 25424 8384 25585 8412
rect 25573 8381 25585 8384
rect 25619 8381 25631 8415
rect 25573 8375 25631 8381
rect 27706 8372 27712 8424
rect 27764 8412 27770 8424
rect 27985 8415 28043 8421
rect 27985 8412 27997 8415
rect 27764 8384 27997 8412
rect 27764 8372 27770 8384
rect 27985 8381 27997 8384
rect 28031 8381 28043 8415
rect 27985 8375 28043 8381
rect 29089 8415 29147 8421
rect 29089 8381 29101 8415
rect 29135 8412 29147 8415
rect 30009 8415 30067 8421
rect 30009 8412 30021 8415
rect 29135 8384 30021 8412
rect 29135 8381 29147 8384
rect 29089 8375 29147 8381
rect 30009 8381 30021 8384
rect 30055 8412 30067 8415
rect 31665 8415 31723 8421
rect 30055 8384 30420 8412
rect 30055 8381 30067 8384
rect 30009 8375 30067 8381
rect 29549 8347 29607 8353
rect 29549 8313 29561 8347
rect 29595 8344 29607 8347
rect 30101 8347 30159 8353
rect 30101 8344 30113 8347
rect 29595 8316 30113 8344
rect 29595 8313 29607 8316
rect 29549 8307 29607 8313
rect 30101 8313 30113 8316
rect 30147 8344 30159 8347
rect 30282 8344 30288 8356
rect 30147 8316 30288 8344
rect 30147 8313 30159 8316
rect 30101 8307 30159 8313
rect 30282 8304 30288 8316
rect 30340 8304 30346 8356
rect 30392 8288 30420 8384
rect 31665 8381 31677 8415
rect 31711 8412 31723 8415
rect 32493 8415 32551 8421
rect 32493 8412 32505 8415
rect 31711 8384 32505 8412
rect 31711 8381 31723 8384
rect 31665 8375 31723 8381
rect 32493 8381 32505 8384
rect 32539 8412 32551 8415
rect 32766 8412 32772 8424
rect 32539 8384 32772 8412
rect 32539 8381 32551 8384
rect 32493 8375 32551 8381
rect 32766 8372 32772 8384
rect 32824 8372 32830 8424
rect 33686 8412 33692 8424
rect 33599 8384 33692 8412
rect 33686 8372 33692 8384
rect 33744 8412 33750 8424
rect 34241 8415 34299 8421
rect 34241 8412 34253 8415
rect 33744 8384 34253 8412
rect 33744 8372 33750 8384
rect 34241 8381 34253 8384
rect 34287 8381 34299 8415
rect 35434 8412 35440 8424
rect 35347 8384 35440 8412
rect 34241 8375 34299 8381
rect 35434 8372 35440 8384
rect 35492 8412 35498 8424
rect 35986 8412 35992 8424
rect 35492 8384 35992 8412
rect 35492 8372 35498 8384
rect 35986 8372 35992 8384
rect 36044 8412 36050 8424
rect 36044 8384 37136 8412
rect 36044 8372 36050 8384
rect 31297 8347 31355 8353
rect 31297 8313 31309 8347
rect 31343 8344 31355 8347
rect 32030 8344 32036 8356
rect 31343 8316 32036 8344
rect 31343 8313 31355 8316
rect 31297 8307 31355 8313
rect 32030 8304 32036 8316
rect 32088 8304 32094 8356
rect 35250 8304 35256 8356
rect 35308 8344 35314 8356
rect 35345 8347 35403 8353
rect 35345 8344 35357 8347
rect 35308 8316 35357 8344
rect 35308 8304 35314 8316
rect 35345 8313 35357 8316
rect 35391 8344 35403 8347
rect 35704 8347 35762 8353
rect 35704 8344 35716 8347
rect 35391 8316 35716 8344
rect 35391 8313 35403 8316
rect 35345 8307 35403 8313
rect 35704 8313 35716 8316
rect 35750 8344 35762 8347
rect 35750 8316 35940 8344
rect 35750 8313 35762 8316
rect 35704 8307 35762 8313
rect 30374 8236 30380 8288
rect 30432 8236 30438 8288
rect 32122 8276 32128 8288
rect 32083 8248 32128 8276
rect 32122 8236 32128 8248
rect 32180 8236 32186 8288
rect 33318 8236 33324 8288
rect 33376 8276 33382 8288
rect 33873 8279 33931 8285
rect 33873 8276 33885 8279
rect 33376 8248 33885 8276
rect 33376 8236 33382 8248
rect 33873 8245 33885 8248
rect 33919 8245 33931 8279
rect 35912 8276 35940 8316
rect 37108 8288 37136 8384
rect 36630 8276 36636 8288
rect 35912 8248 36636 8276
rect 33873 8239 33931 8245
rect 36630 8236 36636 8248
rect 36688 8236 36694 8288
rect 37090 8276 37096 8288
rect 37051 8248 37096 8276
rect 37090 8236 37096 8248
rect 37148 8236 37154 8288
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 24210 8072 24216 8084
rect 24171 8044 24216 8072
rect 24210 8032 24216 8044
rect 24268 8032 24274 8084
rect 27706 8032 27712 8084
rect 27764 8072 27770 8084
rect 28169 8075 28227 8081
rect 28169 8072 28181 8075
rect 27764 8044 28181 8072
rect 27764 8032 27770 8044
rect 28169 8041 28181 8044
rect 28215 8041 28227 8075
rect 28169 8035 28227 8041
rect 28350 8032 28356 8084
rect 28408 8072 28414 8084
rect 28537 8075 28595 8081
rect 28537 8072 28549 8075
rect 28408 8044 28549 8072
rect 28408 8032 28414 8044
rect 28537 8041 28549 8044
rect 28583 8041 28595 8075
rect 30834 8072 30840 8084
rect 30795 8044 30840 8072
rect 28537 8035 28595 8041
rect 30834 8032 30840 8044
rect 30892 8032 30898 8084
rect 31846 8072 31852 8084
rect 31807 8044 31852 8072
rect 31846 8032 31852 8044
rect 31904 8032 31910 8084
rect 32122 8032 32128 8084
rect 32180 8072 32186 8084
rect 32585 8075 32643 8081
rect 32585 8072 32597 8075
rect 32180 8044 32597 8072
rect 32180 8032 32186 8044
rect 32585 8041 32597 8044
rect 32631 8041 32643 8075
rect 33318 8072 33324 8084
rect 33279 8044 33324 8072
rect 32585 8035 32643 8041
rect 33318 8032 33324 8044
rect 33376 8032 33382 8084
rect 33686 8072 33692 8084
rect 33647 8044 33692 8072
rect 33686 8032 33692 8044
rect 33744 8032 33750 8084
rect 34057 8075 34115 8081
rect 34057 8041 34069 8075
rect 34103 8072 34115 8075
rect 34422 8072 34428 8084
rect 34103 8044 34428 8072
rect 34103 8041 34115 8044
rect 34057 8035 34115 8041
rect 34422 8032 34428 8044
rect 34480 8032 34486 8084
rect 36630 8072 36636 8084
rect 36591 8044 36636 8072
rect 36630 8032 36636 8044
rect 36688 8032 36694 8084
rect 26694 7964 26700 8016
rect 26752 8013 26758 8016
rect 26752 8007 26816 8013
rect 26752 7973 26770 8007
rect 26804 7973 26816 8007
rect 35434 8004 35440 8016
rect 26752 7967 26816 7973
rect 35268 7976 35440 8004
rect 26752 7964 26758 7967
rect 28994 7945 29000 7948
rect 28988 7936 29000 7945
rect 28955 7908 29000 7936
rect 28988 7899 29000 7908
rect 28994 7896 29000 7899
rect 29052 7896 29058 7948
rect 32490 7936 32496 7948
rect 32451 7908 32496 7936
rect 32490 7896 32496 7908
rect 32548 7896 32554 7948
rect 35268 7945 35296 7976
rect 35434 7964 35440 7976
rect 35492 7964 35498 8016
rect 34977 7939 35035 7945
rect 34977 7905 34989 7939
rect 35023 7936 35035 7939
rect 35253 7939 35311 7945
rect 35253 7936 35265 7939
rect 35023 7908 35265 7936
rect 35023 7905 35035 7908
rect 34977 7899 35035 7905
rect 35253 7905 35265 7908
rect 35299 7905 35311 7939
rect 35253 7899 35311 7905
rect 35520 7939 35578 7945
rect 35520 7905 35532 7939
rect 35566 7936 35578 7939
rect 36538 7936 36544 7948
rect 35566 7908 36544 7936
rect 35566 7905 35578 7908
rect 35520 7899 35578 7905
rect 36538 7896 36544 7908
rect 36596 7896 36602 7948
rect 25314 7828 25320 7880
rect 25372 7868 25378 7880
rect 25409 7871 25467 7877
rect 25409 7868 25421 7871
rect 25372 7840 25421 7868
rect 25372 7828 25378 7840
rect 25409 7837 25421 7840
rect 25455 7868 25467 7871
rect 26234 7868 26240 7880
rect 25455 7840 26240 7868
rect 25455 7837 25467 7840
rect 25409 7831 25467 7837
rect 26234 7828 26240 7840
rect 26292 7868 26298 7880
rect 26513 7871 26571 7877
rect 26513 7868 26525 7871
rect 26292 7840 26525 7868
rect 26292 7828 26298 7840
rect 26513 7837 26525 7840
rect 26559 7837 26571 7871
rect 28718 7868 28724 7880
rect 28679 7840 28724 7868
rect 26513 7831 26571 7837
rect 28718 7828 28724 7840
rect 28776 7828 28782 7880
rect 31938 7828 31944 7880
rect 31996 7868 32002 7880
rect 32769 7871 32827 7877
rect 32769 7868 32781 7871
rect 31996 7840 32781 7868
rect 31996 7828 32002 7840
rect 32769 7837 32781 7840
rect 32815 7837 32827 7871
rect 34146 7868 34152 7880
rect 34107 7840 34152 7868
rect 32769 7831 32827 7837
rect 32030 7760 32036 7812
rect 32088 7800 32094 7812
rect 32125 7803 32183 7809
rect 32125 7800 32137 7803
rect 32088 7772 32137 7800
rect 32088 7760 32094 7772
rect 32125 7769 32137 7772
rect 32171 7769 32183 7803
rect 32784 7800 32812 7831
rect 34146 7828 34152 7840
rect 34204 7828 34210 7880
rect 34330 7868 34336 7880
rect 34291 7840 34336 7868
rect 34330 7828 34336 7840
rect 34388 7828 34394 7880
rect 34348 7800 34376 7828
rect 32784 7772 34376 7800
rect 32125 7763 32183 7769
rect 27430 7692 27436 7744
rect 27488 7732 27494 7744
rect 27893 7735 27951 7741
rect 27893 7732 27905 7735
rect 27488 7704 27905 7732
rect 27488 7692 27494 7704
rect 27893 7701 27905 7704
rect 27939 7701 27951 7735
rect 30098 7732 30104 7744
rect 30059 7704 30104 7732
rect 27893 7695 27951 7701
rect 30098 7692 30104 7704
rect 30156 7692 30162 7744
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 26234 7528 26240 7540
rect 26195 7500 26240 7528
rect 26234 7488 26240 7500
rect 26292 7488 26298 7540
rect 26605 7531 26663 7537
rect 26605 7497 26617 7531
rect 26651 7528 26663 7531
rect 26694 7528 26700 7540
rect 26651 7500 26700 7528
rect 26651 7497 26663 7500
rect 26605 7491 26663 7497
rect 26694 7488 26700 7500
rect 26752 7488 26758 7540
rect 28166 7488 28172 7540
rect 28224 7528 28230 7540
rect 28261 7531 28319 7537
rect 28261 7528 28273 7531
rect 28224 7500 28273 7528
rect 28224 7488 28230 7500
rect 28261 7497 28273 7500
rect 28307 7497 28319 7531
rect 28261 7491 28319 7497
rect 28721 7531 28779 7537
rect 28721 7497 28733 7531
rect 28767 7528 28779 7531
rect 28994 7528 29000 7540
rect 28767 7500 29000 7528
rect 28767 7497 28779 7500
rect 28721 7491 28779 7497
rect 28994 7488 29000 7500
rect 29052 7528 29058 7540
rect 30653 7531 30711 7537
rect 30653 7528 30665 7531
rect 29052 7500 30665 7528
rect 29052 7488 29058 7500
rect 30653 7497 30665 7500
rect 30699 7497 30711 7531
rect 30653 7491 30711 7497
rect 32490 7488 32496 7540
rect 32548 7528 32554 7540
rect 33137 7531 33195 7537
rect 33137 7528 33149 7531
rect 32548 7500 33149 7528
rect 32548 7488 32554 7500
rect 33137 7497 33149 7500
rect 33183 7528 33195 7531
rect 33226 7528 33232 7540
rect 33183 7500 33232 7528
rect 33183 7497 33195 7500
rect 33137 7491 33195 7497
rect 33226 7488 33232 7500
rect 33284 7488 33290 7540
rect 34149 7531 34207 7537
rect 34149 7497 34161 7531
rect 34195 7528 34207 7531
rect 34422 7528 34428 7540
rect 34195 7500 34428 7528
rect 34195 7497 34207 7500
rect 34149 7491 34207 7497
rect 34422 7488 34428 7500
rect 34480 7488 34486 7540
rect 37001 7531 37059 7537
rect 37001 7497 37013 7531
rect 37047 7528 37059 7531
rect 37090 7528 37096 7540
rect 37047 7500 37096 7528
rect 37047 7497 37059 7500
rect 37001 7491 37059 7497
rect 37090 7488 37096 7500
rect 37148 7488 37154 7540
rect 30374 7420 30380 7472
rect 30432 7460 30438 7472
rect 30926 7460 30932 7472
rect 30432 7432 30932 7460
rect 30432 7420 30438 7432
rect 30926 7420 30932 7432
rect 30984 7460 30990 7472
rect 31297 7463 31355 7469
rect 31297 7460 31309 7463
rect 30984 7432 31309 7460
rect 30984 7420 30990 7432
rect 31297 7429 31309 7432
rect 31343 7429 31355 7463
rect 31297 7423 31355 7429
rect 28810 7352 28816 7404
rect 28868 7392 28874 7404
rect 28997 7395 29055 7401
rect 28997 7392 29009 7395
rect 28868 7364 29009 7392
rect 28868 7352 28874 7364
rect 28997 7361 29009 7364
rect 29043 7392 29055 7395
rect 29043 7364 29408 7392
rect 29043 7361 29055 7364
rect 28997 7355 29055 7361
rect 26881 7327 26939 7333
rect 26881 7293 26893 7327
rect 26927 7293 26939 7327
rect 26881 7287 26939 7293
rect 27148 7327 27206 7333
rect 27148 7293 27160 7327
rect 27194 7324 27206 7327
rect 27430 7324 27436 7336
rect 27194 7296 27436 7324
rect 27194 7293 27206 7296
rect 27148 7287 27206 7293
rect 26896 7256 26924 7287
rect 27430 7284 27436 7296
rect 27488 7284 27494 7336
rect 28718 7284 28724 7336
rect 28776 7324 28782 7336
rect 29270 7324 29276 7336
rect 28776 7296 29276 7324
rect 28776 7284 28782 7296
rect 29270 7284 29276 7296
rect 29328 7284 29334 7336
rect 29380 7324 29408 7364
rect 29529 7327 29587 7333
rect 29529 7324 29541 7327
rect 29380 7296 29541 7324
rect 29529 7293 29541 7296
rect 29575 7293 29587 7327
rect 29529 7287 29587 7293
rect 27246 7256 27252 7268
rect 26896 7228 27252 7256
rect 27246 7216 27252 7228
rect 27304 7216 27310 7268
rect 31312 7256 31340 7423
rect 32582 7420 32588 7472
rect 32640 7460 32646 7472
rect 32861 7463 32919 7469
rect 32861 7460 32873 7463
rect 32640 7432 32873 7460
rect 32640 7420 32646 7432
rect 32861 7429 32873 7432
rect 32907 7429 32919 7463
rect 32861 7423 32919 7429
rect 31478 7324 31484 7336
rect 31439 7296 31484 7324
rect 31478 7284 31484 7296
rect 31536 7284 31542 7336
rect 34882 7324 34888 7336
rect 34795 7296 34888 7324
rect 34882 7284 34888 7296
rect 34940 7324 34946 7336
rect 35434 7324 35440 7336
rect 34940 7296 35440 7324
rect 34940 7284 34946 7296
rect 35434 7284 35440 7296
rect 35492 7284 35498 7336
rect 31726 7259 31784 7265
rect 31726 7256 31738 7259
rect 31312 7228 31738 7256
rect 31726 7225 31738 7228
rect 31772 7225 31784 7259
rect 35130 7259 35188 7265
rect 35130 7256 35142 7259
rect 31726 7219 31784 7225
rect 34624 7228 35142 7256
rect 34624 7200 34652 7228
rect 35130 7225 35142 7228
rect 35176 7225 35188 7259
rect 35130 7219 35188 7225
rect 33781 7191 33839 7197
rect 33781 7157 33793 7191
rect 33827 7188 33839 7191
rect 34146 7188 34152 7200
rect 33827 7160 34152 7188
rect 33827 7157 33839 7160
rect 33781 7151 33839 7157
rect 34146 7148 34152 7160
rect 34204 7188 34210 7200
rect 34422 7188 34428 7200
rect 34204 7160 34428 7188
rect 34204 7148 34210 7160
rect 34422 7148 34428 7160
rect 34480 7148 34486 7200
rect 34606 7188 34612 7200
rect 34567 7160 34612 7188
rect 34606 7148 34612 7160
rect 34664 7148 34670 7200
rect 35894 7148 35900 7200
rect 35952 7188 35958 7200
rect 36265 7191 36323 7197
rect 36265 7188 36277 7191
rect 35952 7160 36277 7188
rect 35952 7148 35958 7160
rect 36265 7157 36277 7160
rect 36311 7157 36323 7191
rect 36538 7188 36544 7200
rect 36499 7160 36544 7188
rect 36265 7151 36323 7157
rect 36538 7148 36544 7160
rect 36596 7148 36602 7200
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 26973 6987 27031 6993
rect 26973 6953 26985 6987
rect 27019 6984 27031 6987
rect 27430 6984 27436 6996
rect 27019 6956 27436 6984
rect 27019 6953 27031 6956
rect 26973 6947 27031 6953
rect 27430 6944 27436 6956
rect 27488 6944 27494 6996
rect 31938 6984 31944 6996
rect 31899 6956 31944 6984
rect 31938 6944 31944 6956
rect 31996 6944 32002 6996
rect 32122 6944 32128 6996
rect 32180 6984 32186 6996
rect 32309 6987 32367 6993
rect 32309 6984 32321 6987
rect 32180 6956 32321 6984
rect 32180 6944 32186 6956
rect 32309 6953 32321 6956
rect 32355 6953 32367 6987
rect 32309 6947 32367 6953
rect 34241 6987 34299 6993
rect 34241 6953 34253 6987
rect 34287 6984 34299 6987
rect 34330 6984 34336 6996
rect 34287 6956 34336 6984
rect 34287 6953 34299 6956
rect 34241 6947 34299 6953
rect 34330 6944 34336 6956
rect 34388 6944 34394 6996
rect 34606 6944 34612 6996
rect 34664 6984 34670 6996
rect 36081 6987 36139 6993
rect 36081 6984 36093 6987
rect 34664 6956 36093 6984
rect 34664 6944 34670 6956
rect 36081 6953 36093 6956
rect 36127 6953 36139 6987
rect 36081 6947 36139 6953
rect 28166 6916 28172 6928
rect 27540 6888 28172 6916
rect 27338 6808 27344 6860
rect 27396 6848 27402 6860
rect 27540 6857 27568 6888
rect 28166 6876 28172 6888
rect 28224 6876 28230 6928
rect 29086 6876 29092 6928
rect 29144 6916 29150 6928
rect 29724 6919 29782 6925
rect 29724 6916 29736 6919
rect 29144 6888 29736 6916
rect 29144 6876 29150 6888
rect 29724 6885 29736 6888
rect 29770 6916 29782 6919
rect 30098 6916 30104 6928
rect 29770 6888 30104 6916
rect 29770 6885 29782 6888
rect 29724 6879 29782 6885
rect 30098 6876 30104 6888
rect 30156 6876 30162 6928
rect 35066 6916 35072 6928
rect 34716 6888 35072 6916
rect 27516 6851 27574 6857
rect 27516 6848 27528 6851
rect 27396 6820 27528 6848
rect 27396 6808 27402 6820
rect 27516 6817 27528 6820
rect 27562 6817 27574 6851
rect 27516 6811 27574 6817
rect 28997 6851 29055 6857
rect 28997 6817 29009 6851
rect 29043 6848 29055 6851
rect 29270 6848 29276 6860
rect 29043 6820 29276 6848
rect 29043 6817 29055 6820
rect 28997 6811 29055 6817
rect 29270 6808 29276 6820
rect 29328 6848 29334 6860
rect 29365 6851 29423 6857
rect 29365 6848 29377 6851
rect 29328 6820 29377 6848
rect 29328 6808 29334 6820
rect 29365 6817 29377 6820
rect 29411 6848 29423 6851
rect 29457 6851 29515 6857
rect 29457 6848 29469 6851
rect 29411 6820 29469 6848
rect 29411 6817 29423 6820
rect 29365 6811 29423 6817
rect 29457 6817 29469 6820
rect 29503 6848 29515 6851
rect 29546 6848 29552 6860
rect 29503 6820 29552 6848
rect 29503 6817 29515 6820
rect 29457 6811 29515 6817
rect 29546 6808 29552 6820
rect 29604 6808 29610 6860
rect 32766 6857 32772 6860
rect 32760 6848 32772 6857
rect 32727 6820 32772 6848
rect 32760 6811 32772 6820
rect 32766 6808 32772 6811
rect 32824 6808 32830 6860
rect 34716 6857 34744 6888
rect 35066 6876 35072 6888
rect 35124 6876 35130 6928
rect 34701 6851 34759 6857
rect 34701 6817 34713 6851
rect 34747 6817 34759 6851
rect 34957 6851 35015 6857
rect 34957 6848 34969 6851
rect 34701 6811 34759 6817
rect 34808 6820 34969 6848
rect 27246 6780 27252 6792
rect 27207 6752 27252 6780
rect 27246 6740 27252 6752
rect 27304 6740 27310 6792
rect 31478 6740 31484 6792
rect 31536 6780 31542 6792
rect 31573 6783 31631 6789
rect 31573 6780 31585 6783
rect 31536 6752 31585 6780
rect 31536 6740 31542 6752
rect 31573 6749 31585 6752
rect 31619 6780 31631 6783
rect 32490 6780 32496 6792
rect 31619 6752 32496 6780
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 32490 6740 32496 6752
rect 32548 6740 32554 6792
rect 34808 6780 34836 6820
rect 34957 6817 34969 6820
rect 35003 6817 35015 6851
rect 34957 6811 35015 6817
rect 34716 6752 34836 6780
rect 28629 6715 28687 6721
rect 28629 6681 28641 6715
rect 28675 6712 28687 6715
rect 28810 6712 28816 6724
rect 28675 6684 28816 6712
rect 28675 6681 28687 6684
rect 28629 6675 28687 6681
rect 28810 6672 28816 6684
rect 28868 6672 28874 6724
rect 34716 6712 34744 6752
rect 33888 6684 34744 6712
rect 30374 6604 30380 6656
rect 30432 6644 30438 6656
rect 30837 6647 30895 6653
rect 30837 6644 30849 6647
rect 30432 6616 30849 6644
rect 30432 6604 30438 6616
rect 30837 6613 30849 6616
rect 30883 6613 30895 6647
rect 30837 6607 30895 6613
rect 33686 6604 33692 6656
rect 33744 6644 33750 6656
rect 33888 6653 33916 6684
rect 33873 6647 33931 6653
rect 33873 6644 33885 6647
rect 33744 6616 33885 6644
rect 33744 6604 33750 6616
rect 33873 6613 33885 6616
rect 33919 6613 33931 6647
rect 33873 6607 33931 6613
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 27338 6440 27344 6452
rect 27299 6412 27344 6440
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 29086 6440 29092 6452
rect 29047 6412 29092 6440
rect 29086 6400 29092 6412
rect 29144 6400 29150 6452
rect 30926 6440 30932 6452
rect 30887 6412 30932 6440
rect 30926 6400 30932 6412
rect 30984 6400 30990 6452
rect 32766 6400 32772 6452
rect 32824 6440 32830 6452
rect 33137 6443 33195 6449
rect 33137 6440 33149 6443
rect 32824 6412 33149 6440
rect 32824 6400 32830 6412
rect 33137 6409 33149 6412
rect 33183 6409 33195 6443
rect 33137 6403 33195 6409
rect 36265 6443 36323 6449
rect 36265 6409 36277 6443
rect 36311 6440 36323 6443
rect 36538 6440 36544 6452
rect 36311 6412 36544 6440
rect 36311 6409 36323 6412
rect 36265 6403 36323 6409
rect 36538 6400 36544 6412
rect 36596 6400 36602 6452
rect 36633 6443 36691 6449
rect 36633 6409 36645 6443
rect 36679 6440 36691 6443
rect 37090 6440 37096 6452
rect 36679 6412 37096 6440
rect 36679 6409 36691 6412
rect 36633 6403 36691 6409
rect 37090 6400 37096 6412
rect 37148 6400 37154 6452
rect 31665 6307 31723 6313
rect 31665 6273 31677 6307
rect 31711 6304 31723 6307
rect 34333 6307 34391 6313
rect 31711 6276 31892 6304
rect 31711 6273 31723 6276
rect 31665 6267 31723 6273
rect 26973 6239 27031 6245
rect 26973 6205 26985 6239
rect 27019 6236 27031 6239
rect 27246 6236 27252 6248
rect 27019 6208 27252 6236
rect 27019 6205 27031 6208
rect 26973 6199 27031 6205
rect 27246 6196 27252 6208
rect 27304 6236 27310 6248
rect 27709 6239 27767 6245
rect 27709 6236 27721 6239
rect 27304 6208 27721 6236
rect 27304 6196 27310 6208
rect 27709 6205 27721 6208
rect 27755 6236 27767 6239
rect 28721 6239 28779 6245
rect 28721 6236 28733 6239
rect 27755 6208 28733 6236
rect 27755 6205 27767 6208
rect 27709 6199 27767 6205
rect 28721 6205 28733 6208
rect 28767 6236 28779 6239
rect 29546 6236 29552 6248
rect 28767 6208 29552 6236
rect 28767 6205 28779 6208
rect 28721 6199 28779 6205
rect 29546 6196 29552 6208
rect 29604 6196 29610 6248
rect 29822 6245 29828 6248
rect 29816 6236 29828 6245
rect 29735 6208 29828 6236
rect 29816 6199 29828 6208
rect 29880 6236 29886 6248
rect 30374 6236 30380 6248
rect 29880 6208 30380 6236
rect 29822 6196 29828 6199
rect 29880 6196 29886 6208
rect 30374 6196 30380 6208
rect 30432 6196 30438 6248
rect 31754 6236 31760 6248
rect 31715 6208 31760 6236
rect 31754 6196 31760 6208
rect 31812 6196 31818 6248
rect 31864 6236 31892 6276
rect 34333 6273 34345 6307
rect 34379 6304 34391 6307
rect 34379 6276 35020 6304
rect 34379 6273 34391 6276
rect 34333 6267 34391 6273
rect 32024 6239 32082 6245
rect 32024 6236 32036 6239
rect 31864 6208 32036 6236
rect 32024 6205 32036 6208
rect 32070 6236 32082 6239
rect 32582 6236 32588 6248
rect 32070 6208 32588 6236
rect 32070 6205 32082 6208
rect 32024 6199 32082 6205
rect 32582 6196 32588 6208
rect 32640 6196 32646 6248
rect 34790 6196 34796 6248
rect 34848 6236 34854 6248
rect 34885 6239 34943 6245
rect 34885 6236 34897 6239
rect 34848 6208 34897 6236
rect 34848 6196 34854 6208
rect 34885 6205 34897 6208
rect 34931 6205 34943 6239
rect 34992 6236 35020 6276
rect 35152 6239 35210 6245
rect 35152 6236 35164 6239
rect 34992 6208 35164 6236
rect 34885 6199 34943 6205
rect 35152 6205 35164 6208
rect 35198 6236 35210 6239
rect 35434 6236 35440 6248
rect 35198 6208 35440 6236
rect 35198 6205 35210 6208
rect 35152 6199 35210 6205
rect 35434 6196 35440 6208
rect 35492 6236 35498 6248
rect 35894 6236 35900 6248
rect 35492 6208 35900 6236
rect 35492 6196 35498 6208
rect 35894 6196 35900 6208
rect 35952 6196 35958 6248
rect 33686 6060 33692 6112
rect 33744 6100 33750 6112
rect 34609 6103 34667 6109
rect 34609 6100 34621 6103
rect 33744 6072 34621 6100
rect 33744 6060 33750 6072
rect 34609 6069 34621 6072
rect 34655 6069 34667 6103
rect 34609 6063 34667 6069
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 28813 5899 28871 5905
rect 28813 5865 28825 5899
rect 28859 5896 28871 5899
rect 28902 5896 28908 5908
rect 28859 5868 28908 5896
rect 28859 5865 28871 5868
rect 28813 5859 28871 5865
rect 28902 5856 28908 5868
rect 28960 5856 28966 5908
rect 29086 5856 29092 5908
rect 29144 5896 29150 5908
rect 29181 5899 29239 5905
rect 29181 5896 29193 5899
rect 29144 5868 29193 5896
rect 29144 5856 29150 5868
rect 29181 5865 29193 5868
rect 29227 5865 29239 5899
rect 29822 5896 29828 5908
rect 29783 5868 29828 5896
rect 29181 5859 29239 5865
rect 29822 5856 29828 5868
rect 29880 5856 29886 5908
rect 32585 5899 32643 5905
rect 32585 5865 32597 5899
rect 32631 5896 32643 5899
rect 32766 5896 32772 5908
rect 32631 5868 32772 5896
rect 32631 5865 32643 5868
rect 32585 5859 32643 5865
rect 32766 5856 32772 5868
rect 32824 5856 32830 5908
rect 33226 5896 33232 5908
rect 33187 5868 33232 5896
rect 33226 5856 33232 5868
rect 33284 5856 33290 5908
rect 34514 5856 34520 5908
rect 34572 5896 34578 5908
rect 34885 5899 34943 5905
rect 34885 5896 34897 5899
rect 34572 5868 34897 5896
rect 34572 5856 34578 5868
rect 34885 5865 34897 5868
rect 34931 5865 34943 5899
rect 34885 5859 34943 5865
rect 35253 5899 35311 5905
rect 35253 5865 35265 5899
rect 35299 5896 35311 5899
rect 35526 5896 35532 5908
rect 35299 5868 35532 5896
rect 35299 5865 35311 5868
rect 35253 5859 35311 5865
rect 35526 5856 35532 5868
rect 35584 5896 35590 5908
rect 36538 5896 36544 5908
rect 35584 5868 36544 5896
rect 35584 5856 35590 5868
rect 36538 5856 36544 5868
rect 36596 5856 36602 5908
rect 28994 5788 29000 5840
rect 29052 5828 29058 5840
rect 29273 5831 29331 5837
rect 29273 5828 29285 5831
rect 29052 5800 29285 5828
rect 29052 5788 29058 5800
rect 29273 5797 29285 5800
rect 29319 5797 29331 5831
rect 29273 5791 29331 5797
rect 29546 5788 29552 5840
rect 29604 5828 29610 5840
rect 30285 5831 30343 5837
rect 30285 5828 30297 5831
rect 29604 5800 30297 5828
rect 29604 5788 29610 5800
rect 30285 5797 30297 5800
rect 30331 5828 30343 5831
rect 31754 5828 31760 5840
rect 30331 5800 31760 5828
rect 30331 5797 30343 5800
rect 30285 5791 30343 5797
rect 31754 5788 31760 5800
rect 31812 5828 31818 5840
rect 31849 5831 31907 5837
rect 31849 5828 31861 5831
rect 31812 5800 31861 5828
rect 31812 5788 31818 5800
rect 31849 5797 31861 5800
rect 31895 5828 31907 5831
rect 32490 5828 32496 5840
rect 31895 5800 32496 5828
rect 31895 5797 31907 5800
rect 31849 5791 31907 5797
rect 32490 5788 32496 5800
rect 32548 5828 32554 5840
rect 32953 5831 33011 5837
rect 32953 5828 32965 5831
rect 32548 5800 32965 5828
rect 32548 5788 32554 5800
rect 32953 5797 32965 5800
rect 32999 5828 33011 5831
rect 34790 5828 34796 5840
rect 32999 5800 34796 5828
rect 32999 5797 33011 5800
rect 32953 5791 33011 5797
rect 34790 5788 34796 5800
rect 34848 5788 34854 5840
rect 35345 5831 35403 5837
rect 35345 5797 35357 5831
rect 35391 5828 35403 5831
rect 35434 5828 35440 5840
rect 35391 5800 35440 5828
rect 35391 5797 35403 5800
rect 35345 5791 35403 5797
rect 35434 5788 35440 5800
rect 35492 5788 35498 5840
rect 33594 5760 33600 5772
rect 33555 5732 33600 5760
rect 33594 5720 33600 5732
rect 33652 5760 33658 5772
rect 34606 5760 34612 5772
rect 33652 5732 34612 5760
rect 33652 5720 33658 5732
rect 34606 5720 34612 5732
rect 34664 5720 34670 5772
rect 28350 5652 28356 5704
rect 28408 5692 28414 5704
rect 29365 5695 29423 5701
rect 29365 5692 29377 5695
rect 28408 5664 29377 5692
rect 28408 5652 28414 5664
rect 29365 5661 29377 5664
rect 29411 5661 29423 5695
rect 33686 5692 33692 5704
rect 33647 5664 33692 5692
rect 29365 5655 29423 5661
rect 33686 5652 33692 5664
rect 33744 5652 33750 5704
rect 33778 5652 33784 5704
rect 33836 5692 33842 5704
rect 35437 5695 35495 5701
rect 35437 5692 35449 5695
rect 33836 5664 35449 5692
rect 33836 5652 33842 5664
rect 35437 5661 35449 5664
rect 35483 5661 35495 5695
rect 35437 5655 35495 5661
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 28350 5312 28356 5364
rect 28408 5352 28414 5364
rect 28537 5355 28595 5361
rect 28537 5352 28549 5355
rect 28408 5324 28549 5352
rect 28408 5312 28414 5324
rect 28537 5321 28549 5324
rect 28583 5321 28595 5355
rect 28902 5352 28908 5364
rect 28863 5324 28908 5352
rect 28537 5315 28595 5321
rect 28902 5312 28908 5324
rect 28960 5312 28966 5364
rect 29086 5312 29092 5364
rect 29144 5352 29150 5364
rect 29457 5355 29515 5361
rect 29457 5352 29469 5355
rect 29144 5324 29469 5352
rect 29144 5312 29150 5324
rect 29457 5321 29469 5324
rect 29503 5321 29515 5355
rect 29457 5315 29515 5321
rect 33321 5355 33379 5361
rect 33321 5321 33333 5355
rect 33367 5352 33379 5355
rect 33686 5352 33692 5364
rect 33367 5324 33692 5352
rect 33367 5321 33379 5324
rect 33321 5315 33379 5321
rect 33686 5312 33692 5324
rect 33744 5312 33750 5364
rect 33778 5312 33784 5364
rect 33836 5352 33842 5364
rect 33965 5355 34023 5361
rect 33965 5352 33977 5355
rect 33836 5324 33977 5352
rect 33836 5312 33842 5324
rect 33965 5321 33977 5324
rect 34011 5352 34023 5355
rect 34609 5355 34667 5361
rect 34609 5352 34621 5355
rect 34011 5324 34621 5352
rect 34011 5321 34023 5324
rect 33965 5315 34023 5321
rect 34609 5321 34621 5324
rect 34655 5321 34667 5355
rect 35526 5352 35532 5364
rect 35487 5324 35532 5352
rect 34609 5315 34667 5321
rect 35526 5312 35532 5324
rect 35584 5312 35590 5364
rect 33594 5284 33600 5296
rect 33555 5256 33600 5284
rect 33594 5244 33600 5256
rect 33652 5244 33658 5296
rect 35161 5287 35219 5293
rect 35161 5253 35173 5287
rect 35207 5284 35219 5287
rect 35434 5284 35440 5296
rect 35207 5256 35440 5284
rect 35207 5253 35219 5256
rect 35161 5247 35219 5253
rect 35434 5244 35440 5256
rect 35492 5244 35498 5296
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 33870 2632 33876 2644
rect 33831 2604 33876 2632
rect 33870 2592 33876 2604
rect 33928 2592 33934 2644
rect 33321 2499 33379 2505
rect 33321 2465 33333 2499
rect 33367 2496 33379 2499
rect 33888 2496 33916 2592
rect 36630 2496 36636 2508
rect 33367 2468 36636 2496
rect 33367 2465 33379 2468
rect 33321 2459 33379 2465
rect 36630 2456 36636 2468
rect 36688 2456 36694 2508
rect 33502 2360 33508 2372
rect 33463 2332 33508 2360
rect 33502 2320 33508 2332
rect 33560 2320 33566 2372
rect 8389 2295 8447 2301
rect 8389 2261 8401 2295
rect 8435 2292 8447 2295
rect 9950 2292 9956 2304
rect 8435 2264 9956 2292
rect 8435 2261 8447 2264
rect 8389 2255 8447 2261
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 7196 36864 7248 36916
rect 7472 36567 7524 36576
rect 7472 36533 7481 36567
rect 7481 36533 7515 36567
rect 7515 36533 7524 36567
rect 7472 36524 7524 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 22836 36252 22888 36304
rect 6828 36227 6880 36236
rect 6828 36193 6837 36227
rect 6837 36193 6871 36227
rect 6871 36193 6880 36227
rect 6828 36184 6880 36193
rect 15660 36227 15712 36236
rect 15660 36193 15669 36227
rect 15669 36193 15703 36227
rect 15703 36193 15712 36227
rect 15660 36184 15712 36193
rect 24768 36184 24820 36236
rect 15752 36159 15804 36168
rect 15752 36125 15761 36159
rect 15761 36125 15795 36159
rect 15795 36125 15804 36159
rect 15752 36116 15804 36125
rect 15936 36159 15988 36168
rect 15936 36125 15945 36159
rect 15945 36125 15979 36159
rect 15979 36125 15988 36159
rect 15936 36116 15988 36125
rect 22468 36116 22520 36168
rect 22928 36159 22980 36168
rect 22928 36125 22937 36159
rect 22937 36125 22971 36159
rect 22971 36125 22980 36159
rect 22928 36116 22980 36125
rect 7380 35980 7432 36032
rect 14004 36023 14056 36032
rect 14004 35989 14013 36023
rect 14013 35989 14047 36023
rect 14047 35989 14056 36023
rect 14004 35980 14056 35989
rect 15200 35980 15252 36032
rect 21732 35980 21784 36032
rect 22284 36023 22336 36032
rect 22284 35989 22293 36023
rect 22293 35989 22327 36023
rect 22327 35989 22336 36023
rect 22284 35980 22336 35989
rect 24216 35980 24268 36032
rect 24952 36023 25004 36032
rect 24952 35989 24961 36023
rect 24961 35989 24995 36023
rect 24995 35989 25004 36023
rect 24952 35980 25004 35989
rect 26240 35980 26292 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 6092 35776 6144 35828
rect 6828 35776 6880 35828
rect 7748 35819 7800 35828
rect 7748 35785 7757 35819
rect 7757 35785 7791 35819
rect 7791 35785 7800 35819
rect 7748 35776 7800 35785
rect 8300 35776 8352 35828
rect 15752 35776 15804 35828
rect 22468 35819 22520 35828
rect 22468 35785 22477 35819
rect 22477 35785 22511 35819
rect 22511 35785 22520 35819
rect 22468 35776 22520 35785
rect 22836 35819 22888 35828
rect 22836 35785 22845 35819
rect 22845 35785 22879 35819
rect 22879 35785 22888 35819
rect 22836 35776 22888 35785
rect 24768 35776 24820 35828
rect 35624 35819 35676 35828
rect 35624 35785 35633 35819
rect 35633 35785 35667 35819
rect 35667 35785 35676 35819
rect 35624 35776 35676 35785
rect 15660 35751 15712 35760
rect 15660 35717 15669 35751
rect 15669 35717 15703 35751
rect 15703 35717 15712 35751
rect 15660 35708 15712 35717
rect 20168 35708 20220 35760
rect 22928 35708 22980 35760
rect 22008 35683 22060 35692
rect 22008 35649 22017 35683
rect 22017 35649 22051 35683
rect 22051 35649 22060 35683
rect 22008 35640 22060 35649
rect 26240 35640 26292 35692
rect 7104 35615 7156 35624
rect 7104 35581 7113 35615
rect 7113 35581 7147 35615
rect 7147 35581 7156 35615
rect 7104 35572 7156 35581
rect 14004 35572 14056 35624
rect 15384 35572 15436 35624
rect 15936 35572 15988 35624
rect 21732 35615 21784 35624
rect 21732 35581 21741 35615
rect 21741 35581 21775 35615
rect 21775 35581 21784 35615
rect 21732 35572 21784 35581
rect 23848 35572 23900 35624
rect 24952 35615 25004 35624
rect 24952 35581 24961 35615
rect 24961 35581 24995 35615
rect 24995 35581 25004 35615
rect 24952 35572 25004 35581
rect 26700 35615 26752 35624
rect 26700 35581 26709 35615
rect 26709 35581 26743 35615
rect 26743 35581 26752 35615
rect 26700 35572 26752 35581
rect 34520 35572 34572 35624
rect 8852 35547 8904 35556
rect 8852 35513 8861 35547
rect 8861 35513 8895 35547
rect 8895 35513 8904 35547
rect 8852 35504 8904 35513
rect 15844 35504 15896 35556
rect 6092 35479 6144 35488
rect 6092 35445 6101 35479
rect 6101 35445 6135 35479
rect 6135 35445 6144 35479
rect 6092 35436 6144 35445
rect 7288 35479 7340 35488
rect 7288 35445 7297 35479
rect 7297 35445 7331 35479
rect 7331 35445 7340 35479
rect 7288 35436 7340 35445
rect 12256 35436 12308 35488
rect 15384 35436 15436 35488
rect 20904 35479 20956 35488
rect 20904 35445 20913 35479
rect 20913 35445 20947 35479
rect 20947 35445 20956 35479
rect 20904 35436 20956 35445
rect 21088 35436 21140 35488
rect 26516 35504 26568 35556
rect 23572 35436 23624 35488
rect 25136 35479 25188 35488
rect 25136 35445 25145 35479
rect 25145 35445 25179 35479
rect 25179 35445 25188 35479
rect 25136 35436 25188 35445
rect 26332 35479 26384 35488
rect 26332 35445 26341 35479
rect 26341 35445 26375 35479
rect 26375 35445 26384 35479
rect 26332 35436 26384 35445
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 1676 35232 1728 35284
rect 4988 35232 5040 35284
rect 7104 35275 7156 35284
rect 7104 35241 7113 35275
rect 7113 35241 7147 35275
rect 7147 35241 7156 35275
rect 7104 35232 7156 35241
rect 12532 35232 12584 35284
rect 14004 35232 14056 35284
rect 14740 35275 14792 35284
rect 14740 35241 14749 35275
rect 14749 35241 14783 35275
rect 14783 35241 14792 35275
rect 14740 35232 14792 35241
rect 15292 35275 15344 35284
rect 15292 35241 15301 35275
rect 15301 35241 15335 35275
rect 15335 35241 15344 35275
rect 15292 35232 15344 35241
rect 20260 35232 20312 35284
rect 20904 35232 20956 35284
rect 22008 35232 22060 35284
rect 22836 35232 22888 35284
rect 23480 35275 23532 35284
rect 23480 35241 23489 35275
rect 23489 35241 23523 35275
rect 23523 35241 23532 35275
rect 23480 35232 23532 35241
rect 24952 35232 25004 35284
rect 25044 35232 25096 35284
rect 26332 35232 26384 35284
rect 35532 35275 35584 35284
rect 35532 35241 35541 35275
rect 35541 35241 35575 35275
rect 35575 35241 35584 35275
rect 35532 35232 35584 35241
rect 9496 35164 9548 35216
rect 10692 35164 10744 35216
rect 22468 35164 22520 35216
rect 1400 35139 1452 35148
rect 1400 35105 1409 35139
rect 1409 35105 1443 35139
rect 1443 35105 1452 35139
rect 1400 35096 1452 35105
rect 4712 35096 4764 35148
rect 5172 35096 5224 35148
rect 9128 35096 9180 35148
rect 9864 35139 9916 35148
rect 9864 35105 9873 35139
rect 9873 35105 9907 35139
rect 9907 35105 9916 35139
rect 9864 35096 9916 35105
rect 11796 35139 11848 35148
rect 11796 35105 11830 35139
rect 11830 35105 11848 35139
rect 11796 35096 11848 35105
rect 14188 35096 14240 35148
rect 14648 35096 14700 35148
rect 17224 35139 17276 35148
rect 17224 35105 17233 35139
rect 17233 35105 17267 35139
rect 17267 35105 17276 35139
rect 17224 35096 17276 35105
rect 19156 35096 19208 35148
rect 20996 35139 21048 35148
rect 20996 35105 21005 35139
rect 21005 35105 21039 35139
rect 21039 35105 21048 35139
rect 20996 35096 21048 35105
rect 26148 35096 26200 35148
rect 35716 35096 35768 35148
rect 11520 35071 11572 35080
rect 11520 35037 11529 35071
rect 11529 35037 11563 35071
rect 11563 35037 11572 35071
rect 11520 35028 11572 35037
rect 15752 35071 15804 35080
rect 15752 35037 15761 35071
rect 15761 35037 15795 35071
rect 15795 35037 15804 35071
rect 15752 35028 15804 35037
rect 15844 35071 15896 35080
rect 15844 35037 15853 35071
rect 15853 35037 15887 35071
rect 15887 35037 15896 35071
rect 17316 35071 17368 35080
rect 15844 35028 15896 35037
rect 17316 35037 17325 35071
rect 17325 35037 17359 35071
rect 17359 35037 17368 35071
rect 17316 35028 17368 35037
rect 16856 35003 16908 35012
rect 16856 34969 16865 35003
rect 16865 34969 16899 35003
rect 16899 34969 16908 35003
rect 16856 34960 16908 34969
rect 17040 34960 17092 35012
rect 18696 34960 18748 35012
rect 5908 34892 5960 34944
rect 6644 34935 6696 34944
rect 6644 34901 6653 34935
rect 6653 34901 6687 34935
rect 6687 34901 6696 34935
rect 6644 34892 6696 34901
rect 7472 34935 7524 34944
rect 7472 34901 7481 34935
rect 7481 34901 7515 34935
rect 7515 34901 7524 34935
rect 7472 34892 7524 34901
rect 8300 34892 8352 34944
rect 9680 34892 9732 34944
rect 10324 34935 10376 34944
rect 10324 34901 10333 34935
rect 10333 34901 10367 34935
rect 10367 34901 10376 34935
rect 10324 34892 10376 34901
rect 12808 34892 12860 34944
rect 13820 34892 13872 34944
rect 18052 34892 18104 34944
rect 20904 34892 20956 34944
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 23572 34960 23624 35012
rect 26424 35028 26476 35080
rect 24032 34935 24084 34944
rect 24032 34901 24041 34935
rect 24041 34901 24075 34935
rect 24075 34901 24084 34935
rect 24032 34892 24084 34901
rect 26516 34892 26568 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 572 34688 624 34740
rect 2044 34731 2096 34740
rect 2044 34697 2053 34731
rect 2053 34697 2087 34731
rect 2087 34697 2096 34731
rect 2044 34688 2096 34697
rect 3884 34688 3936 34740
rect 2688 34663 2740 34672
rect 2688 34629 2697 34663
rect 2697 34629 2731 34663
rect 2731 34629 2740 34663
rect 2688 34620 2740 34629
rect 3148 34595 3200 34604
rect 2044 34484 2096 34536
rect 3148 34561 3157 34595
rect 3157 34561 3191 34595
rect 3191 34561 3200 34595
rect 3148 34552 3200 34561
rect 4620 34688 4672 34740
rect 9128 34731 9180 34740
rect 9128 34697 9137 34731
rect 9137 34697 9171 34731
rect 9171 34697 9180 34731
rect 9128 34688 9180 34697
rect 9496 34731 9548 34740
rect 9496 34697 9505 34731
rect 9505 34697 9539 34731
rect 9539 34697 9548 34731
rect 9496 34688 9548 34697
rect 9864 34688 9916 34740
rect 11796 34688 11848 34740
rect 12440 34688 12492 34740
rect 14188 34731 14240 34740
rect 14188 34697 14197 34731
rect 14197 34697 14231 34731
rect 14231 34697 14240 34731
rect 14188 34688 14240 34697
rect 14648 34731 14700 34740
rect 14648 34697 14657 34731
rect 14657 34697 14691 34731
rect 14691 34697 14700 34731
rect 14648 34688 14700 34697
rect 15844 34688 15896 34740
rect 5448 34620 5500 34672
rect 8852 34620 8904 34672
rect 14280 34620 14332 34672
rect 15752 34620 15804 34672
rect 4712 34552 4764 34604
rect 6092 34552 6144 34604
rect 7288 34552 7340 34604
rect 10140 34595 10192 34604
rect 10140 34561 10149 34595
rect 10149 34561 10183 34595
rect 10183 34561 10192 34595
rect 10140 34552 10192 34561
rect 12348 34552 12400 34604
rect 14740 34595 14792 34604
rect 5908 34484 5960 34536
rect 7472 34484 7524 34536
rect 8392 34484 8444 34536
rect 9772 34484 9824 34536
rect 12532 34527 12584 34536
rect 12532 34493 12541 34527
rect 12541 34493 12575 34527
rect 12575 34493 12584 34527
rect 12532 34484 12584 34493
rect 14740 34561 14749 34595
rect 14749 34561 14783 34595
rect 14783 34561 14792 34595
rect 14740 34552 14792 34561
rect 17224 34688 17276 34740
rect 19156 34731 19208 34740
rect 19156 34697 19165 34731
rect 19165 34697 19199 34731
rect 19199 34697 19208 34731
rect 19156 34688 19208 34697
rect 20996 34731 21048 34740
rect 20996 34697 21005 34731
rect 21005 34697 21039 34731
rect 21039 34697 21048 34731
rect 20996 34688 21048 34697
rect 22468 34688 22520 34740
rect 25044 34688 25096 34740
rect 26148 34731 26200 34740
rect 26148 34697 26157 34731
rect 26157 34697 26191 34731
rect 26191 34697 26200 34731
rect 26148 34688 26200 34697
rect 26516 34731 26568 34740
rect 26516 34697 26525 34731
rect 26525 34697 26559 34731
rect 26559 34697 26568 34731
rect 26516 34688 26568 34697
rect 26792 34688 26844 34740
rect 35808 34688 35860 34740
rect 36728 34731 36780 34740
rect 36728 34697 36737 34731
rect 36737 34697 36771 34731
rect 36771 34697 36780 34731
rect 36728 34688 36780 34697
rect 18144 34620 18196 34672
rect 20536 34620 20588 34672
rect 17960 34552 18012 34604
rect 18696 34595 18748 34604
rect 12808 34527 12860 34536
rect 12808 34493 12842 34527
rect 12842 34493 12860 34527
rect 12808 34484 12860 34493
rect 17684 34484 17736 34536
rect 18696 34561 18705 34595
rect 18705 34561 18739 34595
rect 18739 34561 18748 34595
rect 18696 34552 18748 34561
rect 19156 34552 19208 34604
rect 20076 34552 20128 34604
rect 9312 34416 9364 34468
rect 10324 34416 10376 34468
rect 14280 34416 14332 34468
rect 20260 34484 20312 34536
rect 20904 34484 20956 34536
rect 21732 34484 21784 34536
rect 20168 34416 20220 34468
rect 24032 34484 24084 34536
rect 26608 34527 26660 34536
rect 22284 34416 22336 34468
rect 26608 34493 26617 34527
rect 26617 34493 26651 34527
rect 26651 34493 26660 34527
rect 26608 34484 26660 34493
rect 35532 34484 35584 34536
rect 35716 34484 35768 34536
rect 37096 34527 37148 34536
rect 37096 34493 37105 34527
rect 37105 34493 37139 34527
rect 37139 34493 37148 34527
rect 37096 34484 37148 34493
rect 25044 34416 25096 34468
rect 5172 34348 5224 34400
rect 5632 34391 5684 34400
rect 5632 34357 5641 34391
rect 5641 34357 5675 34391
rect 5675 34357 5684 34391
rect 6276 34391 6328 34400
rect 5632 34348 5684 34357
rect 6276 34357 6285 34391
rect 6285 34357 6319 34391
rect 6319 34357 6328 34391
rect 6276 34348 6328 34357
rect 7196 34391 7248 34400
rect 7196 34357 7205 34391
rect 7205 34357 7239 34391
rect 7239 34357 7248 34391
rect 7196 34348 7248 34357
rect 9588 34391 9640 34400
rect 9588 34357 9597 34391
rect 9597 34357 9631 34391
rect 9631 34357 9640 34391
rect 9588 34348 9640 34357
rect 11152 34391 11204 34400
rect 11152 34357 11161 34391
rect 11161 34357 11195 34391
rect 11195 34357 11204 34391
rect 11152 34348 11204 34357
rect 28632 34348 28684 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 5632 34187 5684 34196
rect 5632 34153 5641 34187
rect 5641 34153 5675 34187
rect 5675 34153 5684 34187
rect 5632 34144 5684 34153
rect 5724 34144 5776 34196
rect 6092 34144 6144 34196
rect 1400 34076 1452 34128
rect 2872 34076 2924 34128
rect 6644 34076 6696 34128
rect 5172 34008 5224 34060
rect 5816 34008 5868 34060
rect 9588 34144 9640 34196
rect 12440 34144 12492 34196
rect 12992 34144 13044 34196
rect 14004 34187 14056 34196
rect 14004 34153 14013 34187
rect 14013 34153 14047 34187
rect 14047 34153 14056 34187
rect 14004 34144 14056 34153
rect 14648 34144 14700 34196
rect 20076 34187 20128 34196
rect 20076 34153 20085 34187
rect 20085 34153 20119 34187
rect 20119 34153 20128 34187
rect 20076 34144 20128 34153
rect 22284 34187 22336 34196
rect 22284 34153 22293 34187
rect 22293 34153 22327 34187
rect 22327 34153 22336 34187
rect 22284 34144 22336 34153
rect 23572 34187 23624 34196
rect 23572 34153 23581 34187
rect 23581 34153 23615 34187
rect 23615 34153 23624 34187
rect 23572 34144 23624 34153
rect 25044 34187 25096 34196
rect 25044 34153 25053 34187
rect 25053 34153 25087 34187
rect 25087 34153 25096 34187
rect 25044 34144 25096 34153
rect 25780 34144 25832 34196
rect 26148 34144 26200 34196
rect 35440 34144 35492 34196
rect 10140 34076 10192 34128
rect 18144 34076 18196 34128
rect 20168 34076 20220 34128
rect 23480 34076 23532 34128
rect 24032 34076 24084 34128
rect 26700 34076 26752 34128
rect 11520 34051 11572 34060
rect 4712 33940 4764 33992
rect 3516 33872 3568 33924
rect 5540 33940 5592 33992
rect 5908 33940 5960 33992
rect 9404 33940 9456 33992
rect 11520 34017 11529 34051
rect 11529 34017 11563 34051
rect 11563 34017 11572 34051
rect 11520 34008 11572 34017
rect 11796 34008 11848 34060
rect 14924 34008 14976 34060
rect 15384 34008 15436 34060
rect 20996 34008 21048 34060
rect 22744 34008 22796 34060
rect 35256 34008 35308 34060
rect 14740 33940 14792 33992
rect 2964 33847 3016 33856
rect 2964 33813 2973 33847
rect 2973 33813 3007 33847
rect 3007 33813 3016 33847
rect 2964 33804 3016 33813
rect 4068 33804 4120 33856
rect 7196 33804 7248 33856
rect 8668 33847 8720 33856
rect 8668 33813 8677 33847
rect 8677 33813 8711 33847
rect 8711 33813 8720 33847
rect 8668 33804 8720 33813
rect 11060 33847 11112 33856
rect 11060 33813 11069 33847
rect 11069 33813 11103 33847
rect 11103 33813 11112 33847
rect 11060 33804 11112 33813
rect 14280 33804 14332 33856
rect 20628 33940 20680 33992
rect 20904 33983 20956 33992
rect 20904 33949 20913 33983
rect 20913 33949 20947 33983
rect 20947 33949 20956 33983
rect 20904 33940 20956 33949
rect 26608 33940 26660 33992
rect 16212 33804 16264 33856
rect 16672 33847 16724 33856
rect 16672 33813 16681 33847
rect 16681 33813 16715 33847
rect 16715 33813 16724 33847
rect 16672 33804 16724 33813
rect 17040 33847 17092 33856
rect 17040 33813 17049 33847
rect 17049 33813 17083 33847
rect 17083 33813 17092 33847
rect 17040 33804 17092 33813
rect 17316 33804 17368 33856
rect 17776 33804 17828 33856
rect 19156 33847 19208 33856
rect 19156 33813 19165 33847
rect 19165 33813 19199 33847
rect 19199 33813 19208 33847
rect 19156 33804 19208 33813
rect 25872 33847 25924 33856
rect 25872 33813 25881 33847
rect 25881 33813 25915 33847
rect 25915 33813 25924 33847
rect 25872 33804 25924 33813
rect 26240 33804 26292 33856
rect 26792 33847 26844 33856
rect 26792 33813 26801 33847
rect 26801 33813 26835 33847
rect 26835 33813 26844 33847
rect 26792 33804 26844 33813
rect 28264 33847 28316 33856
rect 28264 33813 28273 33847
rect 28273 33813 28307 33847
rect 28307 33813 28316 33847
rect 28264 33804 28316 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 5816 33643 5868 33652
rect 5816 33609 5825 33643
rect 5825 33609 5859 33643
rect 5859 33609 5868 33643
rect 5816 33600 5868 33609
rect 6276 33600 6328 33652
rect 10140 33600 10192 33652
rect 15936 33600 15988 33652
rect 17040 33600 17092 33652
rect 18328 33600 18380 33652
rect 19248 33600 19300 33652
rect 20996 33600 21048 33652
rect 22744 33643 22796 33652
rect 6644 33532 6696 33584
rect 10784 33575 10836 33584
rect 10784 33541 10793 33575
rect 10793 33541 10827 33575
rect 10827 33541 10836 33575
rect 10784 33532 10836 33541
rect 3516 33507 3568 33516
rect 3516 33473 3525 33507
rect 3525 33473 3559 33507
rect 3559 33473 3568 33507
rect 3516 33464 3568 33473
rect 7380 33507 7432 33516
rect 7380 33473 7389 33507
rect 7389 33473 7423 33507
rect 7423 33473 7432 33507
rect 7380 33464 7432 33473
rect 2964 33396 3016 33448
rect 4068 33396 4120 33448
rect 5908 33396 5960 33448
rect 6828 33396 6880 33448
rect 8392 33396 8444 33448
rect 11060 33464 11112 33516
rect 11796 33507 11848 33516
rect 11796 33473 11805 33507
rect 11805 33473 11839 33507
rect 11839 33473 11848 33507
rect 11796 33464 11848 33473
rect 12992 33507 13044 33516
rect 12992 33473 13001 33507
rect 13001 33473 13035 33507
rect 13035 33473 13044 33507
rect 12992 33464 13044 33473
rect 15108 33464 15160 33516
rect 15936 33507 15988 33516
rect 15936 33473 15945 33507
rect 15945 33473 15979 33507
rect 15979 33473 15988 33507
rect 15936 33464 15988 33473
rect 22744 33609 22753 33643
rect 22753 33609 22787 33643
rect 22787 33609 22796 33643
rect 22744 33600 22796 33609
rect 23480 33643 23532 33652
rect 23480 33609 23489 33643
rect 23489 33609 23523 33643
rect 23523 33609 23532 33643
rect 23480 33600 23532 33609
rect 25044 33600 25096 33652
rect 8852 33439 8904 33448
rect 8852 33405 8886 33439
rect 8886 33405 8904 33439
rect 8852 33396 8904 33405
rect 11152 33439 11204 33448
rect 11152 33405 11161 33439
rect 11161 33405 11195 33439
rect 11195 33405 11204 33439
rect 11152 33396 11204 33405
rect 11244 33439 11296 33448
rect 11244 33405 11253 33439
rect 11253 33405 11287 33439
rect 11287 33405 11296 33439
rect 12808 33439 12860 33448
rect 11244 33396 11296 33405
rect 12808 33405 12817 33439
rect 12817 33405 12851 33439
rect 12851 33405 12860 33439
rect 12808 33396 12860 33405
rect 4712 33371 4764 33380
rect 4712 33337 4746 33371
rect 4746 33337 4764 33371
rect 4712 33328 4764 33337
rect 6644 33328 6696 33380
rect 12900 33371 12952 33380
rect 12900 33337 12909 33371
rect 12909 33337 12943 33371
rect 12943 33337 12952 33371
rect 12900 33328 12952 33337
rect 15568 33396 15620 33448
rect 18328 33371 18380 33380
rect 18328 33337 18362 33371
rect 18362 33337 18380 33371
rect 18328 33328 18380 33337
rect 1768 33303 1820 33312
rect 1768 33269 1777 33303
rect 1777 33269 1811 33303
rect 1811 33269 1820 33303
rect 1768 33260 1820 33269
rect 2872 33303 2924 33312
rect 2872 33269 2881 33303
rect 2881 33269 2915 33303
rect 2915 33269 2924 33303
rect 2872 33260 2924 33269
rect 3332 33303 3384 33312
rect 3332 33269 3341 33303
rect 3341 33269 3375 33303
rect 3375 33269 3384 33303
rect 3332 33260 3384 33269
rect 7196 33303 7248 33312
rect 7196 33269 7205 33303
rect 7205 33269 7239 33303
rect 7239 33269 7248 33303
rect 7196 33260 7248 33269
rect 12164 33260 12216 33312
rect 14188 33303 14240 33312
rect 14188 33269 14197 33303
rect 14197 33269 14231 33303
rect 14231 33269 14240 33303
rect 14188 33260 14240 33269
rect 15292 33260 15344 33312
rect 17040 33303 17092 33312
rect 17040 33269 17049 33303
rect 17049 33269 17083 33303
rect 17083 33269 17092 33303
rect 17040 33260 17092 33269
rect 18144 33260 18196 33312
rect 20168 33396 20220 33448
rect 20628 33439 20680 33448
rect 20628 33405 20637 33439
rect 20637 33405 20671 33439
rect 20671 33405 20680 33439
rect 20628 33396 20680 33405
rect 21824 33396 21876 33448
rect 24124 33532 24176 33584
rect 23572 33464 23624 33516
rect 24676 33464 24728 33516
rect 23388 33396 23440 33448
rect 21916 33328 21968 33380
rect 24124 33371 24176 33380
rect 24124 33337 24133 33371
rect 24133 33337 24167 33371
rect 24167 33337 24176 33371
rect 24124 33328 24176 33337
rect 19984 33260 20036 33312
rect 23480 33260 23532 33312
rect 25320 33600 25372 33652
rect 26700 33600 26752 33652
rect 35624 33643 35676 33652
rect 35624 33609 35633 33643
rect 35633 33609 35667 33643
rect 35667 33609 35676 33643
rect 35624 33600 35676 33609
rect 25964 33507 26016 33516
rect 25964 33473 25973 33507
rect 25973 33473 26007 33507
rect 26007 33473 26016 33507
rect 25964 33464 26016 33473
rect 35256 33464 35308 33516
rect 25780 33439 25832 33448
rect 25780 33405 25789 33439
rect 25789 33405 25823 33439
rect 25823 33405 25832 33439
rect 25780 33396 25832 33405
rect 26792 33396 26844 33448
rect 27068 33396 27120 33448
rect 28264 33396 28316 33448
rect 27160 33328 27212 33380
rect 28356 33303 28408 33312
rect 28356 33269 28365 33303
rect 28365 33269 28399 33303
rect 28399 33269 28408 33303
rect 28356 33260 28408 33269
rect 28632 33303 28684 33312
rect 28632 33269 28641 33303
rect 28641 33269 28675 33303
rect 28675 33269 28684 33303
rect 28632 33260 28684 33269
rect 35348 33303 35400 33312
rect 35348 33269 35357 33303
rect 35357 33269 35391 33303
rect 35391 33269 35400 33303
rect 35348 33260 35400 33269
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 2872 33056 2924 33108
rect 3792 33099 3844 33108
rect 3792 33065 3801 33099
rect 3801 33065 3835 33099
rect 3835 33065 3844 33099
rect 3792 33056 3844 33065
rect 4712 33056 4764 33108
rect 5540 33056 5592 33108
rect 6828 33056 6880 33108
rect 7196 33056 7248 33108
rect 8392 33056 8444 33108
rect 8668 33056 8720 33108
rect 10968 33056 11020 33108
rect 11244 33099 11296 33108
rect 11244 33065 11253 33099
rect 11253 33065 11287 33099
rect 11287 33065 11296 33099
rect 11244 33056 11296 33065
rect 12164 33056 12216 33108
rect 12808 33056 12860 33108
rect 13636 33099 13688 33108
rect 13636 33065 13645 33099
rect 13645 33065 13679 33099
rect 13679 33065 13688 33099
rect 13636 33056 13688 33065
rect 14924 33056 14976 33108
rect 15108 33099 15160 33108
rect 15108 33065 15117 33099
rect 15117 33065 15151 33099
rect 15151 33065 15160 33099
rect 15108 33056 15160 33065
rect 19340 33099 19392 33108
rect 19340 33065 19349 33099
rect 19349 33065 19383 33099
rect 19383 33065 19392 33099
rect 19340 33056 19392 33065
rect 22100 33056 22152 33108
rect 24676 33099 24728 33108
rect 24676 33065 24685 33099
rect 24685 33065 24719 33099
rect 24719 33065 24728 33099
rect 24676 33056 24728 33065
rect 24860 33099 24912 33108
rect 24860 33065 24869 33099
rect 24869 33065 24903 33099
rect 24903 33065 24912 33099
rect 24860 33056 24912 33065
rect 27068 33099 27120 33108
rect 27068 33065 27077 33099
rect 27077 33065 27111 33099
rect 27111 33065 27120 33099
rect 27068 33056 27120 33065
rect 5908 32988 5960 33040
rect 9404 33031 9456 33040
rect 9404 32997 9413 33031
rect 9413 32997 9447 33031
rect 9447 32997 9456 33031
rect 9404 32988 9456 32997
rect 12256 33031 12308 33040
rect 12256 32997 12265 33031
rect 12265 32997 12299 33031
rect 12299 32997 12308 33031
rect 12256 32988 12308 32997
rect 1860 32920 1912 32972
rect 3332 32920 3384 32972
rect 1768 32895 1820 32904
rect 1400 32716 1452 32768
rect 1768 32861 1777 32895
rect 1777 32861 1811 32895
rect 1811 32861 1820 32895
rect 1768 32852 1820 32861
rect 2964 32784 3016 32836
rect 7288 32920 7340 32972
rect 8392 32920 8444 32972
rect 9680 32963 9732 32972
rect 9680 32929 9689 32963
rect 9689 32929 9723 32963
rect 9723 32929 9732 32963
rect 9680 32920 9732 32929
rect 13268 32920 13320 32972
rect 15292 32963 15344 32972
rect 15292 32929 15301 32963
rect 15301 32929 15335 32963
rect 15335 32929 15344 32963
rect 15292 32920 15344 32929
rect 15568 32920 15620 32972
rect 16028 32963 16080 32972
rect 16028 32929 16037 32963
rect 16037 32929 16071 32963
rect 16071 32929 16080 32963
rect 16028 32920 16080 32929
rect 18236 32963 18288 32972
rect 18236 32929 18270 32963
rect 18270 32929 18288 32963
rect 18236 32920 18288 32929
rect 20628 32920 20680 32972
rect 22928 32920 22980 32972
rect 25228 32963 25280 32972
rect 4068 32895 4120 32904
rect 4068 32861 4077 32895
rect 4077 32861 4111 32895
rect 4111 32861 4120 32895
rect 4068 32852 4120 32861
rect 6276 32852 6328 32904
rect 7380 32852 7432 32904
rect 8208 32852 8260 32904
rect 12348 32852 12400 32904
rect 12532 32895 12584 32904
rect 12532 32861 12541 32895
rect 12541 32861 12575 32895
rect 12575 32861 12584 32895
rect 12532 32852 12584 32861
rect 14096 32895 14148 32904
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 14280 32895 14332 32904
rect 14280 32861 14289 32895
rect 14289 32861 14323 32895
rect 14323 32861 14332 32895
rect 14280 32852 14332 32861
rect 15752 32895 15804 32904
rect 15752 32861 15764 32895
rect 15764 32861 15798 32895
rect 15798 32861 15804 32895
rect 15752 32852 15804 32861
rect 16212 32852 16264 32904
rect 17592 32852 17644 32904
rect 23572 32895 23624 32904
rect 3516 32759 3568 32768
rect 3516 32725 3525 32759
rect 3525 32725 3559 32759
rect 3559 32725 3568 32759
rect 3516 32716 3568 32725
rect 3700 32716 3752 32768
rect 9588 32784 9640 32836
rect 11612 32784 11664 32836
rect 12624 32784 12676 32836
rect 7840 32716 7892 32768
rect 9864 32759 9916 32768
rect 9864 32725 9873 32759
rect 9873 32725 9907 32759
rect 9907 32725 9916 32759
rect 9864 32716 9916 32725
rect 11520 32716 11572 32768
rect 16764 32716 16816 32768
rect 18144 32716 18196 32768
rect 20168 32716 20220 32768
rect 23572 32861 23581 32895
rect 23581 32861 23615 32895
rect 23615 32861 23624 32895
rect 23572 32852 23624 32861
rect 25228 32929 25237 32963
rect 25237 32929 25271 32963
rect 25271 32929 25280 32963
rect 25228 32920 25280 32929
rect 25044 32852 25096 32904
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 27804 32988 27856 33040
rect 28356 32988 28408 33040
rect 27160 32963 27212 32972
rect 27160 32929 27169 32963
rect 27169 32929 27203 32963
rect 27203 32929 27212 32963
rect 27160 32920 27212 32929
rect 28632 32920 28684 32972
rect 29368 32963 29420 32972
rect 29368 32929 29377 32963
rect 29377 32929 29411 32963
rect 29411 32929 29420 32963
rect 29368 32920 29420 32929
rect 23388 32784 23440 32836
rect 21088 32716 21140 32768
rect 24124 32759 24176 32768
rect 24124 32725 24133 32759
rect 24133 32725 24167 32759
rect 24167 32725 24176 32759
rect 24124 32716 24176 32725
rect 28540 32759 28592 32768
rect 28540 32725 28549 32759
rect 28549 32725 28583 32759
rect 28583 32725 28592 32759
rect 28540 32716 28592 32725
rect 29552 32759 29604 32768
rect 29552 32725 29561 32759
rect 29561 32725 29595 32759
rect 29595 32725 29604 32759
rect 29552 32716 29604 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 1860 32512 1912 32564
rect 3332 32512 3384 32564
rect 5540 32555 5592 32564
rect 5540 32521 5549 32555
rect 5549 32521 5583 32555
rect 5583 32521 5592 32555
rect 5540 32512 5592 32521
rect 6276 32555 6328 32564
rect 6276 32521 6285 32555
rect 6285 32521 6319 32555
rect 6319 32521 6328 32555
rect 6276 32512 6328 32521
rect 2964 32444 3016 32496
rect 7288 32512 7340 32564
rect 7840 32555 7892 32564
rect 7840 32521 7849 32555
rect 7849 32521 7883 32555
rect 7883 32521 7892 32555
rect 7840 32512 7892 32521
rect 12164 32512 12216 32564
rect 12532 32512 12584 32564
rect 13268 32555 13320 32564
rect 13268 32521 13277 32555
rect 13277 32521 13311 32555
rect 13311 32521 13320 32555
rect 13268 32512 13320 32521
rect 14188 32555 14240 32564
rect 14188 32521 14197 32555
rect 14197 32521 14231 32555
rect 14231 32521 14240 32555
rect 14188 32512 14240 32521
rect 15108 32512 15160 32564
rect 15568 32512 15620 32564
rect 16212 32555 16264 32564
rect 16212 32521 16221 32555
rect 16221 32521 16255 32555
rect 16255 32521 16264 32555
rect 16212 32512 16264 32521
rect 20168 32555 20220 32564
rect 20168 32521 20177 32555
rect 20177 32521 20211 32555
rect 20211 32521 20220 32555
rect 20168 32512 20220 32521
rect 20628 32555 20680 32564
rect 20628 32521 20637 32555
rect 20637 32521 20671 32555
rect 20671 32521 20680 32555
rect 20628 32512 20680 32521
rect 23572 32512 23624 32564
rect 25228 32555 25280 32564
rect 25228 32521 25237 32555
rect 25237 32521 25271 32555
rect 25271 32521 25280 32555
rect 25228 32512 25280 32521
rect 25320 32512 25372 32564
rect 27804 32555 27856 32564
rect 27804 32521 27813 32555
rect 27813 32521 27847 32555
rect 27847 32521 27856 32555
rect 27804 32512 27856 32521
rect 28632 32555 28684 32564
rect 28632 32521 28641 32555
rect 28641 32521 28675 32555
rect 28675 32521 28684 32555
rect 28632 32512 28684 32521
rect 29368 32512 29420 32564
rect 8484 32444 8536 32496
rect 12256 32444 12308 32496
rect 15752 32487 15804 32496
rect 15752 32453 15761 32487
rect 15761 32453 15795 32487
rect 15795 32453 15804 32487
rect 15752 32444 15804 32453
rect 22100 32444 22152 32496
rect 3516 32376 3568 32428
rect 3976 32376 4028 32428
rect 5172 32376 5224 32428
rect 7380 32419 7432 32428
rect 7380 32385 7389 32419
rect 7389 32385 7423 32419
rect 7423 32385 7432 32419
rect 7380 32376 7432 32385
rect 8668 32376 8720 32428
rect 14096 32376 14148 32428
rect 14924 32419 14976 32428
rect 14924 32385 14933 32419
rect 14933 32385 14967 32419
rect 14967 32385 14976 32419
rect 14924 32376 14976 32385
rect 17684 32376 17736 32428
rect 21088 32419 21140 32428
rect 21088 32385 21097 32419
rect 21097 32385 21131 32419
rect 21131 32385 21140 32419
rect 21088 32376 21140 32385
rect 24216 32419 24268 32428
rect 24216 32385 24225 32419
rect 24225 32385 24259 32419
rect 24259 32385 24268 32419
rect 24216 32376 24268 32385
rect 25044 32376 25096 32428
rect 25872 32376 25924 32428
rect 27068 32376 27120 32428
rect 1400 32308 1452 32360
rect 3240 32308 3292 32360
rect 3700 32308 3752 32360
rect 3792 32308 3844 32360
rect 5540 32308 5592 32360
rect 7840 32308 7892 32360
rect 9680 32351 9732 32360
rect 9680 32317 9689 32351
rect 9689 32317 9723 32351
rect 9723 32317 9732 32351
rect 9680 32308 9732 32317
rect 14188 32308 14240 32360
rect 15108 32308 15160 32360
rect 16580 32308 16632 32360
rect 18144 32308 18196 32360
rect 18880 32308 18932 32360
rect 19984 32308 20036 32360
rect 20904 32308 20956 32360
rect 23296 32308 23348 32360
rect 24124 32308 24176 32360
rect 26884 32308 26936 32360
rect 27804 32308 27856 32360
rect 2780 32240 2832 32292
rect 3700 32172 3752 32224
rect 4068 32215 4120 32224
rect 4068 32181 4077 32215
rect 4077 32181 4111 32215
rect 4111 32181 4120 32215
rect 4068 32172 4120 32181
rect 4528 32215 4580 32224
rect 4528 32181 4537 32215
rect 4537 32181 4571 32215
rect 4571 32181 4580 32215
rect 4528 32172 4580 32181
rect 5540 32172 5592 32224
rect 8484 32240 8536 32292
rect 19156 32240 19208 32292
rect 7196 32215 7248 32224
rect 7196 32181 7205 32215
rect 7205 32181 7239 32215
rect 7239 32181 7248 32215
rect 7196 32172 7248 32181
rect 8392 32215 8444 32224
rect 8392 32181 8401 32215
rect 8401 32181 8435 32215
rect 8435 32181 8444 32215
rect 8392 32172 8444 32181
rect 18144 32172 18196 32224
rect 19432 32215 19484 32224
rect 19432 32181 19441 32215
rect 19441 32181 19475 32215
rect 19475 32181 19484 32215
rect 19432 32172 19484 32181
rect 20812 32172 20864 32224
rect 26240 32240 26292 32292
rect 23664 32215 23716 32224
rect 23664 32181 23673 32215
rect 23673 32181 23707 32215
rect 23707 32181 23716 32215
rect 23664 32172 23716 32181
rect 24124 32215 24176 32224
rect 24124 32181 24133 32215
rect 24133 32181 24167 32215
rect 24167 32181 24176 32215
rect 24124 32172 24176 32181
rect 26700 32172 26752 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 2780 32011 2832 32020
rect 2780 31977 2789 32011
rect 2789 31977 2823 32011
rect 2823 31977 2832 32011
rect 3240 32011 3292 32020
rect 2780 31968 2832 31977
rect 3240 31977 3249 32011
rect 3249 31977 3283 32011
rect 3283 31977 3292 32011
rect 3240 31968 3292 31977
rect 4528 31968 4580 32020
rect 5172 32011 5224 32020
rect 5172 31977 5181 32011
rect 5181 31977 5215 32011
rect 5215 31977 5224 32011
rect 5172 31968 5224 31977
rect 6276 31968 6328 32020
rect 7196 31968 7248 32020
rect 7288 32011 7340 32020
rect 7288 31977 7297 32011
rect 7297 31977 7331 32011
rect 7331 31977 7340 32011
rect 7288 31968 7340 31977
rect 8392 31968 8444 32020
rect 14280 31968 14332 32020
rect 15108 31968 15160 32020
rect 15568 31968 15620 32020
rect 17868 31968 17920 32020
rect 18880 32011 18932 32020
rect 18880 31977 18889 32011
rect 18889 31977 18923 32011
rect 18923 31977 18932 32011
rect 18880 31968 18932 31977
rect 20812 31968 20864 32020
rect 22928 31968 22980 32020
rect 24124 31968 24176 32020
rect 24216 32011 24268 32020
rect 24216 31977 24225 32011
rect 24225 31977 24259 32011
rect 24259 31977 24268 32011
rect 24216 31968 24268 31977
rect 25228 31968 25280 32020
rect 25872 32011 25924 32020
rect 25872 31977 25881 32011
rect 25881 31977 25915 32011
rect 25915 31977 25924 32011
rect 25872 31968 25924 31977
rect 26884 32011 26936 32020
rect 26884 31977 26893 32011
rect 26893 31977 26927 32011
rect 26927 31977 26936 32011
rect 26884 31968 26936 31977
rect 35808 31968 35860 32020
rect 3424 31900 3476 31952
rect 3700 31900 3752 31952
rect 7380 31900 7432 31952
rect 11060 31900 11112 31952
rect 14924 31900 14976 31952
rect 16028 31900 16080 31952
rect 21088 31900 21140 31952
rect 22008 31900 22060 31952
rect 25136 31900 25188 31952
rect 26700 31900 26752 31952
rect 28540 31900 28592 31952
rect 2504 31832 2556 31884
rect 4712 31832 4764 31884
rect 5632 31875 5684 31884
rect 5632 31841 5641 31875
rect 5641 31841 5675 31875
rect 5675 31841 5684 31875
rect 5632 31832 5684 31841
rect 8484 31875 8536 31884
rect 8484 31841 8493 31875
rect 8493 31841 8527 31875
rect 8527 31841 8536 31875
rect 8484 31832 8536 31841
rect 9404 31832 9456 31884
rect 11520 31832 11572 31884
rect 18144 31875 18196 31884
rect 18144 31841 18153 31875
rect 18153 31841 18187 31875
rect 18187 31841 18196 31875
rect 18144 31832 18196 31841
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 5172 31764 5224 31816
rect 4896 31696 4948 31748
rect 9312 31764 9364 31816
rect 9588 31764 9640 31816
rect 15292 31807 15344 31816
rect 15292 31773 15301 31807
rect 15301 31773 15335 31807
rect 15335 31773 15344 31807
rect 15292 31764 15344 31773
rect 18420 31832 18472 31884
rect 21640 31832 21692 31884
rect 23388 31832 23440 31884
rect 24768 31832 24820 31884
rect 25228 31875 25280 31884
rect 25228 31841 25237 31875
rect 25237 31841 25271 31875
rect 25271 31841 25280 31875
rect 25228 31832 25280 31841
rect 3700 31671 3752 31680
rect 3700 31637 3709 31671
rect 3709 31637 3743 31671
rect 3743 31637 3752 31671
rect 3700 31628 3752 31637
rect 17868 31696 17920 31748
rect 18052 31696 18104 31748
rect 20904 31764 20956 31816
rect 24216 31764 24268 31816
rect 26792 31832 26844 31884
rect 27160 31832 27212 31884
rect 35440 31875 35492 31884
rect 35440 31841 35449 31875
rect 35449 31841 35483 31875
rect 35483 31841 35492 31875
rect 35440 31832 35492 31841
rect 25504 31807 25556 31816
rect 25504 31773 25513 31807
rect 25513 31773 25547 31807
rect 25547 31773 25556 31807
rect 25504 31764 25556 31773
rect 18604 31696 18656 31748
rect 5724 31628 5776 31680
rect 5908 31628 5960 31680
rect 12348 31671 12400 31680
rect 12348 31637 12357 31671
rect 12357 31637 12391 31671
rect 12391 31637 12400 31671
rect 12348 31628 12400 31637
rect 24860 31671 24912 31680
rect 24860 31637 24869 31671
rect 24869 31637 24903 31671
rect 24903 31637 24912 31671
rect 24860 31628 24912 31637
rect 28448 31671 28500 31680
rect 28448 31637 28457 31671
rect 28457 31637 28491 31671
rect 28491 31637 28500 31671
rect 28448 31628 28500 31637
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 3424 31467 3476 31476
rect 3424 31433 3433 31467
rect 3433 31433 3467 31467
rect 3467 31433 3476 31467
rect 3424 31424 3476 31433
rect 4712 31467 4764 31476
rect 4712 31433 4721 31467
rect 4721 31433 4755 31467
rect 4755 31433 4764 31467
rect 4712 31424 4764 31433
rect 5632 31424 5684 31476
rect 7196 31424 7248 31476
rect 8484 31467 8536 31476
rect 8484 31433 8493 31467
rect 8493 31433 8527 31467
rect 8527 31433 8536 31467
rect 8484 31424 8536 31433
rect 8576 31424 8628 31476
rect 9404 31424 9456 31476
rect 10968 31424 11020 31476
rect 11888 31467 11940 31476
rect 11888 31433 11897 31467
rect 11897 31433 11931 31467
rect 11931 31433 11940 31467
rect 11888 31424 11940 31433
rect 2504 31356 2556 31408
rect 11520 31356 11572 31408
rect 1400 31331 1452 31340
rect 1400 31297 1409 31331
rect 1409 31297 1443 31331
rect 1443 31297 1452 31331
rect 1400 31288 1452 31297
rect 3976 31288 4028 31340
rect 5724 31331 5776 31340
rect 5724 31297 5733 31331
rect 5733 31297 5767 31331
rect 5767 31297 5776 31331
rect 5724 31288 5776 31297
rect 9220 31288 9272 31340
rect 9588 31288 9640 31340
rect 1676 31195 1728 31204
rect 1676 31161 1710 31195
rect 1710 31161 1728 31195
rect 1676 31152 1728 31161
rect 2964 31152 3016 31204
rect 3700 31152 3752 31204
rect 3608 31127 3660 31136
rect 3608 31093 3617 31127
rect 3617 31093 3651 31127
rect 3651 31093 3660 31127
rect 3608 31084 3660 31093
rect 4068 31127 4120 31136
rect 4068 31093 4077 31127
rect 4077 31093 4111 31127
rect 4111 31093 4120 31127
rect 4068 31084 4120 31093
rect 5080 31127 5132 31136
rect 5080 31093 5089 31127
rect 5089 31093 5123 31127
rect 5123 31093 5132 31127
rect 5080 31084 5132 31093
rect 8668 31220 8720 31272
rect 5264 31152 5316 31204
rect 9864 31195 9916 31204
rect 9864 31161 9873 31195
rect 9873 31161 9907 31195
rect 9907 31161 9916 31195
rect 9864 31152 9916 31161
rect 11152 31263 11204 31272
rect 11152 31229 11161 31263
rect 11161 31229 11195 31263
rect 11195 31229 11204 31263
rect 11152 31220 11204 31229
rect 11888 31220 11940 31272
rect 13912 31424 13964 31476
rect 16488 31467 16540 31476
rect 16488 31433 16497 31467
rect 16497 31433 16531 31467
rect 16531 31433 16540 31467
rect 16488 31424 16540 31433
rect 17040 31467 17092 31476
rect 17040 31433 17049 31467
rect 17049 31433 17083 31467
rect 17083 31433 17092 31467
rect 17040 31424 17092 31433
rect 17868 31467 17920 31476
rect 17868 31433 17877 31467
rect 17877 31433 17911 31467
rect 17911 31433 17920 31467
rect 17868 31424 17920 31433
rect 18604 31467 18656 31476
rect 18604 31433 18613 31467
rect 18613 31433 18647 31467
rect 18647 31433 18656 31467
rect 18604 31424 18656 31433
rect 20812 31467 20864 31476
rect 20812 31433 20821 31467
rect 20821 31433 20855 31467
rect 20855 31433 20864 31467
rect 20812 31424 20864 31433
rect 21824 31424 21876 31476
rect 23388 31467 23440 31476
rect 23388 31433 23397 31467
rect 23397 31433 23431 31467
rect 23431 31433 23440 31467
rect 23388 31424 23440 31433
rect 24768 31424 24820 31476
rect 25136 31424 25188 31476
rect 26240 31467 26292 31476
rect 26240 31433 26249 31467
rect 26249 31433 26283 31467
rect 26283 31433 26292 31467
rect 26240 31424 26292 31433
rect 26700 31467 26752 31476
rect 26700 31433 26709 31467
rect 26709 31433 26743 31467
rect 26743 31433 26752 31467
rect 26700 31424 26752 31433
rect 16580 31356 16632 31408
rect 13544 31263 13596 31272
rect 13544 31229 13553 31263
rect 13553 31229 13587 31263
rect 13587 31229 13596 31263
rect 13544 31220 13596 31229
rect 14372 31220 14424 31272
rect 15476 31263 15528 31272
rect 15476 31229 15485 31263
rect 15485 31229 15519 31263
rect 15519 31229 15528 31263
rect 15476 31220 15528 31229
rect 22008 31331 22060 31340
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 20812 31220 20864 31272
rect 26056 31356 26108 31408
rect 26608 31220 26660 31272
rect 26792 31263 26844 31272
rect 26792 31229 26801 31263
rect 26801 31229 26835 31263
rect 26835 31229 26844 31263
rect 26792 31220 26844 31229
rect 28448 31220 28500 31272
rect 5356 31084 5408 31136
rect 9588 31084 9640 31136
rect 9772 31127 9824 31136
rect 9772 31093 9781 31127
rect 9781 31093 9815 31127
rect 9815 31093 9824 31127
rect 9772 31084 9824 31093
rect 11336 31084 11388 31136
rect 13084 31084 13136 31136
rect 18144 31152 18196 31204
rect 21640 31152 21692 31204
rect 24768 31195 24820 31204
rect 24768 31161 24777 31195
rect 24777 31161 24811 31195
rect 24811 31161 24820 31195
rect 24768 31152 24820 31161
rect 25136 31084 25188 31136
rect 28172 31127 28224 31136
rect 28172 31093 28181 31127
rect 28181 31093 28215 31127
rect 28215 31093 28224 31127
rect 28172 31084 28224 31093
rect 35440 31127 35492 31136
rect 35440 31093 35449 31127
rect 35449 31093 35483 31127
rect 35483 31093 35492 31127
rect 35440 31084 35492 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 2504 30880 2556 30932
rect 2780 30880 2832 30932
rect 4068 30880 4120 30932
rect 5448 30880 5500 30932
rect 1400 30812 1452 30864
rect 6276 30812 6328 30864
rect 3608 30744 3660 30796
rect 3976 30744 4028 30796
rect 4896 30787 4948 30796
rect 4896 30753 4905 30787
rect 4905 30753 4939 30787
rect 4939 30753 4948 30787
rect 4896 30744 4948 30753
rect 5448 30744 5500 30796
rect 8668 30787 8720 30796
rect 8668 30753 8677 30787
rect 8677 30753 8711 30787
rect 8711 30753 8720 30787
rect 8668 30744 8720 30753
rect 9956 30744 10008 30796
rect 11520 30880 11572 30932
rect 12716 30923 12768 30932
rect 12716 30889 12725 30923
rect 12725 30889 12759 30923
rect 12759 30889 12768 30923
rect 12716 30880 12768 30889
rect 13084 30923 13136 30932
rect 13084 30889 13093 30923
rect 13093 30889 13127 30923
rect 13127 30889 13136 30923
rect 13084 30880 13136 30889
rect 13544 30923 13596 30932
rect 13544 30889 13553 30923
rect 13553 30889 13587 30923
rect 13587 30889 13596 30923
rect 13544 30880 13596 30889
rect 14372 30923 14424 30932
rect 14372 30889 14381 30923
rect 14381 30889 14415 30923
rect 14415 30889 14424 30923
rect 14372 30880 14424 30889
rect 17776 30923 17828 30932
rect 17776 30889 17785 30923
rect 17785 30889 17819 30923
rect 17819 30889 17828 30923
rect 17776 30880 17828 30889
rect 20904 30880 20956 30932
rect 21640 30880 21692 30932
rect 22008 30880 22060 30932
rect 23296 30880 23348 30932
rect 23940 30880 23992 30932
rect 24768 30923 24820 30932
rect 24768 30889 24777 30923
rect 24777 30889 24811 30923
rect 24811 30889 24820 30923
rect 24768 30880 24820 30889
rect 25504 30923 25556 30932
rect 25504 30889 25513 30923
rect 25513 30889 25547 30923
rect 25547 30889 25556 30923
rect 25504 30880 25556 30889
rect 35624 30923 35676 30932
rect 35624 30889 35633 30923
rect 35633 30889 35667 30923
rect 35667 30889 35676 30923
rect 35624 30880 35676 30889
rect 15568 30812 15620 30864
rect 5356 30719 5408 30728
rect 5356 30685 5365 30719
rect 5365 30685 5399 30719
rect 5399 30685 5408 30719
rect 5356 30676 5408 30685
rect 9772 30676 9824 30728
rect 10692 30676 10744 30728
rect 13728 30744 13780 30796
rect 14556 30787 14608 30796
rect 14556 30753 14565 30787
rect 14565 30753 14599 30787
rect 14599 30753 14608 30787
rect 14556 30744 14608 30753
rect 17040 30744 17092 30796
rect 18788 30744 18840 30796
rect 22560 30787 22612 30796
rect 22560 30753 22569 30787
rect 22569 30753 22603 30787
rect 22603 30753 22612 30787
rect 22560 30744 22612 30753
rect 25136 30744 25188 30796
rect 26516 30787 26568 30796
rect 26516 30753 26525 30787
rect 26525 30753 26559 30787
rect 26559 30753 26568 30787
rect 26516 30744 26568 30753
rect 35624 30744 35676 30796
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 7012 30651 7064 30660
rect 7012 30617 7021 30651
rect 7021 30617 7055 30651
rect 7055 30617 7064 30651
rect 7012 30608 7064 30617
rect 3056 30583 3108 30592
rect 3056 30549 3065 30583
rect 3065 30549 3099 30583
rect 3099 30549 3108 30583
rect 3056 30540 3108 30549
rect 5264 30583 5316 30592
rect 5264 30549 5273 30583
rect 5273 30549 5307 30583
rect 5307 30549 5316 30583
rect 5264 30540 5316 30549
rect 6736 30583 6788 30592
rect 6736 30549 6745 30583
rect 6745 30549 6779 30583
rect 6779 30549 6788 30583
rect 6736 30540 6788 30549
rect 8484 30583 8536 30592
rect 8484 30549 8493 30583
rect 8493 30549 8527 30583
rect 8527 30549 8536 30583
rect 8484 30540 8536 30549
rect 12900 30651 12952 30660
rect 12900 30617 12909 30651
rect 12909 30617 12943 30651
rect 12943 30617 12952 30651
rect 12900 30608 12952 30617
rect 17776 30676 17828 30728
rect 18328 30719 18380 30728
rect 18328 30685 18337 30719
rect 18337 30685 18371 30719
rect 18371 30685 18380 30719
rect 18328 30676 18380 30685
rect 23664 30676 23716 30728
rect 24124 30608 24176 30660
rect 11060 30540 11112 30592
rect 14280 30583 14332 30592
rect 14280 30549 14289 30583
rect 14289 30549 14323 30583
rect 14323 30549 14332 30583
rect 14280 30540 14332 30549
rect 16580 30540 16632 30592
rect 18880 30583 18932 30592
rect 18880 30549 18889 30583
rect 18889 30549 18923 30583
rect 18923 30549 18932 30583
rect 18880 30540 18932 30549
rect 24400 30583 24452 30592
rect 24400 30549 24409 30583
rect 24409 30549 24443 30583
rect 24443 30549 24452 30583
rect 24400 30540 24452 30549
rect 26608 30540 26660 30592
rect 33048 30540 33100 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 1400 30336 1452 30388
rect 2964 30379 3016 30388
rect 2964 30345 2973 30379
rect 2973 30345 3007 30379
rect 3007 30345 3016 30379
rect 2964 30336 3016 30345
rect 3976 30379 4028 30388
rect 3976 30345 3985 30379
rect 3985 30345 4019 30379
rect 4019 30345 4028 30379
rect 3976 30336 4028 30345
rect 2320 30268 2372 30320
rect 4896 30336 4948 30388
rect 5264 30336 5316 30388
rect 9864 30379 9916 30388
rect 9864 30345 9873 30379
rect 9873 30345 9907 30379
rect 9907 30345 9916 30379
rect 9864 30336 9916 30345
rect 13728 30379 13780 30388
rect 13728 30345 13737 30379
rect 13737 30345 13771 30379
rect 13771 30345 13780 30379
rect 13728 30336 13780 30345
rect 5908 30311 5960 30320
rect 5908 30277 5917 30311
rect 5917 30277 5951 30311
rect 5951 30277 5960 30311
rect 5908 30268 5960 30277
rect 10784 30311 10836 30320
rect 10784 30277 10793 30311
rect 10793 30277 10827 30311
rect 10827 30277 10836 30311
rect 10784 30268 10836 30277
rect 5540 30200 5592 30252
rect 6000 30200 6052 30252
rect 11428 30243 11480 30252
rect 11428 30209 11437 30243
rect 11437 30209 11471 30243
rect 11471 30209 11480 30243
rect 11428 30200 11480 30209
rect 13084 30200 13136 30252
rect 16488 30200 16540 30252
rect 17316 30200 17368 30252
rect 18880 30336 18932 30388
rect 21640 30336 21692 30388
rect 22560 30379 22612 30388
rect 22560 30345 22569 30379
rect 22569 30345 22603 30379
rect 22603 30345 22612 30379
rect 22560 30336 22612 30345
rect 24676 30379 24728 30388
rect 24676 30345 24685 30379
rect 24685 30345 24719 30379
rect 24719 30345 24728 30379
rect 24676 30336 24728 30345
rect 26516 30379 26568 30388
rect 26516 30345 26525 30379
rect 26525 30345 26559 30379
rect 26559 30345 26568 30379
rect 26516 30336 26568 30345
rect 18236 30200 18288 30252
rect 18788 30243 18840 30252
rect 18788 30209 18797 30243
rect 18797 30209 18831 30243
rect 18831 30209 18840 30243
rect 18788 30200 18840 30209
rect 35716 30268 35768 30320
rect 33048 30243 33100 30252
rect 3056 30132 3108 30184
rect 5356 30132 5408 30184
rect 6460 30132 6512 30184
rect 7012 30132 7064 30184
rect 8576 30132 8628 30184
rect 11060 30132 11112 30184
rect 12900 30132 12952 30184
rect 14188 30175 14240 30184
rect 14188 30141 14197 30175
rect 14197 30141 14231 30175
rect 14231 30141 14240 30175
rect 14188 30132 14240 30141
rect 14280 30132 14332 30184
rect 16764 30175 16816 30184
rect 16764 30141 16773 30175
rect 16773 30141 16807 30175
rect 16807 30141 16816 30175
rect 16764 30132 16816 30141
rect 18420 30132 18472 30184
rect 4068 30064 4120 30116
rect 6736 30064 6788 30116
rect 12440 30064 12492 30116
rect 15660 30064 15712 30116
rect 6276 30039 6328 30048
rect 6276 30005 6285 30039
rect 6285 30005 6319 30039
rect 6319 30005 6328 30039
rect 6276 29996 6328 30005
rect 8392 30039 8444 30048
rect 8392 30005 8401 30039
rect 8401 30005 8435 30039
rect 8435 30005 8444 30039
rect 8392 29996 8444 30005
rect 10232 30039 10284 30048
rect 10232 30005 10241 30039
rect 10241 30005 10275 30039
rect 10275 30005 10284 30039
rect 10232 29996 10284 30005
rect 10692 30039 10744 30048
rect 10692 30005 10701 30039
rect 10701 30005 10735 30039
rect 10735 30005 10744 30039
rect 10692 29996 10744 30005
rect 12624 30039 12676 30048
rect 12624 30005 12633 30039
rect 12633 30005 12667 30039
rect 12667 30005 12676 30039
rect 12624 29996 12676 30005
rect 12716 29996 12768 30048
rect 15568 30039 15620 30048
rect 15568 30005 15577 30039
rect 15577 30005 15611 30039
rect 15611 30005 15620 30039
rect 15568 29996 15620 30005
rect 16396 30039 16448 30048
rect 16396 30005 16405 30039
rect 16405 30005 16439 30039
rect 16439 30005 16448 30039
rect 16396 29996 16448 30005
rect 16580 29996 16632 30048
rect 17500 30039 17552 30048
rect 17500 30005 17509 30039
rect 17509 30005 17543 30039
rect 17543 30005 17552 30039
rect 17500 29996 17552 30005
rect 19156 29996 19208 30048
rect 20812 30132 20864 30184
rect 23664 30175 23716 30184
rect 23664 30141 23673 30175
rect 23673 30141 23707 30175
rect 23707 30141 23716 30175
rect 23664 30132 23716 30141
rect 24400 30132 24452 30184
rect 33048 30209 33057 30243
rect 33057 30209 33091 30243
rect 33091 30209 33100 30243
rect 33048 30200 33100 30209
rect 26976 30175 27028 30184
rect 24032 30064 24084 30116
rect 26976 30141 26985 30175
rect 26985 30141 27019 30175
rect 27019 30141 27028 30175
rect 26976 30132 27028 30141
rect 35716 30132 35768 30184
rect 20076 29996 20128 30048
rect 20536 30039 20588 30048
rect 20536 30005 20545 30039
rect 20545 30005 20579 30039
rect 20579 30005 20588 30039
rect 20536 29996 20588 30005
rect 23848 30039 23900 30048
rect 23848 30005 23857 30039
rect 23857 30005 23891 30039
rect 23891 30005 23900 30039
rect 23848 29996 23900 30005
rect 26148 30039 26200 30048
rect 26148 30005 26157 30039
rect 26157 30005 26191 30039
rect 26191 30005 26200 30039
rect 26148 29996 26200 30005
rect 27160 30039 27212 30048
rect 27160 30005 27169 30039
rect 27169 30005 27203 30039
rect 27203 30005 27212 30039
rect 27160 29996 27212 30005
rect 32220 30039 32272 30048
rect 32220 30005 32229 30039
rect 32229 30005 32263 30039
rect 32263 30005 32272 30039
rect 32220 29996 32272 30005
rect 32496 29996 32548 30048
rect 32772 30039 32824 30048
rect 32772 30005 32781 30039
rect 32781 30005 32815 30039
rect 32815 30005 32824 30039
rect 32772 29996 32824 30005
rect 35624 29996 35676 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 2320 29835 2372 29844
rect 2320 29801 2329 29835
rect 2329 29801 2363 29835
rect 2363 29801 2372 29835
rect 2320 29792 2372 29801
rect 2688 29792 2740 29844
rect 6000 29835 6052 29844
rect 6000 29801 6009 29835
rect 6009 29801 6043 29835
rect 6043 29801 6052 29835
rect 6000 29792 6052 29801
rect 6276 29792 6328 29844
rect 8576 29792 8628 29844
rect 10692 29792 10744 29844
rect 11428 29835 11480 29844
rect 11428 29801 11437 29835
rect 11437 29801 11471 29835
rect 11471 29801 11480 29835
rect 11428 29792 11480 29801
rect 14280 29792 14332 29844
rect 15660 29792 15712 29844
rect 17500 29835 17552 29844
rect 17500 29801 17509 29835
rect 17509 29801 17543 29835
rect 17543 29801 17552 29835
rect 17500 29792 17552 29801
rect 18788 29792 18840 29844
rect 20536 29792 20588 29844
rect 23848 29792 23900 29844
rect 24584 29792 24636 29844
rect 2780 29699 2832 29708
rect 2780 29665 2789 29699
rect 2789 29665 2823 29699
rect 2823 29665 2832 29699
rect 2780 29656 2832 29665
rect 2504 29588 2556 29640
rect 3056 29724 3108 29776
rect 4620 29724 4672 29776
rect 9864 29724 9916 29776
rect 12900 29724 12952 29776
rect 18144 29767 18196 29776
rect 18144 29733 18153 29767
rect 18153 29733 18187 29767
rect 18187 29733 18196 29767
rect 18144 29724 18196 29733
rect 24124 29767 24176 29776
rect 24124 29733 24133 29767
rect 24133 29733 24167 29767
rect 24167 29733 24176 29767
rect 24124 29724 24176 29733
rect 24400 29767 24452 29776
rect 24400 29733 24409 29767
rect 24409 29733 24443 29767
rect 24443 29733 24452 29767
rect 24400 29724 24452 29733
rect 24492 29724 24544 29776
rect 27160 29792 27212 29844
rect 35900 29835 35952 29844
rect 35900 29801 35909 29835
rect 35909 29801 35943 29835
rect 35943 29801 35952 29835
rect 35900 29792 35952 29801
rect 3884 29699 3936 29708
rect 3884 29665 3893 29699
rect 3893 29665 3927 29699
rect 3927 29665 3936 29699
rect 3884 29656 3936 29665
rect 5356 29656 5408 29708
rect 6552 29656 6604 29708
rect 8668 29656 8720 29708
rect 6460 29631 6512 29640
rect 6460 29597 6469 29631
rect 6469 29597 6503 29631
rect 6503 29597 6512 29631
rect 6460 29588 6512 29597
rect 7748 29588 7800 29640
rect 8484 29588 8536 29640
rect 9772 29656 9824 29708
rect 14188 29656 14240 29708
rect 15016 29656 15068 29708
rect 15384 29656 15436 29708
rect 16764 29656 16816 29708
rect 19616 29699 19668 29708
rect 19616 29665 19625 29699
rect 19625 29665 19659 29699
rect 19659 29665 19668 29699
rect 19616 29656 19668 29665
rect 20812 29656 20864 29708
rect 21180 29699 21232 29708
rect 21180 29665 21214 29699
rect 21214 29665 21232 29699
rect 21180 29656 21232 29665
rect 32772 29656 32824 29708
rect 33600 29656 33652 29708
rect 34520 29656 34572 29708
rect 35532 29656 35584 29708
rect 35808 29656 35860 29708
rect 11060 29588 11112 29640
rect 15476 29588 15528 29640
rect 15844 29588 15896 29640
rect 16304 29588 16356 29640
rect 19340 29588 19392 29640
rect 5632 29563 5684 29572
rect 5632 29529 5641 29563
rect 5641 29529 5675 29563
rect 5675 29529 5684 29563
rect 5632 29520 5684 29529
rect 19064 29520 19116 29572
rect 20536 29588 20588 29640
rect 25136 29631 25188 29640
rect 25136 29597 25145 29631
rect 25145 29597 25179 29631
rect 25179 29597 25188 29631
rect 25136 29588 25188 29597
rect 26148 29588 26200 29640
rect 26792 29588 26844 29640
rect 33508 29631 33560 29640
rect 33508 29597 33517 29631
rect 33517 29597 33551 29631
rect 33551 29597 33560 29631
rect 33508 29588 33560 29597
rect 12716 29452 12768 29504
rect 14004 29452 14056 29504
rect 14556 29452 14608 29504
rect 19248 29495 19300 29504
rect 19248 29461 19257 29495
rect 19257 29461 19291 29495
rect 19291 29461 19300 29495
rect 19248 29452 19300 29461
rect 24768 29452 24820 29504
rect 26148 29452 26200 29504
rect 27068 29495 27120 29504
rect 27068 29461 27077 29495
rect 27077 29461 27111 29495
rect 27111 29461 27120 29495
rect 27068 29452 27120 29461
rect 34704 29452 34756 29504
rect 35900 29452 35952 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 2504 29291 2556 29300
rect 2504 29257 2513 29291
rect 2513 29257 2547 29291
rect 2547 29257 2556 29291
rect 2504 29248 2556 29257
rect 4068 29291 4120 29300
rect 4068 29257 4077 29291
rect 4077 29257 4111 29291
rect 4111 29257 4120 29291
rect 4068 29248 4120 29257
rect 4620 29248 4672 29300
rect 5080 29248 5132 29300
rect 6552 29291 6604 29300
rect 6552 29257 6561 29291
rect 6561 29257 6595 29291
rect 6595 29257 6604 29291
rect 6552 29248 6604 29257
rect 9956 29291 10008 29300
rect 9956 29257 9965 29291
rect 9965 29257 9999 29291
rect 9999 29257 10008 29291
rect 9956 29248 10008 29257
rect 11336 29291 11388 29300
rect 11336 29257 11345 29291
rect 11345 29257 11379 29291
rect 11379 29257 11388 29291
rect 11336 29248 11388 29257
rect 11428 29248 11480 29300
rect 9864 29180 9916 29232
rect 5632 29155 5684 29164
rect 5632 29121 5641 29155
rect 5641 29121 5675 29155
rect 5675 29121 5684 29155
rect 5632 29112 5684 29121
rect 6000 29112 6052 29164
rect 6460 29112 6512 29164
rect 7748 29155 7800 29164
rect 7748 29121 7757 29155
rect 7757 29121 7791 29155
rect 7791 29121 7800 29155
rect 7748 29112 7800 29121
rect 10600 29155 10652 29164
rect 10600 29121 10609 29155
rect 10609 29121 10643 29155
rect 10643 29121 10652 29155
rect 12900 29248 12952 29300
rect 15660 29248 15712 29300
rect 16580 29248 16632 29300
rect 17316 29291 17368 29300
rect 17316 29257 17325 29291
rect 17325 29257 17359 29291
rect 17359 29257 17368 29291
rect 17316 29248 17368 29257
rect 17776 29291 17828 29300
rect 17776 29257 17785 29291
rect 17785 29257 17819 29291
rect 17819 29257 17828 29291
rect 17776 29248 17828 29257
rect 18420 29291 18472 29300
rect 18420 29257 18429 29291
rect 18429 29257 18463 29291
rect 18463 29257 18472 29291
rect 18420 29248 18472 29257
rect 19616 29248 19668 29300
rect 20812 29248 20864 29300
rect 21824 29291 21876 29300
rect 21824 29257 21833 29291
rect 21833 29257 21867 29291
rect 21867 29257 21876 29291
rect 21824 29248 21876 29257
rect 24584 29291 24636 29300
rect 24584 29257 24593 29291
rect 24593 29257 24627 29291
rect 24627 29257 24636 29291
rect 24584 29248 24636 29257
rect 26148 29291 26200 29300
rect 26148 29257 26157 29291
rect 26157 29257 26191 29291
rect 26191 29257 26200 29291
rect 26148 29248 26200 29257
rect 26424 29291 26476 29300
rect 26424 29257 26433 29291
rect 26433 29257 26467 29291
rect 26467 29257 26476 29291
rect 26424 29248 26476 29257
rect 26792 29291 26844 29300
rect 26792 29257 26801 29291
rect 26801 29257 26835 29291
rect 26835 29257 26844 29291
rect 26792 29248 26844 29257
rect 12440 29223 12492 29232
rect 12440 29189 12449 29223
rect 12449 29189 12483 29223
rect 12483 29189 12492 29223
rect 12440 29180 12492 29189
rect 15200 29180 15252 29232
rect 19156 29223 19208 29232
rect 19156 29189 19165 29223
rect 19165 29189 19199 29223
rect 19199 29189 19208 29223
rect 19156 29180 19208 29189
rect 21548 29180 21600 29232
rect 24216 29180 24268 29232
rect 24492 29180 24544 29232
rect 10600 29112 10652 29121
rect 13728 29112 13780 29164
rect 14280 29112 14332 29164
rect 15016 29112 15068 29164
rect 19248 29112 19300 29164
rect 20076 29155 20128 29164
rect 20076 29121 20085 29155
rect 20085 29121 20119 29155
rect 20119 29121 20128 29155
rect 20076 29112 20128 29121
rect 2044 29044 2096 29096
rect 5816 29044 5868 29096
rect 6276 29044 6328 29096
rect 9680 29044 9732 29096
rect 12716 29044 12768 29096
rect 15384 29044 15436 29096
rect 17316 29044 17368 29096
rect 18880 29044 18932 29096
rect 20352 29044 20404 29096
rect 20720 29044 20772 29096
rect 21180 29044 21232 29096
rect 21916 29044 21968 29096
rect 23940 29044 23992 29096
rect 24032 29044 24084 29096
rect 26884 29180 26936 29232
rect 34796 29180 34848 29232
rect 34980 29180 35032 29232
rect 35716 29180 35768 29232
rect 27068 29112 27120 29164
rect 35900 29112 35952 29164
rect 2780 28976 2832 29028
rect 8300 28976 8352 29028
rect 13820 29019 13872 29028
rect 13820 28985 13829 29019
rect 13829 28985 13863 29019
rect 13863 28985 13872 29019
rect 13820 28976 13872 28985
rect 19156 28976 19208 29028
rect 9128 28951 9180 28960
rect 9128 28917 9137 28951
rect 9137 28917 9171 28951
rect 9171 28917 9180 28951
rect 9128 28908 9180 28917
rect 10416 28951 10468 28960
rect 10416 28917 10425 28951
rect 10425 28917 10459 28951
rect 10459 28917 10468 28951
rect 10416 28908 10468 28917
rect 10968 28908 11020 28960
rect 14464 28951 14516 28960
rect 14464 28917 14473 28951
rect 14473 28917 14507 28951
rect 14507 28917 14516 28951
rect 21272 28976 21324 29028
rect 25136 28976 25188 29028
rect 14464 28908 14516 28917
rect 20536 28908 20588 28960
rect 24768 28908 24820 28960
rect 31484 29087 31536 29096
rect 31484 29053 31493 29087
rect 31493 29053 31527 29087
rect 31527 29053 31536 29087
rect 31484 29044 31536 29053
rect 35716 29044 35768 29096
rect 26424 28976 26476 29028
rect 25504 28908 25556 28960
rect 31208 28908 31260 28960
rect 33508 28976 33560 29028
rect 32680 28908 32732 28960
rect 33600 28951 33652 28960
rect 33600 28917 33609 28951
rect 33609 28917 33643 28951
rect 33643 28917 33652 28951
rect 33600 28908 33652 28917
rect 35808 28976 35860 29028
rect 34244 28908 34296 28960
rect 34704 28951 34756 28960
rect 34704 28917 34713 28951
rect 34713 28917 34747 28951
rect 34747 28917 34756 28951
rect 34704 28908 34756 28917
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 2780 28704 2832 28756
rect 3884 28747 3936 28756
rect 3884 28713 3893 28747
rect 3893 28713 3927 28747
rect 3927 28713 3936 28747
rect 3884 28704 3936 28713
rect 4620 28704 4672 28756
rect 5816 28747 5868 28756
rect 5816 28713 5825 28747
rect 5825 28713 5859 28747
rect 5859 28713 5868 28747
rect 5816 28704 5868 28713
rect 8300 28704 8352 28756
rect 10232 28704 10284 28756
rect 10600 28747 10652 28756
rect 10600 28713 10609 28747
rect 10609 28713 10643 28747
rect 10643 28713 10652 28747
rect 10600 28704 10652 28713
rect 14464 28704 14516 28756
rect 15292 28704 15344 28756
rect 19248 28747 19300 28756
rect 19248 28713 19257 28747
rect 19257 28713 19291 28747
rect 19291 28713 19300 28747
rect 19248 28704 19300 28713
rect 1860 28636 1912 28688
rect 2504 28636 2556 28688
rect 4160 28636 4212 28688
rect 12348 28636 12400 28688
rect 14280 28636 14332 28688
rect 15200 28636 15252 28688
rect 15844 28636 15896 28688
rect 19064 28679 19116 28688
rect 19064 28645 19073 28679
rect 19073 28645 19107 28679
rect 19107 28645 19116 28679
rect 19064 28636 19116 28645
rect 19524 28636 19576 28688
rect 20076 28704 20128 28756
rect 20812 28704 20864 28756
rect 22100 28704 22152 28756
rect 23664 28747 23716 28756
rect 23664 28713 23673 28747
rect 23673 28713 23707 28747
rect 23707 28713 23716 28747
rect 23664 28704 23716 28713
rect 24768 28704 24820 28756
rect 31208 28747 31260 28756
rect 31208 28713 31217 28747
rect 31217 28713 31251 28747
rect 31251 28713 31260 28747
rect 31208 28704 31260 28713
rect 33600 28704 33652 28756
rect 35716 28704 35768 28756
rect 7288 28568 7340 28620
rect 8392 28611 8444 28620
rect 8392 28577 8401 28611
rect 8401 28577 8435 28611
rect 8435 28577 8444 28611
rect 8392 28568 8444 28577
rect 9128 28568 9180 28620
rect 10232 28568 10284 28620
rect 12624 28568 12676 28620
rect 13452 28568 13504 28620
rect 21180 28611 21232 28620
rect 21180 28577 21214 28611
rect 21214 28577 21232 28611
rect 21180 28568 21232 28577
rect 26148 28636 26200 28688
rect 34152 28636 34204 28688
rect 34980 28636 35032 28688
rect 25596 28568 25648 28620
rect 27252 28568 27304 28620
rect 29920 28568 29972 28620
rect 32220 28568 32272 28620
rect 32680 28611 32732 28620
rect 32680 28577 32703 28611
rect 32703 28577 32732 28611
rect 32680 28568 32732 28577
rect 34704 28568 34756 28620
rect 8668 28543 8720 28552
rect 8668 28509 8677 28543
rect 8677 28509 8711 28543
rect 8711 28509 8720 28543
rect 8668 28500 8720 28509
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 9772 28500 9824 28552
rect 14648 28500 14700 28552
rect 15568 28500 15620 28552
rect 16856 28543 16908 28552
rect 16856 28509 16865 28543
rect 16865 28509 16899 28543
rect 16899 28509 16908 28543
rect 16856 28500 16908 28509
rect 19708 28543 19760 28552
rect 19708 28509 19717 28543
rect 19717 28509 19751 28543
rect 19751 28509 19760 28543
rect 19708 28500 19760 28509
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 20720 28500 20772 28552
rect 23848 28500 23900 28552
rect 26516 28543 26568 28552
rect 26516 28509 26525 28543
rect 26525 28509 26559 28543
rect 26559 28509 26568 28543
rect 26516 28500 26568 28509
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 29828 28500 29880 28509
rect 10416 28432 10468 28484
rect 16488 28432 16540 28484
rect 25504 28432 25556 28484
rect 2044 28364 2096 28416
rect 7840 28407 7892 28416
rect 7840 28373 7849 28407
rect 7849 28373 7883 28407
rect 7883 28373 7892 28407
rect 7840 28364 7892 28373
rect 12808 28364 12860 28416
rect 12992 28407 13044 28416
rect 12992 28373 13001 28407
rect 13001 28373 13035 28407
rect 13035 28373 13044 28407
rect 12992 28364 13044 28373
rect 15016 28364 15068 28416
rect 15384 28364 15436 28416
rect 16304 28407 16356 28416
rect 16304 28373 16313 28407
rect 16313 28373 16347 28407
rect 16347 28373 16356 28407
rect 16304 28364 16356 28373
rect 20352 28407 20404 28416
rect 20352 28373 20361 28407
rect 20361 28373 20395 28407
rect 20395 28373 20404 28407
rect 20352 28364 20404 28373
rect 20536 28364 20588 28416
rect 25596 28407 25648 28416
rect 25596 28373 25605 28407
rect 25605 28373 25639 28407
rect 25639 28373 25648 28407
rect 25596 28364 25648 28373
rect 27896 28407 27948 28416
rect 27896 28373 27905 28407
rect 27905 28373 27939 28407
rect 27939 28373 27948 28407
rect 27896 28364 27948 28373
rect 31484 28364 31536 28416
rect 34244 28364 34296 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 1860 28203 1912 28212
rect 1860 28169 1869 28203
rect 1869 28169 1903 28203
rect 1903 28169 1912 28203
rect 1860 28160 1912 28169
rect 4068 28160 4120 28212
rect 5356 28160 5408 28212
rect 7288 28203 7340 28212
rect 7288 28169 7297 28203
rect 7297 28169 7331 28203
rect 7331 28169 7340 28203
rect 7288 28160 7340 28169
rect 8300 28160 8352 28212
rect 10968 28160 11020 28212
rect 12348 28160 12400 28212
rect 13452 28203 13504 28212
rect 8668 28024 8720 28076
rect 9220 28024 9272 28076
rect 7564 27956 7616 28008
rect 11336 28067 11388 28076
rect 11336 28033 11345 28067
rect 11345 28033 11379 28067
rect 11379 28033 11388 28067
rect 13452 28169 13461 28203
rect 13461 28169 13495 28203
rect 13495 28169 13504 28203
rect 13452 28160 13504 28169
rect 14648 28203 14700 28212
rect 14648 28169 14657 28203
rect 14657 28169 14691 28203
rect 14691 28169 14700 28203
rect 14648 28160 14700 28169
rect 15292 28203 15344 28212
rect 15292 28169 15301 28203
rect 15301 28169 15335 28203
rect 15335 28169 15344 28203
rect 15292 28160 15344 28169
rect 16304 28160 16356 28212
rect 16396 28160 16448 28212
rect 19524 28160 19576 28212
rect 19708 28160 19760 28212
rect 19984 28160 20036 28212
rect 23848 28203 23900 28212
rect 23848 28169 23857 28203
rect 23857 28169 23891 28203
rect 23891 28169 23900 28203
rect 23848 28160 23900 28169
rect 27252 28203 27304 28212
rect 27252 28169 27261 28203
rect 27261 28169 27295 28203
rect 27295 28169 27304 28203
rect 27252 28160 27304 28169
rect 29920 28160 29972 28212
rect 32220 28203 32272 28212
rect 11336 28024 11388 28033
rect 12992 28067 13044 28076
rect 12992 28033 13001 28067
rect 13001 28033 13035 28067
rect 13035 28033 13044 28067
rect 19800 28092 19852 28144
rect 23756 28092 23808 28144
rect 12992 28024 13044 28033
rect 16488 28024 16540 28076
rect 19432 28024 19484 28076
rect 32220 28169 32229 28203
rect 32229 28169 32263 28203
rect 32263 28169 32272 28203
rect 32220 28160 32272 28169
rect 34704 28203 34756 28212
rect 34704 28169 34713 28203
rect 34713 28169 34747 28203
rect 34747 28169 34756 28203
rect 34704 28160 34756 28169
rect 12808 27999 12860 28008
rect 12808 27965 12817 27999
rect 12817 27965 12851 27999
rect 12851 27965 12860 27999
rect 12808 27956 12860 27965
rect 15568 27956 15620 28008
rect 16856 27956 16908 28008
rect 20812 27956 20864 28008
rect 23848 27956 23900 28008
rect 25412 27956 25464 28008
rect 32772 28024 32824 28076
rect 33048 28024 33100 28076
rect 33784 28024 33836 28076
rect 25872 27999 25924 28008
rect 25872 27965 25906 27999
rect 25906 27965 25924 27999
rect 25872 27956 25924 27965
rect 29828 27956 29880 28008
rect 7288 27888 7340 27940
rect 7840 27888 7892 27940
rect 15292 27888 15344 27940
rect 21824 27888 21876 27940
rect 26148 27888 26200 27940
rect 31024 27888 31076 27940
rect 31208 27956 31260 28008
rect 31484 27888 31536 27940
rect 2044 27820 2096 27872
rect 7564 27863 7616 27872
rect 7564 27829 7573 27863
rect 7573 27829 7607 27863
rect 7607 27829 7616 27863
rect 7564 27820 7616 27829
rect 7748 27863 7800 27872
rect 7748 27829 7757 27863
rect 7757 27829 7791 27863
rect 7791 27829 7800 27863
rect 7748 27820 7800 27829
rect 9220 27863 9272 27872
rect 9220 27829 9229 27863
rect 9229 27829 9263 27863
rect 9263 27829 9272 27863
rect 9220 27820 9272 27829
rect 10232 27863 10284 27872
rect 10232 27829 10241 27863
rect 10241 27829 10275 27863
rect 10275 27829 10284 27863
rect 10232 27820 10284 27829
rect 11152 27863 11204 27872
rect 11152 27829 11161 27863
rect 11161 27829 11195 27863
rect 11195 27829 11204 27863
rect 11152 27820 11204 27829
rect 21180 27820 21232 27872
rect 22100 27863 22152 27872
rect 22100 27829 22109 27863
rect 22109 27829 22143 27863
rect 22143 27829 22152 27863
rect 22100 27820 22152 27829
rect 24492 27863 24544 27872
rect 24492 27829 24501 27863
rect 24501 27829 24535 27863
rect 24535 27829 24544 27863
rect 24492 27820 24544 27829
rect 27068 27820 27120 27872
rect 32312 27863 32364 27872
rect 32312 27829 32321 27863
rect 32321 27829 32355 27863
rect 32355 27829 32364 27863
rect 32312 27820 32364 27829
rect 33968 27888 34020 27940
rect 34612 27888 34664 27940
rect 35072 27956 35124 28008
rect 35716 27956 35768 28008
rect 37464 27888 37516 27940
rect 33784 27863 33836 27872
rect 33784 27829 33793 27863
rect 33793 27829 33827 27863
rect 33827 27829 33836 27863
rect 33784 27820 33836 27829
rect 34244 27820 34296 27872
rect 34704 27820 34756 27872
rect 36360 27863 36412 27872
rect 36360 27829 36369 27863
rect 36369 27829 36403 27863
rect 36403 27829 36412 27863
rect 36360 27820 36412 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 2504 27616 2556 27668
rect 8300 27616 8352 27668
rect 9496 27659 9548 27668
rect 9496 27625 9505 27659
rect 9505 27625 9539 27659
rect 9539 27625 9548 27659
rect 9496 27616 9548 27625
rect 2044 27548 2096 27600
rect 1676 27523 1728 27532
rect 1676 27489 1710 27523
rect 1710 27489 1728 27523
rect 1676 27480 1728 27489
rect 6644 27480 6696 27532
rect 11152 27616 11204 27668
rect 12256 27616 12308 27668
rect 12348 27616 12400 27668
rect 12808 27616 12860 27668
rect 15568 27659 15620 27668
rect 15568 27625 15577 27659
rect 15577 27625 15611 27659
rect 15611 27625 15620 27659
rect 15568 27616 15620 27625
rect 15844 27659 15896 27668
rect 15844 27625 15853 27659
rect 15853 27625 15887 27659
rect 15887 27625 15896 27659
rect 15844 27616 15896 27625
rect 20812 27616 20864 27668
rect 24492 27616 24544 27668
rect 31024 27659 31076 27668
rect 31024 27625 31033 27659
rect 31033 27625 31067 27659
rect 31067 27625 31076 27659
rect 31024 27616 31076 27625
rect 32312 27616 32364 27668
rect 35072 27659 35124 27668
rect 35072 27625 35081 27659
rect 35081 27625 35115 27659
rect 35115 27625 35124 27659
rect 35072 27616 35124 27625
rect 21272 27591 21324 27600
rect 21272 27557 21281 27591
rect 21281 27557 21315 27591
rect 21315 27557 21324 27591
rect 21272 27548 21324 27557
rect 25412 27548 25464 27600
rect 26884 27548 26936 27600
rect 7288 27480 7340 27532
rect 9956 27523 10008 27532
rect 9956 27489 9965 27523
rect 9965 27489 9999 27523
rect 9999 27489 10008 27523
rect 9956 27480 10008 27489
rect 11060 27523 11112 27532
rect 11060 27489 11069 27523
rect 11069 27489 11103 27523
rect 11103 27489 11112 27523
rect 11060 27480 11112 27489
rect 11796 27480 11848 27532
rect 12348 27480 12400 27532
rect 12440 27480 12492 27532
rect 13452 27480 13504 27532
rect 16488 27523 16540 27532
rect 16488 27489 16497 27523
rect 16497 27489 16531 27523
rect 16531 27489 16540 27523
rect 16488 27480 16540 27489
rect 19340 27480 19392 27532
rect 22836 27523 22888 27532
rect 22836 27489 22845 27523
rect 22845 27489 22879 27523
rect 22879 27489 22888 27523
rect 22836 27480 22888 27489
rect 29460 27480 29512 27532
rect 29828 27548 29880 27600
rect 32496 27591 32548 27600
rect 32496 27557 32505 27591
rect 32505 27557 32539 27591
rect 32539 27557 32548 27591
rect 32496 27548 32548 27557
rect 32772 27548 32824 27600
rect 34612 27548 34664 27600
rect 35348 27548 35400 27600
rect 35900 27548 35952 27600
rect 37004 27548 37056 27600
rect 30840 27480 30892 27532
rect 34428 27480 34480 27532
rect 36360 27480 36412 27532
rect 19064 27412 19116 27464
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 10140 27387 10192 27396
rect 10140 27353 10149 27387
rect 10149 27353 10183 27387
rect 10183 27353 10192 27387
rect 10140 27344 10192 27353
rect 13728 27344 13780 27396
rect 18972 27344 19024 27396
rect 21088 27344 21140 27396
rect 22100 27412 22152 27464
rect 22652 27412 22704 27464
rect 23112 27455 23164 27464
rect 23112 27421 23121 27455
rect 23121 27421 23155 27455
rect 23155 27421 23164 27455
rect 23112 27412 23164 27421
rect 25320 27455 25372 27464
rect 25320 27421 25329 27455
rect 25329 27421 25363 27455
rect 25363 27421 25372 27455
rect 25320 27412 25372 27421
rect 25596 27412 25648 27464
rect 26516 27455 26568 27464
rect 26516 27421 26525 27455
rect 26525 27421 26559 27455
rect 26559 27421 26568 27455
rect 26516 27412 26568 27421
rect 33508 27412 33560 27464
rect 34704 27412 34756 27464
rect 12348 27276 12400 27328
rect 12900 27276 12952 27328
rect 15384 27276 15436 27328
rect 16672 27319 16724 27328
rect 16672 27285 16681 27319
rect 16681 27285 16715 27319
rect 16715 27285 16724 27319
rect 16672 27276 16724 27285
rect 20996 27276 21048 27328
rect 25596 27276 25648 27328
rect 27804 27276 27856 27328
rect 32128 27319 32180 27328
rect 32128 27285 32137 27319
rect 32137 27285 32171 27319
rect 32171 27285 32180 27319
rect 32128 27276 32180 27285
rect 33232 27319 33284 27328
rect 33232 27285 33241 27319
rect 33241 27285 33275 27319
rect 33275 27285 33284 27319
rect 33232 27276 33284 27285
rect 34244 27319 34296 27328
rect 34244 27285 34253 27319
rect 34253 27285 34287 27319
rect 34287 27285 34296 27319
rect 34244 27276 34296 27285
rect 36820 27319 36872 27328
rect 36820 27285 36829 27319
rect 36829 27285 36863 27319
rect 36863 27285 36872 27319
rect 36820 27276 36872 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 2044 27115 2096 27124
rect 2044 27081 2053 27115
rect 2053 27081 2087 27115
rect 2087 27081 2096 27115
rect 2044 27072 2096 27081
rect 6644 27115 6696 27124
rect 6644 27081 6653 27115
rect 6653 27081 6687 27115
rect 6687 27081 6696 27115
rect 6644 27072 6696 27081
rect 7748 27115 7800 27124
rect 7748 27081 7757 27115
rect 7757 27081 7791 27115
rect 7791 27081 7800 27115
rect 7748 27072 7800 27081
rect 8208 27115 8260 27124
rect 8208 27081 8217 27115
rect 8217 27081 8251 27115
rect 8251 27081 8260 27115
rect 8208 27072 8260 27081
rect 9956 27115 10008 27124
rect 9956 27081 9965 27115
rect 9965 27081 9999 27115
rect 9999 27081 10008 27115
rect 9956 27072 10008 27081
rect 11796 27115 11848 27124
rect 11796 27081 11805 27115
rect 11805 27081 11839 27115
rect 11839 27081 11848 27115
rect 11796 27072 11848 27081
rect 12256 27072 12308 27124
rect 13452 27115 13504 27124
rect 13452 27081 13461 27115
rect 13461 27081 13495 27115
rect 13495 27081 13504 27115
rect 13452 27072 13504 27081
rect 15292 27115 15344 27124
rect 15292 27081 15301 27115
rect 15301 27081 15335 27115
rect 15335 27081 15344 27115
rect 15292 27072 15344 27081
rect 16488 27072 16540 27124
rect 18512 27072 18564 27124
rect 19064 27072 19116 27124
rect 19340 27115 19392 27124
rect 19340 27081 19349 27115
rect 19349 27081 19383 27115
rect 19383 27081 19392 27115
rect 19340 27072 19392 27081
rect 21180 27072 21232 27124
rect 21824 27115 21876 27124
rect 21824 27081 21833 27115
rect 21833 27081 21867 27115
rect 21867 27081 21876 27115
rect 21824 27072 21876 27081
rect 23112 27072 23164 27124
rect 25412 27115 25464 27124
rect 25412 27081 25421 27115
rect 25421 27081 25455 27115
rect 25455 27081 25464 27115
rect 25412 27072 25464 27081
rect 27804 27115 27856 27124
rect 27804 27081 27813 27115
rect 27813 27081 27847 27115
rect 27847 27081 27856 27115
rect 27804 27072 27856 27081
rect 30840 27115 30892 27124
rect 30840 27081 30849 27115
rect 30849 27081 30883 27115
rect 30883 27081 30892 27115
rect 30840 27072 30892 27081
rect 31668 27115 31720 27124
rect 12900 27004 12952 27056
rect 8852 26979 8904 26988
rect 8852 26945 8861 26979
rect 8861 26945 8895 26979
rect 8895 26945 8904 26979
rect 8852 26936 8904 26945
rect 11336 26979 11388 26988
rect 11336 26945 11345 26979
rect 11345 26945 11379 26979
rect 11379 26945 11388 26979
rect 11336 26936 11388 26945
rect 12348 26936 12400 26988
rect 22100 27047 22152 27056
rect 22100 27013 22109 27047
rect 22109 27013 22143 27047
rect 22143 27013 22152 27047
rect 22100 27004 22152 27013
rect 7748 26868 7800 26920
rect 10968 26868 11020 26920
rect 11796 26868 11848 26920
rect 1676 26843 1728 26852
rect 1676 26809 1685 26843
rect 1685 26809 1719 26843
rect 1719 26809 1728 26843
rect 1676 26800 1728 26809
rect 2688 26800 2740 26852
rect 7288 26775 7340 26784
rect 7288 26741 7297 26775
rect 7297 26741 7331 26775
rect 7331 26741 7340 26775
rect 7288 26732 7340 26741
rect 7840 26732 7892 26784
rect 12348 26800 12400 26852
rect 15292 26868 15344 26920
rect 24584 26979 24636 26988
rect 24584 26945 24593 26979
rect 24593 26945 24627 26979
rect 24627 26945 24636 26979
rect 24584 26936 24636 26945
rect 31668 27081 31677 27115
rect 31677 27081 31711 27115
rect 31711 27081 31720 27115
rect 31668 27072 31720 27081
rect 32312 27072 32364 27124
rect 34428 27072 34480 27124
rect 34796 27072 34848 27124
rect 20996 26868 21048 26920
rect 25412 26868 25464 26920
rect 25596 26911 25648 26920
rect 25596 26877 25605 26911
rect 25605 26877 25639 26911
rect 25639 26877 25648 26911
rect 25596 26868 25648 26877
rect 27712 26868 27764 26920
rect 32772 26936 32824 26988
rect 33508 26936 33560 26988
rect 36360 27115 36412 27124
rect 36360 27081 36369 27115
rect 36369 27081 36403 27115
rect 36403 27081 36412 27115
rect 36360 27072 36412 27081
rect 37464 27115 37516 27124
rect 37464 27081 37473 27115
rect 37473 27081 37507 27115
rect 37507 27081 37516 27115
rect 37464 27072 37516 27081
rect 29552 26868 29604 26920
rect 33232 26868 33284 26920
rect 19892 26800 19944 26852
rect 20720 26843 20772 26852
rect 20720 26809 20754 26843
rect 20754 26809 20772 26843
rect 20720 26800 20772 26809
rect 22100 26800 22152 26852
rect 22836 26843 22888 26852
rect 22836 26809 22845 26843
rect 22845 26809 22879 26843
rect 22879 26809 22888 26843
rect 22836 26800 22888 26809
rect 11060 26775 11112 26784
rect 11060 26741 11069 26775
rect 11069 26741 11103 26775
rect 11103 26741 11112 26775
rect 11060 26732 11112 26741
rect 11796 26732 11848 26784
rect 12532 26732 12584 26784
rect 14004 26732 14056 26784
rect 14740 26775 14792 26784
rect 14740 26741 14749 26775
rect 14749 26741 14783 26775
rect 14783 26741 14792 26775
rect 14740 26732 14792 26741
rect 15936 26732 15988 26784
rect 22652 26732 22704 26784
rect 25320 26800 25372 26852
rect 24032 26775 24084 26784
rect 24032 26741 24041 26775
rect 24041 26741 24075 26775
rect 24075 26741 24084 26775
rect 24400 26775 24452 26784
rect 24032 26732 24084 26741
rect 24400 26741 24409 26775
rect 24409 26741 24443 26775
rect 24443 26741 24452 26775
rect 24400 26732 24452 26741
rect 25872 26843 25924 26852
rect 25872 26809 25906 26843
rect 25906 26809 25924 26843
rect 25872 26800 25924 26809
rect 30840 26800 30892 26852
rect 36636 26936 36688 26988
rect 37004 26979 37056 26988
rect 37004 26945 37013 26979
rect 37013 26945 37047 26979
rect 37047 26945 37056 26979
rect 37004 26936 37056 26945
rect 36360 26868 36412 26920
rect 34980 26800 35032 26852
rect 25964 26732 26016 26784
rect 26056 26732 26108 26784
rect 32036 26775 32088 26784
rect 32036 26741 32045 26775
rect 32045 26741 32079 26775
rect 32079 26741 32088 26775
rect 32036 26732 32088 26741
rect 33048 26775 33100 26784
rect 33048 26741 33057 26775
rect 33057 26741 33091 26775
rect 33091 26741 33100 26775
rect 33048 26732 33100 26741
rect 33232 26775 33284 26784
rect 33232 26741 33241 26775
rect 33241 26741 33275 26775
rect 33275 26741 33284 26775
rect 33232 26732 33284 26741
rect 34428 26732 34480 26784
rect 36820 26775 36872 26784
rect 36820 26741 36829 26775
rect 36829 26741 36863 26775
rect 36863 26741 36872 26775
rect 36820 26732 36872 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 7288 26528 7340 26580
rect 8852 26528 8904 26580
rect 11336 26528 11388 26580
rect 15936 26571 15988 26580
rect 15936 26537 15945 26571
rect 15945 26537 15979 26571
rect 15979 26537 15988 26571
rect 15936 26528 15988 26537
rect 19064 26528 19116 26580
rect 6920 26460 6972 26512
rect 7564 26460 7616 26512
rect 8208 26460 8260 26512
rect 11060 26460 11112 26512
rect 12348 26460 12400 26512
rect 19156 26503 19208 26512
rect 19156 26469 19165 26503
rect 19165 26469 19199 26503
rect 19199 26469 19208 26503
rect 19984 26528 20036 26580
rect 20720 26528 20772 26580
rect 23940 26528 23992 26580
rect 24584 26528 24636 26580
rect 24952 26528 25004 26580
rect 19156 26460 19208 26469
rect 26516 26528 26568 26580
rect 30840 26571 30892 26580
rect 30840 26537 30849 26571
rect 30849 26537 30883 26571
rect 30883 26537 30892 26571
rect 30840 26528 30892 26537
rect 31024 26528 31076 26580
rect 32036 26528 32088 26580
rect 33048 26528 33100 26580
rect 34980 26571 35032 26580
rect 34980 26537 34989 26571
rect 34989 26537 35023 26571
rect 35023 26537 35032 26571
rect 34980 26528 35032 26537
rect 32680 26460 32732 26512
rect 33784 26460 33836 26512
rect 7012 26392 7064 26444
rect 11796 26392 11848 26444
rect 15844 26435 15896 26444
rect 15844 26401 15853 26435
rect 15853 26401 15887 26435
rect 15887 26401 15896 26435
rect 15844 26392 15896 26401
rect 17040 26435 17092 26444
rect 17040 26401 17049 26435
rect 17049 26401 17083 26435
rect 17083 26401 17092 26435
rect 17040 26392 17092 26401
rect 10968 26324 11020 26376
rect 15752 26324 15804 26376
rect 16672 26324 16724 26376
rect 19708 26367 19760 26376
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 20720 26392 20772 26444
rect 24676 26392 24728 26444
rect 20904 26367 20956 26376
rect 20904 26333 20913 26367
rect 20913 26333 20947 26367
rect 20947 26333 20956 26367
rect 20904 26324 20956 26333
rect 25320 26367 25372 26376
rect 25320 26333 25329 26367
rect 25329 26333 25363 26367
rect 25363 26333 25372 26367
rect 25320 26324 25372 26333
rect 25964 26392 26016 26444
rect 27528 26392 27580 26444
rect 29000 26392 29052 26444
rect 30288 26392 30340 26444
rect 33508 26435 33560 26444
rect 33508 26401 33517 26435
rect 33517 26401 33551 26435
rect 33551 26401 33560 26435
rect 33508 26392 33560 26401
rect 33876 26392 33928 26444
rect 34704 26392 34756 26444
rect 36820 26392 36872 26444
rect 26056 26324 26108 26376
rect 26240 26367 26292 26376
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 26332 26324 26384 26376
rect 26700 26324 26752 26376
rect 26976 26367 27028 26376
rect 26976 26333 26988 26367
rect 26988 26333 27022 26367
rect 27022 26333 27028 26367
rect 26976 26324 27028 26333
rect 12532 26256 12584 26308
rect 17224 26299 17276 26308
rect 17224 26265 17233 26299
rect 17233 26265 17267 26299
rect 17267 26265 17276 26299
rect 17224 26256 17276 26265
rect 24400 26256 24452 26308
rect 15108 26188 15160 26240
rect 25872 26256 25924 26308
rect 24860 26188 24912 26240
rect 26240 26188 26292 26240
rect 27252 26188 27304 26240
rect 28816 26256 28868 26308
rect 29460 26367 29512 26376
rect 29460 26333 29469 26367
rect 29469 26333 29503 26367
rect 29503 26333 29512 26367
rect 29460 26324 29512 26333
rect 31300 26367 31352 26376
rect 31300 26333 31309 26367
rect 31309 26333 31343 26367
rect 31343 26333 31352 26367
rect 31300 26324 31352 26333
rect 32312 26324 32364 26376
rect 32772 26367 32824 26376
rect 32772 26333 32781 26367
rect 32781 26333 32815 26367
rect 32815 26333 32824 26367
rect 32772 26324 32824 26333
rect 34244 26367 34296 26376
rect 34244 26333 34253 26367
rect 34253 26333 34287 26367
rect 34287 26333 34296 26367
rect 34244 26324 34296 26333
rect 34796 26324 34848 26376
rect 31208 26188 31260 26240
rect 31760 26188 31812 26240
rect 33140 26231 33192 26240
rect 33140 26197 33149 26231
rect 33149 26197 33183 26231
rect 33183 26197 33192 26231
rect 33140 26188 33192 26197
rect 33692 26231 33744 26240
rect 33692 26197 33701 26231
rect 33701 26197 33735 26231
rect 33735 26197 33744 26231
rect 33692 26188 33744 26197
rect 35624 26188 35676 26240
rect 36912 26299 36964 26308
rect 36912 26265 36921 26299
rect 36921 26265 36955 26299
rect 36955 26265 36964 26299
rect 36912 26256 36964 26265
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 6920 25984 6972 26036
rect 8300 26027 8352 26036
rect 8300 25993 8309 26027
rect 8309 25993 8343 26027
rect 8343 25993 8352 26027
rect 8300 25984 8352 25993
rect 11796 26027 11848 26036
rect 11796 25993 11805 26027
rect 11805 25993 11839 26027
rect 11839 25993 11848 26027
rect 11796 25984 11848 25993
rect 12440 26027 12492 26036
rect 12440 25993 12449 26027
rect 12449 25993 12483 26027
rect 12483 25993 12492 26027
rect 17040 26027 17092 26036
rect 12440 25984 12492 25993
rect 17040 25993 17049 26027
rect 17049 25993 17083 26027
rect 17083 25993 17092 26027
rect 17040 25984 17092 25993
rect 20812 25984 20864 26036
rect 22652 26027 22704 26036
rect 22652 25993 22661 26027
rect 22661 25993 22695 26027
rect 22695 25993 22704 26027
rect 22652 25984 22704 25993
rect 25320 25984 25372 26036
rect 27620 25984 27672 26036
rect 29000 25984 29052 26036
rect 30380 25984 30432 26036
rect 31208 26027 31260 26036
rect 18972 25916 19024 25968
rect 25964 25959 26016 25968
rect 25964 25925 25973 25959
rect 25973 25925 26007 25959
rect 26007 25925 26016 25959
rect 25964 25916 26016 25925
rect 31208 25993 31217 26027
rect 31217 25993 31251 26027
rect 31251 25993 31260 26027
rect 31208 25984 31260 25993
rect 31576 26027 31628 26036
rect 31576 25993 31585 26027
rect 31585 25993 31619 26027
rect 31619 25993 31628 26027
rect 31576 25984 31628 25993
rect 32312 26027 32364 26036
rect 32312 25993 32321 26027
rect 32321 25993 32355 26027
rect 32355 25993 32364 26027
rect 32312 25984 32364 25993
rect 32680 26027 32732 26036
rect 32680 25993 32689 26027
rect 32689 25993 32723 26027
rect 32723 25993 32732 26027
rect 34704 26027 34756 26036
rect 32680 25984 32732 25993
rect 34704 25993 34713 26027
rect 34713 25993 34747 26027
rect 34747 25993 34756 26027
rect 34704 25984 34756 25993
rect 35532 25984 35584 26036
rect 33140 25916 33192 25968
rect 7012 25780 7064 25832
rect 9680 25823 9732 25832
rect 9680 25789 9689 25823
rect 9689 25789 9723 25823
rect 9723 25789 9732 25823
rect 9680 25780 9732 25789
rect 12900 25848 12952 25900
rect 10416 25823 10468 25832
rect 10416 25789 10450 25823
rect 10450 25789 10468 25823
rect 7104 25712 7156 25764
rect 10416 25780 10468 25789
rect 15292 25823 15344 25832
rect 15292 25789 15301 25823
rect 15301 25789 15335 25823
rect 15335 25789 15344 25823
rect 15292 25780 15344 25789
rect 21088 25848 21140 25900
rect 22008 25848 22060 25900
rect 24308 25848 24360 25900
rect 24860 25891 24912 25900
rect 24860 25857 24869 25891
rect 24869 25857 24903 25891
rect 24903 25857 24912 25891
rect 24860 25848 24912 25857
rect 26240 25848 26292 25900
rect 27068 25848 27120 25900
rect 27528 25848 27580 25900
rect 29460 25891 29512 25900
rect 29460 25857 29469 25891
rect 29469 25857 29503 25891
rect 29503 25857 29512 25891
rect 29460 25848 29512 25857
rect 34244 25848 34296 25900
rect 15936 25780 15988 25832
rect 18328 25780 18380 25832
rect 10692 25712 10744 25764
rect 11520 25687 11572 25696
rect 11520 25653 11529 25687
rect 11529 25653 11563 25687
rect 11563 25653 11572 25687
rect 11520 25644 11572 25653
rect 12532 25644 12584 25696
rect 15844 25644 15896 25696
rect 18788 25644 18840 25696
rect 20628 25780 20680 25832
rect 21548 25823 21600 25832
rect 19708 25712 19760 25764
rect 21548 25789 21557 25823
rect 21557 25789 21591 25823
rect 21591 25789 21600 25823
rect 21548 25780 21600 25789
rect 23664 25780 23716 25832
rect 27252 25823 27304 25832
rect 27252 25789 27261 25823
rect 27261 25789 27295 25823
rect 27295 25789 27304 25823
rect 27252 25780 27304 25789
rect 31576 25780 31628 25832
rect 33140 25823 33192 25832
rect 33140 25789 33149 25823
rect 33149 25789 33183 25823
rect 33183 25789 33192 25823
rect 33140 25780 33192 25789
rect 35624 25823 35676 25832
rect 35624 25789 35633 25823
rect 35633 25789 35667 25823
rect 35667 25789 35676 25823
rect 35624 25780 35676 25789
rect 26976 25712 27028 25764
rect 30748 25712 30800 25764
rect 35532 25712 35584 25764
rect 19248 25644 19300 25696
rect 20812 25644 20864 25696
rect 26608 25687 26660 25696
rect 26608 25653 26617 25687
rect 26617 25653 26651 25687
rect 26651 25653 26660 25687
rect 26608 25644 26660 25653
rect 32772 25687 32824 25696
rect 32772 25653 32781 25687
rect 32781 25653 32815 25687
rect 32815 25653 32824 25687
rect 32772 25644 32824 25653
rect 32864 25644 32916 25696
rect 33784 25687 33836 25696
rect 33784 25653 33793 25687
rect 33793 25653 33827 25687
rect 33827 25653 33836 25687
rect 33784 25644 33836 25653
rect 33876 25644 33928 25696
rect 34796 25644 34848 25696
rect 36820 25687 36872 25696
rect 36820 25653 36829 25687
rect 36829 25653 36863 25687
rect 36863 25653 36872 25687
rect 36820 25644 36872 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 10692 25440 10744 25492
rect 10968 25440 11020 25492
rect 12532 25483 12584 25492
rect 12532 25449 12541 25483
rect 12541 25449 12575 25483
rect 12575 25449 12584 25483
rect 12532 25440 12584 25449
rect 19156 25440 19208 25492
rect 20720 25483 20772 25492
rect 20720 25449 20729 25483
rect 20729 25449 20763 25483
rect 20763 25449 20772 25483
rect 20720 25440 20772 25449
rect 21088 25483 21140 25492
rect 21088 25449 21097 25483
rect 21097 25449 21131 25483
rect 21131 25449 21140 25483
rect 21088 25440 21140 25449
rect 21548 25483 21600 25492
rect 21548 25449 21557 25483
rect 21557 25449 21591 25483
rect 21591 25449 21600 25483
rect 21548 25440 21600 25449
rect 23664 25483 23716 25492
rect 23664 25449 23673 25483
rect 23673 25449 23707 25483
rect 23707 25449 23716 25483
rect 23664 25440 23716 25449
rect 25320 25440 25372 25492
rect 26240 25483 26292 25492
rect 26240 25449 26249 25483
rect 26249 25449 26283 25483
rect 26283 25449 26292 25483
rect 26240 25440 26292 25449
rect 27252 25440 27304 25492
rect 27528 25483 27580 25492
rect 27528 25449 27537 25483
rect 27537 25449 27571 25483
rect 27571 25449 27580 25483
rect 27528 25440 27580 25449
rect 29460 25440 29512 25492
rect 30748 25483 30800 25492
rect 30748 25449 30757 25483
rect 30757 25449 30791 25483
rect 30791 25449 30800 25483
rect 30748 25440 30800 25449
rect 33784 25440 33836 25492
rect 34244 25440 34296 25492
rect 14096 25372 14148 25424
rect 20628 25372 20680 25424
rect 20996 25372 21048 25424
rect 24216 25372 24268 25424
rect 24676 25372 24728 25424
rect 26976 25372 27028 25424
rect 34704 25372 34756 25424
rect 35624 25372 35676 25424
rect 7012 25304 7064 25356
rect 7196 25304 7248 25356
rect 10048 25304 10100 25356
rect 11520 25304 11572 25356
rect 10692 25279 10744 25288
rect 10692 25245 10701 25279
rect 10701 25245 10735 25279
rect 10735 25245 10744 25279
rect 10692 25236 10744 25245
rect 13728 25236 13780 25288
rect 15108 25304 15160 25356
rect 14464 25236 14516 25288
rect 7104 25100 7156 25152
rect 8208 25100 8260 25152
rect 10140 25143 10192 25152
rect 10140 25109 10149 25143
rect 10149 25109 10183 25143
rect 10183 25109 10192 25143
rect 10140 25100 10192 25109
rect 11060 25100 11112 25152
rect 12532 25100 12584 25152
rect 12900 25143 12952 25152
rect 12900 25109 12909 25143
rect 12909 25109 12943 25143
rect 12943 25109 12952 25143
rect 12900 25100 12952 25109
rect 13636 25143 13688 25152
rect 13636 25109 13645 25143
rect 13645 25109 13679 25143
rect 13679 25109 13688 25143
rect 13636 25100 13688 25109
rect 14740 25143 14792 25152
rect 14740 25109 14749 25143
rect 14749 25109 14783 25143
rect 14783 25109 14792 25143
rect 14740 25100 14792 25109
rect 15016 25143 15068 25152
rect 15016 25109 15025 25143
rect 15025 25109 15059 25143
rect 15059 25109 15068 25143
rect 15844 25304 15896 25356
rect 18144 25347 18196 25356
rect 18144 25313 18153 25347
rect 18153 25313 18187 25347
rect 18187 25313 18196 25347
rect 18144 25304 18196 25313
rect 19616 25347 19668 25356
rect 19616 25313 19625 25347
rect 19625 25313 19659 25347
rect 19659 25313 19668 25347
rect 19616 25304 19668 25313
rect 20260 25304 20312 25356
rect 20904 25347 20956 25356
rect 20904 25313 20913 25347
rect 20913 25313 20947 25347
rect 20947 25313 20956 25347
rect 20904 25304 20956 25313
rect 28172 25347 28224 25356
rect 28172 25313 28181 25347
rect 28181 25313 28215 25347
rect 28215 25313 28224 25347
rect 28172 25304 28224 25313
rect 28816 25304 28868 25356
rect 29000 25304 29052 25356
rect 31944 25304 31996 25356
rect 32128 25304 32180 25356
rect 33692 25304 33744 25356
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 15292 25236 15344 25245
rect 16672 25236 16724 25288
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 23480 25236 23532 25288
rect 23848 25236 23900 25288
rect 28448 25279 28500 25288
rect 28448 25245 28457 25279
rect 28457 25245 28491 25279
rect 28491 25245 28500 25279
rect 28448 25236 28500 25245
rect 29368 25279 29420 25288
rect 29368 25245 29377 25279
rect 29377 25245 29411 25279
rect 29411 25245 29420 25279
rect 29368 25236 29420 25245
rect 32772 25236 32824 25288
rect 34060 25279 34112 25288
rect 34060 25245 34069 25279
rect 34069 25245 34103 25279
rect 34103 25245 34112 25279
rect 34060 25236 34112 25245
rect 15016 25100 15068 25109
rect 15936 25100 15988 25152
rect 16580 25100 16632 25152
rect 17408 25143 17460 25152
rect 17408 25109 17417 25143
rect 17417 25109 17451 25143
rect 17451 25109 17460 25143
rect 17408 25100 17460 25109
rect 18604 25100 18656 25152
rect 18696 25143 18748 25152
rect 18696 25109 18705 25143
rect 18705 25109 18739 25143
rect 18739 25109 18748 25143
rect 18696 25100 18748 25109
rect 24860 25100 24912 25152
rect 27804 25143 27856 25152
rect 27804 25109 27813 25143
rect 27813 25109 27847 25143
rect 27847 25109 27856 25143
rect 27804 25100 27856 25109
rect 32864 25143 32916 25152
rect 32864 25109 32873 25143
rect 32873 25109 32907 25143
rect 32907 25109 32916 25143
rect 32864 25100 32916 25109
rect 33416 25143 33468 25152
rect 33416 25109 33425 25143
rect 33425 25109 33459 25143
rect 33459 25109 33468 25143
rect 33416 25100 33468 25109
rect 34796 25143 34848 25152
rect 34796 25109 34805 25143
rect 34805 25109 34839 25143
rect 34839 25109 34848 25143
rect 34796 25100 34848 25109
rect 36360 25143 36412 25152
rect 36360 25109 36369 25143
rect 36369 25109 36403 25143
rect 36403 25109 36412 25143
rect 36360 25100 36412 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 7012 24896 7064 24948
rect 9680 24939 9732 24948
rect 9680 24905 9689 24939
rect 9689 24905 9723 24939
rect 9723 24905 9732 24939
rect 9680 24896 9732 24905
rect 10048 24939 10100 24948
rect 10048 24905 10057 24939
rect 10057 24905 10091 24939
rect 10091 24905 10100 24939
rect 10048 24896 10100 24905
rect 12440 24939 12492 24948
rect 12440 24905 12449 24939
rect 12449 24905 12483 24939
rect 12483 24905 12492 24939
rect 12440 24896 12492 24905
rect 15016 24896 15068 24948
rect 18328 24939 18380 24948
rect 18328 24905 18337 24939
rect 18337 24905 18371 24939
rect 18371 24905 18380 24939
rect 18328 24896 18380 24905
rect 19800 24939 19852 24948
rect 19800 24905 19809 24939
rect 19809 24905 19843 24939
rect 19843 24905 19852 24939
rect 19800 24896 19852 24905
rect 20812 24896 20864 24948
rect 23848 24896 23900 24948
rect 24216 24939 24268 24948
rect 24216 24905 24225 24939
rect 24225 24905 24259 24939
rect 24259 24905 24268 24939
rect 24216 24896 24268 24905
rect 28448 24896 28500 24948
rect 29000 24896 29052 24948
rect 12900 24828 12952 24880
rect 11888 24803 11940 24812
rect 11888 24769 11897 24803
rect 11897 24769 11931 24803
rect 11931 24769 11940 24803
rect 11888 24760 11940 24769
rect 15936 24828 15988 24880
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 7380 24735 7432 24744
rect 7380 24701 7389 24735
rect 7389 24701 7423 24735
rect 7423 24701 7432 24735
rect 7380 24692 7432 24701
rect 10140 24735 10192 24744
rect 10140 24701 10149 24735
rect 10149 24701 10183 24735
rect 10183 24701 10192 24735
rect 10140 24692 10192 24701
rect 14740 24692 14792 24744
rect 17500 24760 17552 24812
rect 17868 24760 17920 24812
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 20904 24828 20956 24880
rect 20996 24760 21048 24812
rect 23940 24803 23992 24812
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 17408 24692 17460 24744
rect 18604 24692 18656 24744
rect 19892 24735 19944 24744
rect 19892 24701 19901 24735
rect 19901 24701 19935 24735
rect 19935 24701 19944 24735
rect 19892 24692 19944 24701
rect 19984 24692 20036 24744
rect 29000 24760 29052 24812
rect 32128 24896 32180 24948
rect 32772 24896 32824 24948
rect 33140 24939 33192 24948
rect 33140 24905 33149 24939
rect 33149 24905 33183 24939
rect 33183 24905 33192 24939
rect 33140 24896 33192 24905
rect 33876 24939 33928 24948
rect 33876 24905 33885 24939
rect 33885 24905 33919 24939
rect 33919 24905 33928 24939
rect 33876 24896 33928 24905
rect 34704 24939 34756 24948
rect 34704 24905 34713 24939
rect 34713 24905 34747 24939
rect 34747 24905 34756 24939
rect 34704 24896 34756 24905
rect 36360 24939 36412 24948
rect 36360 24905 36369 24939
rect 36369 24905 36403 24939
rect 36403 24905 36412 24939
rect 36360 24896 36412 24905
rect 36636 24939 36688 24948
rect 36636 24905 36645 24939
rect 36645 24905 36679 24939
rect 36679 24905 36688 24939
rect 36636 24896 36688 24905
rect 31300 24828 31352 24880
rect 31760 24828 31812 24880
rect 32772 24760 32824 24812
rect 24768 24735 24820 24744
rect 24768 24701 24791 24735
rect 24791 24701 24820 24735
rect 7656 24667 7708 24676
rect 7656 24633 7690 24667
rect 7690 24633 7708 24667
rect 7656 24624 7708 24633
rect 10232 24624 10284 24676
rect 15108 24667 15160 24676
rect 15108 24633 15142 24667
rect 15142 24633 15160 24667
rect 15108 24624 15160 24633
rect 18144 24624 18196 24676
rect 19616 24624 19668 24676
rect 24768 24692 24820 24701
rect 29368 24692 29420 24744
rect 34428 24692 34480 24744
rect 35900 24760 35952 24812
rect 37188 24760 37240 24812
rect 24584 24624 24636 24676
rect 28816 24624 28868 24676
rect 30564 24624 30616 24676
rect 33876 24624 33928 24676
rect 8760 24599 8812 24608
rect 8760 24565 8769 24599
rect 8769 24565 8803 24599
rect 8803 24565 8812 24599
rect 8760 24556 8812 24565
rect 11520 24599 11572 24608
rect 11520 24565 11529 24599
rect 11529 24565 11563 24599
rect 11563 24565 11572 24599
rect 11520 24556 11572 24565
rect 12164 24599 12216 24608
rect 12164 24565 12173 24599
rect 12173 24565 12207 24599
rect 12207 24565 12216 24599
rect 12164 24556 12216 24565
rect 12532 24556 12584 24608
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 15660 24556 15712 24608
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 18696 24599 18748 24608
rect 18696 24565 18705 24599
rect 18705 24565 18739 24599
rect 18739 24565 18748 24599
rect 18696 24556 18748 24565
rect 25872 24599 25924 24608
rect 25872 24565 25881 24599
rect 25881 24565 25915 24599
rect 25915 24565 25924 24599
rect 25872 24556 25924 24565
rect 28172 24556 28224 24608
rect 31852 24599 31904 24608
rect 31852 24565 31861 24599
rect 31861 24565 31895 24599
rect 31895 24565 31904 24599
rect 31852 24556 31904 24565
rect 34796 24556 34848 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 7196 24395 7248 24404
rect 7196 24361 7205 24395
rect 7205 24361 7239 24395
rect 7239 24361 7248 24395
rect 7196 24352 7248 24361
rect 7840 24395 7892 24404
rect 7840 24361 7849 24395
rect 7849 24361 7883 24395
rect 7883 24361 7892 24395
rect 7840 24352 7892 24361
rect 10232 24395 10284 24404
rect 10232 24361 10241 24395
rect 10241 24361 10275 24395
rect 10275 24361 10284 24395
rect 10232 24352 10284 24361
rect 12164 24352 12216 24404
rect 14096 24352 14148 24404
rect 15660 24395 15712 24404
rect 15660 24361 15669 24395
rect 15669 24361 15703 24395
rect 15703 24361 15712 24395
rect 15660 24352 15712 24361
rect 7932 24284 7984 24336
rect 8760 24284 8812 24336
rect 10968 24284 11020 24336
rect 11520 24284 11572 24336
rect 12532 24327 12584 24336
rect 12532 24293 12541 24327
rect 12541 24293 12575 24327
rect 12575 24293 12584 24327
rect 12532 24284 12584 24293
rect 15108 24284 15160 24336
rect 16488 24352 16540 24404
rect 17776 24352 17828 24404
rect 18972 24352 19024 24404
rect 19984 24395 20036 24404
rect 19984 24361 19993 24395
rect 19993 24361 20027 24395
rect 20027 24361 20036 24395
rect 19984 24352 20036 24361
rect 20260 24395 20312 24404
rect 20260 24361 20269 24395
rect 20269 24361 20303 24395
rect 20303 24361 20312 24395
rect 20260 24352 20312 24361
rect 24308 24395 24360 24404
rect 24308 24361 24317 24395
rect 24317 24361 24351 24395
rect 24351 24361 24360 24395
rect 24308 24352 24360 24361
rect 27528 24352 27580 24404
rect 29368 24352 29420 24404
rect 30564 24352 30616 24404
rect 30748 24352 30800 24404
rect 31852 24352 31904 24404
rect 31944 24395 31996 24404
rect 31944 24361 31953 24395
rect 31953 24361 31987 24395
rect 31987 24361 31996 24395
rect 31944 24352 31996 24361
rect 32864 24352 32916 24404
rect 33048 24352 33100 24404
rect 33692 24352 33744 24404
rect 34060 24352 34112 24404
rect 36912 24352 36964 24404
rect 19892 24284 19944 24336
rect 8208 24259 8260 24268
rect 8208 24225 8217 24259
rect 8217 24225 8251 24259
rect 8251 24225 8260 24259
rect 8208 24216 8260 24225
rect 10692 24216 10744 24268
rect 13268 24216 13320 24268
rect 13636 24216 13688 24268
rect 17776 24216 17828 24268
rect 18880 24259 18932 24268
rect 18880 24225 18914 24259
rect 18914 24225 18932 24259
rect 18880 24216 18932 24225
rect 20720 24284 20772 24336
rect 23480 24284 23532 24336
rect 35900 24284 35952 24336
rect 20996 24216 21048 24268
rect 24032 24216 24084 24268
rect 27436 24259 27488 24268
rect 27436 24225 27445 24259
rect 27445 24225 27479 24259
rect 27479 24225 27488 24259
rect 27436 24216 27488 24225
rect 29552 24259 29604 24268
rect 29552 24225 29586 24259
rect 29586 24225 29604 24259
rect 29552 24216 29604 24225
rect 32036 24216 32088 24268
rect 34888 24216 34940 24268
rect 35532 24216 35584 24268
rect 36452 24259 36504 24268
rect 36452 24225 36461 24259
rect 36461 24225 36495 24259
rect 36495 24225 36504 24259
rect 36452 24216 36504 24225
rect 8484 24191 8536 24200
rect 8484 24157 8493 24191
rect 8493 24157 8527 24191
rect 8527 24157 8536 24191
rect 8484 24148 8536 24157
rect 10140 24148 10192 24200
rect 10416 24148 10468 24200
rect 15200 24148 15252 24200
rect 15752 24148 15804 24200
rect 17316 24191 17368 24200
rect 7380 24080 7432 24132
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 21364 24191 21416 24200
rect 21364 24157 21373 24191
rect 21373 24157 21407 24191
rect 21407 24157 21416 24191
rect 21364 24148 21416 24157
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 24216 24148 24268 24200
rect 25872 24148 25924 24200
rect 29000 24148 29052 24200
rect 16948 24080 17000 24132
rect 14464 24012 14516 24064
rect 25136 24012 25188 24064
rect 35624 24055 35676 24064
rect 35624 24021 35633 24055
rect 35633 24021 35667 24055
rect 35667 24021 35676 24055
rect 35624 24012 35676 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 7932 23851 7984 23860
rect 7932 23817 7941 23851
rect 7941 23817 7975 23851
rect 7975 23817 7984 23851
rect 7932 23808 7984 23817
rect 8208 23851 8260 23860
rect 8208 23817 8217 23851
rect 8217 23817 8251 23851
rect 8251 23817 8260 23851
rect 8208 23808 8260 23817
rect 8484 23808 8536 23860
rect 10692 23851 10744 23860
rect 10692 23817 10701 23851
rect 10701 23817 10735 23851
rect 10735 23817 10744 23851
rect 10692 23808 10744 23817
rect 10784 23808 10836 23860
rect 13268 23851 13320 23860
rect 13268 23817 13277 23851
rect 13277 23817 13311 23851
rect 13311 23817 13320 23851
rect 13268 23808 13320 23817
rect 15108 23808 15160 23860
rect 15660 23808 15712 23860
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 17316 23808 17368 23860
rect 17776 23851 17828 23860
rect 17776 23817 17785 23851
rect 17785 23817 17819 23851
rect 17819 23817 17828 23851
rect 17776 23808 17828 23817
rect 19340 23808 19392 23860
rect 19984 23851 20036 23860
rect 19984 23817 19993 23851
rect 19993 23817 20027 23851
rect 20027 23817 20036 23851
rect 19984 23808 20036 23817
rect 20720 23851 20772 23860
rect 20720 23817 20729 23851
rect 20729 23817 20763 23851
rect 20763 23817 20772 23851
rect 20720 23808 20772 23817
rect 22008 23808 22060 23860
rect 23480 23808 23532 23860
rect 24584 23808 24636 23860
rect 27436 23808 27488 23860
rect 28080 23808 28132 23860
rect 28908 23851 28960 23860
rect 10416 23740 10468 23792
rect 11796 23740 11848 23792
rect 18788 23740 18840 23792
rect 21364 23740 21416 23792
rect 11060 23604 11112 23656
rect 12348 23604 12400 23656
rect 15660 23604 15712 23656
rect 16488 23604 16540 23656
rect 17408 23672 17460 23724
rect 24032 23672 24084 23724
rect 27528 23740 27580 23792
rect 17500 23604 17552 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 19432 23647 19484 23656
rect 19432 23613 19441 23647
rect 19441 23613 19475 23647
rect 19475 23613 19484 23647
rect 19432 23604 19484 23613
rect 25136 23647 25188 23656
rect 25136 23613 25145 23647
rect 25145 23613 25179 23647
rect 25179 23613 25188 23647
rect 25136 23604 25188 23613
rect 14740 23536 14792 23588
rect 16948 23536 17000 23588
rect 19984 23536 20036 23588
rect 21548 23536 21600 23588
rect 25044 23536 25096 23588
rect 14372 23468 14424 23520
rect 16580 23468 16632 23520
rect 24860 23468 24912 23520
rect 28908 23817 28917 23851
rect 28917 23817 28951 23851
rect 28951 23817 28960 23851
rect 28908 23808 28960 23817
rect 29552 23851 29604 23860
rect 29552 23817 29561 23851
rect 29561 23817 29595 23851
rect 29595 23817 29604 23851
rect 31300 23851 31352 23860
rect 29552 23808 29604 23817
rect 28816 23740 28868 23792
rect 31300 23817 31309 23851
rect 31309 23817 31343 23851
rect 31343 23817 31352 23851
rect 31300 23808 31352 23817
rect 32036 23808 32088 23860
rect 32772 23851 32824 23860
rect 32772 23817 32781 23851
rect 32781 23817 32815 23851
rect 32815 23817 32824 23851
rect 32772 23808 32824 23817
rect 33140 23851 33192 23860
rect 33140 23817 33149 23851
rect 33149 23817 33183 23851
rect 33183 23817 33192 23851
rect 33140 23808 33192 23817
rect 33416 23808 33468 23860
rect 33876 23851 33928 23860
rect 30288 23672 30340 23724
rect 33140 23604 33192 23656
rect 33876 23817 33885 23851
rect 33885 23817 33919 23851
rect 33919 23817 33928 23851
rect 33876 23808 33928 23817
rect 35900 23851 35952 23860
rect 35900 23817 35909 23851
rect 35909 23817 35943 23851
rect 35943 23817 35952 23851
rect 35900 23808 35952 23817
rect 36452 23851 36504 23860
rect 36452 23817 36461 23851
rect 36461 23817 36495 23851
rect 36495 23817 36504 23851
rect 36452 23808 36504 23817
rect 34428 23672 34480 23724
rect 35624 23672 35676 23724
rect 34520 23604 34572 23656
rect 34796 23604 34848 23656
rect 26148 23536 26200 23588
rect 30564 23536 30616 23588
rect 35992 23536 36044 23588
rect 25596 23511 25648 23520
rect 25596 23477 25605 23511
rect 25605 23477 25639 23511
rect 25639 23477 25648 23511
rect 25596 23468 25648 23477
rect 28908 23468 28960 23520
rect 34244 23468 34296 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 10416 23307 10468 23316
rect 10416 23273 10425 23307
rect 10425 23273 10459 23307
rect 10459 23273 10468 23307
rect 10416 23264 10468 23273
rect 12440 23264 12492 23316
rect 15108 23307 15160 23316
rect 15108 23273 15117 23307
rect 15117 23273 15151 23307
rect 15151 23273 15160 23307
rect 15108 23264 15160 23273
rect 15292 23307 15344 23316
rect 15292 23273 15301 23307
rect 15301 23273 15335 23307
rect 15335 23273 15344 23307
rect 15292 23264 15344 23273
rect 18880 23264 18932 23316
rect 21456 23264 21508 23316
rect 28080 23307 28132 23316
rect 28080 23273 28089 23307
rect 28089 23273 28123 23307
rect 28123 23273 28132 23307
rect 28080 23264 28132 23273
rect 30288 23307 30340 23316
rect 30288 23273 30297 23307
rect 30297 23273 30331 23307
rect 30331 23273 30340 23307
rect 30288 23264 30340 23273
rect 30564 23307 30616 23316
rect 30564 23273 30573 23307
rect 30573 23273 30607 23307
rect 30607 23273 30616 23307
rect 30564 23264 30616 23273
rect 34520 23264 34572 23316
rect 35532 23264 35584 23316
rect 35992 23264 36044 23316
rect 19432 23239 19484 23248
rect 19432 23205 19466 23239
rect 19466 23205 19484 23239
rect 19432 23196 19484 23205
rect 25136 23196 25188 23248
rect 33600 23196 33652 23248
rect 34244 23196 34296 23248
rect 34428 23239 34480 23248
rect 34428 23205 34462 23239
rect 34462 23205 34480 23239
rect 34428 23196 34480 23205
rect 10508 23128 10560 23180
rect 11060 23128 11112 23180
rect 12716 23171 12768 23180
rect 12716 23137 12725 23171
rect 12725 23137 12759 23171
rect 12759 23137 12768 23171
rect 12716 23128 12768 23137
rect 13268 23171 13320 23180
rect 13268 23137 13302 23171
rect 13302 23137 13320 23171
rect 13268 23128 13320 23137
rect 15660 23171 15712 23180
rect 15660 23137 15669 23171
rect 15669 23137 15703 23171
rect 15703 23137 15712 23171
rect 15660 23128 15712 23137
rect 17592 23128 17644 23180
rect 18604 23128 18656 23180
rect 24676 23171 24728 23180
rect 24676 23137 24685 23171
rect 24685 23137 24719 23171
rect 24719 23137 24728 23171
rect 24676 23128 24728 23137
rect 27804 23128 27856 23180
rect 29184 23171 29236 23180
rect 29184 23137 29218 23171
rect 29218 23137 29236 23171
rect 29184 23128 29236 23137
rect 33048 23171 33100 23180
rect 33048 23137 33057 23171
rect 33057 23137 33091 23171
rect 33091 23137 33100 23171
rect 33048 23128 33100 23137
rect 15384 23060 15436 23112
rect 17316 23103 17368 23112
rect 14464 22992 14516 23044
rect 15016 22992 15068 23044
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 28908 23103 28960 23112
rect 16028 22992 16080 23044
rect 17224 22992 17276 23044
rect 28908 23069 28917 23103
rect 28917 23069 28951 23103
rect 28951 23069 28960 23103
rect 28908 23060 28960 23069
rect 31208 23060 31260 23112
rect 34060 23060 34112 23112
rect 13636 22924 13688 22976
rect 14280 22924 14332 22976
rect 16396 22967 16448 22976
rect 16396 22933 16405 22967
rect 16405 22933 16439 22967
rect 16439 22933 16448 22967
rect 16396 22924 16448 22933
rect 16672 22924 16724 22976
rect 18420 22967 18472 22976
rect 18420 22933 18429 22967
rect 18429 22933 18463 22967
rect 18463 22933 18472 22967
rect 18420 22924 18472 22933
rect 21548 22967 21600 22976
rect 21548 22933 21557 22967
rect 21557 22933 21591 22967
rect 21591 22933 21600 22967
rect 21548 22924 21600 22933
rect 22100 22967 22152 22976
rect 22100 22933 22109 22967
rect 22109 22933 22143 22967
rect 22143 22933 22152 22967
rect 22100 22924 22152 22933
rect 24216 22924 24268 22976
rect 25872 22924 25924 22976
rect 33232 22967 33284 22976
rect 33232 22933 33241 22967
rect 33241 22933 33275 22967
rect 33275 22933 33284 22967
rect 33232 22924 33284 22933
rect 35532 22967 35584 22976
rect 35532 22933 35541 22967
rect 35541 22933 35575 22967
rect 35575 22933 35584 22967
rect 35532 22924 35584 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 10508 22763 10560 22772
rect 10508 22729 10517 22763
rect 10517 22729 10551 22763
rect 10551 22729 10560 22763
rect 10508 22720 10560 22729
rect 12624 22720 12676 22772
rect 12992 22763 13044 22772
rect 12992 22729 13001 22763
rect 13001 22729 13035 22763
rect 13035 22729 13044 22763
rect 12992 22720 13044 22729
rect 15384 22763 15436 22772
rect 15384 22729 15393 22763
rect 15393 22729 15427 22763
rect 15427 22729 15436 22763
rect 15384 22720 15436 22729
rect 15660 22720 15712 22772
rect 17316 22763 17368 22772
rect 17316 22729 17325 22763
rect 17325 22729 17359 22763
rect 17359 22729 17368 22763
rect 17316 22720 17368 22729
rect 17592 22763 17644 22772
rect 17592 22729 17601 22763
rect 17601 22729 17635 22763
rect 17635 22729 17644 22763
rect 17592 22720 17644 22729
rect 19432 22720 19484 22772
rect 20996 22720 21048 22772
rect 25136 22720 25188 22772
rect 25688 22763 25740 22772
rect 25688 22729 25697 22763
rect 25697 22729 25731 22763
rect 25731 22729 25740 22763
rect 25688 22720 25740 22729
rect 30748 22763 30800 22772
rect 30748 22729 30757 22763
rect 30757 22729 30791 22763
rect 30791 22729 30800 22763
rect 31208 22763 31260 22772
rect 30748 22720 30800 22729
rect 31208 22729 31217 22763
rect 31217 22729 31251 22763
rect 31251 22729 31260 22763
rect 31208 22720 31260 22729
rect 13268 22584 13320 22636
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 14648 22584 14700 22636
rect 15108 22584 15160 22636
rect 16028 22627 16080 22636
rect 16028 22593 16037 22627
rect 16037 22593 16071 22627
rect 16071 22593 16080 22627
rect 16028 22584 16080 22593
rect 23388 22584 23440 22636
rect 30104 22584 30156 22636
rect 15844 22491 15896 22500
rect 15844 22457 15853 22491
rect 15853 22457 15887 22491
rect 15887 22457 15896 22491
rect 15844 22448 15896 22457
rect 13820 22380 13872 22432
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 16304 22380 16356 22432
rect 18052 22380 18104 22432
rect 18420 22516 18472 22568
rect 22100 22516 22152 22568
rect 26884 22559 26936 22568
rect 26884 22525 26893 22559
rect 26893 22525 26927 22559
rect 26927 22525 26936 22559
rect 26884 22516 26936 22525
rect 29184 22516 29236 22568
rect 31944 22720 31996 22772
rect 33048 22720 33100 22772
rect 34428 22720 34480 22772
rect 34244 22516 34296 22568
rect 34888 22559 34940 22568
rect 34888 22525 34897 22559
rect 34897 22525 34931 22559
rect 34931 22525 34940 22559
rect 34888 22516 34940 22525
rect 35532 22516 35584 22568
rect 20352 22423 20404 22432
rect 20352 22389 20361 22423
rect 20361 22389 20395 22423
rect 20395 22389 20404 22423
rect 20352 22380 20404 22389
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 22744 22380 22796 22432
rect 23940 22380 23992 22432
rect 30012 22448 30064 22500
rect 33600 22491 33652 22500
rect 33600 22457 33609 22491
rect 33609 22457 33643 22491
rect 33643 22457 33652 22491
rect 33600 22448 33652 22457
rect 34152 22448 34204 22500
rect 36636 22448 36688 22500
rect 25228 22380 25280 22432
rect 27804 22380 27856 22432
rect 29276 22423 29328 22432
rect 29276 22389 29285 22423
rect 29285 22389 29319 22423
rect 29319 22389 29328 22423
rect 29276 22380 29328 22389
rect 29736 22423 29788 22432
rect 29736 22389 29745 22423
rect 29745 22389 29779 22423
rect 29779 22389 29788 22423
rect 29736 22380 29788 22389
rect 33140 22380 33192 22432
rect 36268 22423 36320 22432
rect 36268 22389 36277 22423
rect 36277 22389 36311 22423
rect 36311 22389 36320 22423
rect 36268 22380 36320 22389
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 12624 22219 12676 22228
rect 12624 22185 12633 22219
rect 12633 22185 12667 22219
rect 12667 22185 12676 22219
rect 12624 22176 12676 22185
rect 14648 22219 14700 22228
rect 14648 22185 14657 22219
rect 14657 22185 14691 22219
rect 14691 22185 14700 22219
rect 14648 22176 14700 22185
rect 15016 22219 15068 22228
rect 15016 22185 15025 22219
rect 15025 22185 15059 22219
rect 15059 22185 15068 22219
rect 15016 22176 15068 22185
rect 15660 22176 15712 22228
rect 17316 22176 17368 22228
rect 17592 22176 17644 22228
rect 18512 22176 18564 22228
rect 19340 22176 19392 22228
rect 20352 22176 20404 22228
rect 25136 22176 25188 22228
rect 11796 22040 11848 22092
rect 12808 22083 12860 22092
rect 12808 22049 12817 22083
rect 12817 22049 12851 22083
rect 12851 22049 12860 22083
rect 12808 22040 12860 22049
rect 12992 22040 13044 22092
rect 13728 22040 13780 22092
rect 14740 22040 14792 22092
rect 22100 22108 22152 22160
rect 27620 22151 27672 22160
rect 15108 21972 15160 22024
rect 15936 22040 15988 22092
rect 14280 21947 14332 21956
rect 14280 21913 14289 21947
rect 14289 21913 14323 21947
rect 14323 21913 14332 21947
rect 14280 21904 14332 21913
rect 14648 21904 14700 21956
rect 17684 22040 17736 22092
rect 20996 22040 21048 22092
rect 27620 22117 27629 22151
rect 27629 22117 27663 22151
rect 27663 22117 27672 22151
rect 27620 22108 27672 22117
rect 29276 22176 29328 22228
rect 33968 22176 34020 22228
rect 34060 22176 34112 22228
rect 34888 22176 34940 22228
rect 23756 22083 23808 22092
rect 23756 22049 23779 22083
rect 23779 22049 23808 22083
rect 23756 22040 23808 22049
rect 26240 22040 26292 22092
rect 26516 22083 26568 22092
rect 26516 22049 26525 22083
rect 26525 22049 26559 22083
rect 26559 22049 26568 22083
rect 26516 22040 26568 22049
rect 17316 22015 17368 22024
rect 17316 21981 17325 22015
rect 17325 21981 17359 22015
rect 17359 21981 17368 22015
rect 17316 21972 17368 21981
rect 18880 22015 18932 22024
rect 18880 21981 18889 22015
rect 18889 21981 18923 22015
rect 18923 21981 18932 22015
rect 18880 21972 18932 21981
rect 12900 21836 12952 21888
rect 16304 21879 16356 21888
rect 16304 21845 16313 21879
rect 16313 21845 16347 21879
rect 16347 21845 16356 21879
rect 16304 21836 16356 21845
rect 21272 21836 21324 21888
rect 21640 21836 21692 21888
rect 23112 21836 23164 21888
rect 28816 21972 28868 22024
rect 29460 22040 29512 22092
rect 29736 22083 29788 22092
rect 29736 22049 29745 22083
rect 29745 22049 29779 22083
rect 29779 22049 29788 22083
rect 29736 22040 29788 22049
rect 33600 22083 33652 22092
rect 33600 22049 33609 22083
rect 33609 22049 33643 22083
rect 33643 22049 33652 22083
rect 33600 22040 33652 22049
rect 29184 22015 29236 22024
rect 29184 21981 29193 22015
rect 29193 21981 29227 22015
rect 29227 21981 29236 22015
rect 29184 21972 29236 21981
rect 32956 21972 33008 22024
rect 33140 21972 33192 22024
rect 34704 22040 34756 22092
rect 36268 22108 36320 22160
rect 34796 22015 34848 22024
rect 34796 21981 34805 22015
rect 34805 21981 34839 22015
rect 34839 21981 34848 22015
rect 34796 21972 34848 21981
rect 24676 21836 24728 21888
rect 25504 21836 25556 21888
rect 26700 21879 26752 21888
rect 26700 21845 26709 21879
rect 26709 21845 26743 21879
rect 26743 21845 26752 21879
rect 26700 21836 26752 21845
rect 28632 21879 28684 21888
rect 28632 21845 28641 21879
rect 28641 21845 28675 21879
rect 28675 21845 28684 21879
rect 28632 21836 28684 21845
rect 30104 21879 30156 21888
rect 30104 21845 30113 21879
rect 30113 21845 30147 21879
rect 30147 21845 30156 21879
rect 30104 21836 30156 21845
rect 31208 21836 31260 21888
rect 33140 21879 33192 21888
rect 33140 21845 33149 21879
rect 33149 21845 33183 21879
rect 33183 21845 33192 21879
rect 33140 21836 33192 21845
rect 35716 21836 35768 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12992 21632 13044 21684
rect 14740 21675 14792 21684
rect 14740 21641 14749 21675
rect 14749 21641 14783 21675
rect 14783 21641 14792 21675
rect 14740 21632 14792 21641
rect 15108 21675 15160 21684
rect 15108 21641 15117 21675
rect 15117 21641 15151 21675
rect 15151 21641 15160 21675
rect 15108 21632 15160 21641
rect 16304 21632 16356 21684
rect 16672 21675 16724 21684
rect 16672 21641 16681 21675
rect 16681 21641 16715 21675
rect 16715 21641 16724 21675
rect 16672 21632 16724 21641
rect 16948 21675 17000 21684
rect 16948 21641 16957 21675
rect 16957 21641 16991 21675
rect 16991 21641 17000 21675
rect 16948 21632 17000 21641
rect 17684 21675 17736 21684
rect 17684 21641 17693 21675
rect 17693 21641 17727 21675
rect 17727 21641 17736 21675
rect 17684 21632 17736 21641
rect 19340 21632 19392 21684
rect 22744 21675 22796 21684
rect 22744 21641 22753 21675
rect 22753 21641 22787 21675
rect 22787 21641 22796 21675
rect 22744 21632 22796 21641
rect 23112 21675 23164 21684
rect 23112 21641 23121 21675
rect 23121 21641 23155 21675
rect 23155 21641 23164 21675
rect 23112 21632 23164 21641
rect 23756 21632 23808 21684
rect 24768 21632 24820 21684
rect 26516 21632 26568 21684
rect 28448 21675 28500 21684
rect 28448 21641 28457 21675
rect 28457 21641 28491 21675
rect 28491 21641 28500 21675
rect 28448 21632 28500 21641
rect 28816 21675 28868 21684
rect 28816 21641 28825 21675
rect 28825 21641 28859 21675
rect 28859 21641 28868 21675
rect 28816 21632 28868 21641
rect 29184 21632 29236 21684
rect 33232 21632 33284 21684
rect 34704 21675 34756 21684
rect 34704 21641 34713 21675
rect 34713 21641 34747 21675
rect 34747 21641 34756 21675
rect 34704 21632 34756 21641
rect 36636 21675 36688 21684
rect 36636 21641 36645 21675
rect 36645 21641 36679 21675
rect 36679 21641 36688 21675
rect 36636 21632 36688 21641
rect 34520 21564 34572 21616
rect 12992 21471 13044 21480
rect 12992 21437 13001 21471
rect 13001 21437 13035 21471
rect 13035 21437 13044 21471
rect 12992 21428 13044 21437
rect 15936 21496 15988 21548
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 24676 21539 24728 21548
rect 24676 21505 24685 21539
rect 24685 21505 24719 21539
rect 24719 21505 24728 21539
rect 24676 21496 24728 21505
rect 31576 21496 31628 21548
rect 33140 21496 33192 21548
rect 14280 21428 14332 21480
rect 16672 21428 16724 21480
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 21364 21471 21416 21480
rect 21364 21437 21373 21471
rect 21373 21437 21407 21471
rect 21407 21437 21416 21471
rect 21364 21428 21416 21437
rect 21640 21471 21692 21480
rect 15292 21360 15344 21412
rect 18880 21360 18932 21412
rect 19892 21360 19944 21412
rect 21640 21437 21674 21471
rect 21674 21437 21692 21471
rect 21640 21428 21692 21437
rect 25504 21428 25556 21480
rect 26792 21428 26844 21480
rect 28448 21428 28500 21480
rect 28908 21428 28960 21480
rect 25872 21403 25924 21412
rect 15660 21335 15712 21344
rect 15660 21301 15669 21335
rect 15669 21301 15703 21335
rect 15703 21301 15712 21335
rect 15660 21292 15712 21301
rect 17316 21335 17368 21344
rect 17316 21301 17325 21335
rect 17325 21301 17359 21335
rect 17359 21301 17368 21335
rect 17316 21292 17368 21301
rect 19432 21292 19484 21344
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 23848 21292 23900 21344
rect 25136 21292 25188 21344
rect 25872 21369 25884 21403
rect 25884 21369 25924 21403
rect 25872 21360 25924 21369
rect 30104 21428 30156 21480
rect 31852 21471 31904 21480
rect 31852 21437 31861 21471
rect 31861 21437 31895 21471
rect 31895 21437 31904 21471
rect 31852 21428 31904 21437
rect 33232 21428 33284 21480
rect 33968 21428 34020 21480
rect 34060 21428 34112 21480
rect 34520 21428 34572 21480
rect 34704 21428 34756 21480
rect 34796 21428 34848 21480
rect 29828 21360 29880 21412
rect 30748 21360 30800 21412
rect 31668 21360 31720 21412
rect 27068 21292 27120 21344
rect 27988 21335 28040 21344
rect 27988 21301 27997 21335
rect 27997 21301 28031 21335
rect 28031 21301 28040 21335
rect 27988 21292 28040 21301
rect 31208 21292 31260 21344
rect 33232 21335 33284 21344
rect 33232 21301 33241 21335
rect 33241 21301 33275 21335
rect 33275 21301 33284 21335
rect 33232 21292 33284 21301
rect 34612 21360 34664 21412
rect 35624 21428 35676 21480
rect 35440 21360 35492 21412
rect 33876 21292 33928 21344
rect 35164 21292 35216 21344
rect 35900 21292 35952 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 12808 21088 12860 21140
rect 14188 21088 14240 21140
rect 15660 21088 15712 21140
rect 15936 21131 15988 21140
rect 15936 21097 15945 21131
rect 15945 21097 15979 21131
rect 15979 21097 15988 21131
rect 15936 21088 15988 21097
rect 17684 21088 17736 21140
rect 18144 21088 18196 21140
rect 23756 21088 23808 21140
rect 24032 21088 24084 21140
rect 24492 21088 24544 21140
rect 25228 21131 25280 21140
rect 25228 21097 25237 21131
rect 25237 21097 25271 21131
rect 25271 21097 25280 21131
rect 25228 21088 25280 21097
rect 25596 21088 25648 21140
rect 28632 21088 28684 21140
rect 29736 21088 29788 21140
rect 30104 21088 30156 21140
rect 31576 21131 31628 21140
rect 31576 21097 31585 21131
rect 31585 21097 31619 21131
rect 31619 21097 31628 21131
rect 31576 21088 31628 21097
rect 31852 21088 31904 21140
rect 32956 21131 33008 21140
rect 32956 21097 32965 21131
rect 32965 21097 32999 21131
rect 32999 21097 33008 21131
rect 32956 21088 33008 21097
rect 33600 21088 33652 21140
rect 13084 21020 13136 21072
rect 14740 21020 14792 21072
rect 22744 21020 22796 21072
rect 29184 21020 29236 21072
rect 35164 21088 35216 21140
rect 35624 21131 35676 21140
rect 35624 21097 35633 21131
rect 35633 21097 35667 21131
rect 35667 21097 35676 21131
rect 35624 21088 35676 21097
rect 17316 20952 17368 21004
rect 17960 20952 18012 21004
rect 21180 20995 21232 21004
rect 21180 20961 21189 20995
rect 21189 20961 21223 20995
rect 21223 20961 21232 20995
rect 21180 20952 21232 20961
rect 12992 20927 13044 20936
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 16212 20927 16264 20936
rect 16212 20893 16221 20927
rect 16221 20893 16255 20927
rect 16255 20893 16264 20927
rect 16212 20884 16264 20893
rect 20168 20927 20220 20936
rect 20168 20893 20177 20927
rect 20177 20893 20211 20927
rect 20211 20893 20220 20927
rect 20168 20884 20220 20893
rect 20352 20884 20404 20936
rect 21364 20884 21416 20936
rect 23112 20952 23164 21004
rect 24676 20952 24728 21004
rect 27068 20995 27120 21004
rect 27068 20961 27102 20995
rect 27102 20961 27120 20995
rect 27068 20952 27120 20961
rect 34244 20995 34296 21004
rect 34244 20961 34253 20995
rect 34253 20961 34287 20995
rect 34287 20961 34296 20995
rect 34244 20952 34296 20961
rect 25136 20884 25188 20936
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 21364 20791 21416 20800
rect 21364 20757 21373 20791
rect 21373 20757 21407 20791
rect 21407 20757 21416 20791
rect 21364 20748 21416 20757
rect 26240 20748 26292 20800
rect 27896 20748 27948 20800
rect 33140 20884 33192 20936
rect 33692 20884 33744 20936
rect 33968 20927 34020 20936
rect 33968 20893 33980 20927
rect 33980 20893 34014 20927
rect 34014 20893 34020 20927
rect 33968 20884 34020 20893
rect 29828 20748 29880 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 12992 20544 13044 20596
rect 15292 20587 15344 20596
rect 15292 20553 15301 20587
rect 15301 20553 15335 20587
rect 15335 20553 15344 20587
rect 15292 20544 15344 20553
rect 15844 20544 15896 20596
rect 16212 20544 16264 20596
rect 18052 20544 18104 20596
rect 19432 20587 19484 20596
rect 19432 20553 19441 20587
rect 19441 20553 19475 20587
rect 19475 20553 19484 20587
rect 19432 20544 19484 20553
rect 19984 20544 20036 20596
rect 20904 20544 20956 20596
rect 22744 20544 22796 20596
rect 25228 20544 25280 20596
rect 25596 20544 25648 20596
rect 27620 20587 27672 20596
rect 27620 20553 27629 20587
rect 27629 20553 27663 20587
rect 27663 20553 27672 20587
rect 27620 20544 27672 20553
rect 28724 20544 28776 20596
rect 13084 20519 13136 20528
rect 13084 20485 13093 20519
rect 13093 20485 13127 20519
rect 13127 20485 13136 20519
rect 13084 20476 13136 20485
rect 17316 20476 17368 20528
rect 17868 20476 17920 20528
rect 13636 20340 13688 20392
rect 13912 20383 13964 20392
rect 13912 20349 13921 20383
rect 13921 20349 13955 20383
rect 13955 20349 13964 20383
rect 13912 20340 13964 20349
rect 15936 20408 15988 20460
rect 16948 20408 17000 20460
rect 19524 20519 19576 20528
rect 19524 20485 19533 20519
rect 19533 20485 19567 20519
rect 19567 20485 19576 20519
rect 19524 20476 19576 20485
rect 20076 20451 20128 20460
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 26240 20408 26292 20460
rect 26608 20451 26660 20460
rect 26608 20417 26617 20451
rect 26617 20417 26651 20451
rect 26651 20417 26660 20451
rect 27068 20451 27120 20460
rect 26608 20408 26660 20417
rect 27068 20417 27077 20451
rect 27077 20417 27111 20451
rect 27111 20417 27120 20451
rect 27068 20408 27120 20417
rect 27528 20408 27580 20460
rect 14188 20383 14240 20392
rect 14188 20349 14222 20383
rect 14222 20349 14240 20383
rect 14188 20340 14240 20349
rect 17408 20340 17460 20392
rect 18144 20340 18196 20392
rect 19892 20383 19944 20392
rect 19892 20349 19901 20383
rect 19901 20349 19935 20383
rect 19935 20349 19944 20383
rect 19892 20340 19944 20349
rect 20352 20340 20404 20392
rect 23664 20340 23716 20392
rect 29000 20340 29052 20392
rect 16028 20315 16080 20324
rect 16028 20281 16037 20315
rect 16037 20281 16071 20315
rect 16071 20281 16080 20315
rect 16028 20272 16080 20281
rect 17960 20272 18012 20324
rect 23112 20272 23164 20324
rect 28172 20272 28224 20324
rect 16672 20204 16724 20256
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 20536 20204 20588 20256
rect 23480 20247 23532 20256
rect 23480 20213 23489 20247
rect 23489 20213 23523 20247
rect 23523 20213 23532 20247
rect 23480 20204 23532 20213
rect 23756 20204 23808 20256
rect 26056 20247 26108 20256
rect 26056 20213 26065 20247
rect 26065 20213 26099 20247
rect 26099 20213 26108 20247
rect 26056 20204 26108 20213
rect 28080 20247 28132 20256
rect 28080 20213 28089 20247
rect 28089 20213 28123 20247
rect 28123 20213 28132 20247
rect 28080 20204 28132 20213
rect 29276 20544 29328 20596
rect 33692 20587 33744 20596
rect 33692 20553 33701 20587
rect 33701 20553 33735 20587
rect 33735 20553 33744 20587
rect 33692 20544 33744 20553
rect 33968 20587 34020 20596
rect 33968 20553 33977 20587
rect 33977 20553 34011 20587
rect 34011 20553 34020 20587
rect 33968 20544 34020 20553
rect 34244 20544 34296 20596
rect 34796 20544 34848 20596
rect 36084 20544 36136 20596
rect 29736 20451 29788 20460
rect 29736 20417 29748 20451
rect 29748 20417 29782 20451
rect 29782 20417 29788 20451
rect 29736 20408 29788 20417
rect 31668 20408 31720 20460
rect 31852 20408 31904 20460
rect 29276 20383 29328 20392
rect 29276 20349 29285 20383
rect 29285 20349 29319 20383
rect 29319 20349 29328 20383
rect 29276 20340 29328 20349
rect 29368 20340 29420 20392
rect 30012 20383 30064 20392
rect 30012 20349 30021 20383
rect 30021 20349 30055 20383
rect 30055 20349 30064 20383
rect 30012 20340 30064 20349
rect 31760 20315 31812 20324
rect 31760 20281 31769 20315
rect 31769 20281 31803 20315
rect 31803 20281 31812 20315
rect 31760 20272 31812 20281
rect 35164 20340 35216 20392
rect 35900 20340 35952 20392
rect 35440 20272 35492 20324
rect 29736 20247 29788 20256
rect 29736 20213 29751 20247
rect 29751 20213 29785 20247
rect 29785 20213 29788 20247
rect 31116 20247 31168 20256
rect 29736 20204 29788 20213
rect 31116 20213 31125 20247
rect 31125 20213 31159 20247
rect 31159 20213 31168 20247
rect 31116 20204 31168 20213
rect 32956 20204 33008 20256
rect 33324 20247 33376 20256
rect 33324 20213 33333 20247
rect 33333 20213 33367 20247
rect 33367 20213 33376 20247
rect 33324 20204 33376 20213
rect 36084 20204 36136 20256
rect 37280 20247 37332 20256
rect 37280 20213 37289 20247
rect 37289 20213 37323 20247
rect 37323 20213 37332 20247
rect 37280 20204 37332 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 17868 20000 17920 20052
rect 19984 20000 20036 20052
rect 21180 20043 21232 20052
rect 21180 20009 21189 20043
rect 21189 20009 21223 20043
rect 21223 20009 21232 20043
rect 21180 20000 21232 20009
rect 23664 20043 23716 20052
rect 23664 20009 23673 20043
rect 23673 20009 23707 20043
rect 23707 20009 23716 20043
rect 23664 20000 23716 20009
rect 24032 20043 24084 20052
rect 24032 20009 24041 20043
rect 24041 20009 24075 20043
rect 24075 20009 24084 20043
rect 24032 20000 24084 20009
rect 25136 20043 25188 20052
rect 25136 20009 25145 20043
rect 25145 20009 25179 20043
rect 25179 20009 25188 20043
rect 25136 20000 25188 20009
rect 26608 20000 26660 20052
rect 29000 20043 29052 20052
rect 29000 20009 29009 20043
rect 29009 20009 29043 20043
rect 29043 20009 29052 20043
rect 29000 20000 29052 20009
rect 31576 20000 31628 20052
rect 31852 20000 31904 20052
rect 33232 20000 33284 20052
rect 33692 20000 33744 20052
rect 34336 20000 34388 20052
rect 35164 20043 35216 20052
rect 35164 20009 35173 20043
rect 35173 20009 35207 20043
rect 35207 20009 35216 20043
rect 35164 20000 35216 20009
rect 16028 19932 16080 19984
rect 16212 19932 16264 19984
rect 17592 19932 17644 19984
rect 19892 19975 19944 19984
rect 19892 19941 19901 19975
rect 19901 19941 19935 19975
rect 19935 19941 19944 19975
rect 19892 19932 19944 19941
rect 24308 19932 24360 19984
rect 22100 19864 22152 19916
rect 22284 19907 22336 19916
rect 22284 19873 22293 19907
rect 22293 19873 22327 19907
rect 22327 19873 22336 19907
rect 22284 19864 22336 19873
rect 24400 19907 24452 19916
rect 24400 19873 24409 19907
rect 24409 19873 24443 19907
rect 24443 19873 24452 19907
rect 24400 19864 24452 19873
rect 14556 19796 14608 19848
rect 22192 19796 22244 19848
rect 22560 19839 22612 19848
rect 22560 19805 22569 19839
rect 22569 19805 22603 19839
rect 22603 19805 22612 19839
rect 22560 19796 22612 19805
rect 24032 19796 24084 19848
rect 28080 19932 28132 19984
rect 30104 19975 30156 19984
rect 30104 19941 30138 19975
rect 30138 19941 30156 19975
rect 30104 19932 30156 19941
rect 26516 19907 26568 19916
rect 26516 19873 26525 19907
rect 26525 19873 26559 19907
rect 26559 19873 26568 19907
rect 26516 19864 26568 19873
rect 27896 19907 27948 19916
rect 27896 19873 27930 19907
rect 27930 19873 27948 19907
rect 27896 19864 27948 19873
rect 29828 19907 29880 19916
rect 29828 19873 29837 19907
rect 29837 19873 29871 19907
rect 29871 19873 29880 19907
rect 29828 19864 29880 19873
rect 35992 19907 36044 19916
rect 26792 19796 26844 19848
rect 27620 19839 27672 19848
rect 27620 19805 27629 19839
rect 27629 19805 27663 19839
rect 27663 19805 27672 19839
rect 27620 19796 27672 19805
rect 33416 19796 33468 19848
rect 33692 19839 33744 19848
rect 33692 19805 33701 19839
rect 33701 19805 33735 19839
rect 33735 19805 33744 19839
rect 33692 19796 33744 19805
rect 34428 19728 34480 19780
rect 35992 19873 36001 19907
rect 36001 19873 36035 19907
rect 36035 19873 36044 19907
rect 35992 19864 36044 19873
rect 19984 19660 20036 19712
rect 20536 19703 20588 19712
rect 20536 19669 20545 19703
rect 20545 19669 20579 19703
rect 20579 19669 20588 19703
rect 20536 19660 20588 19669
rect 26240 19660 26292 19712
rect 29368 19703 29420 19712
rect 29368 19669 29377 19703
rect 29377 19669 29411 19703
rect 29411 19669 29420 19703
rect 29368 19660 29420 19669
rect 32956 19660 33008 19712
rect 36912 19796 36964 19848
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 16028 19456 16080 19508
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 18052 19456 18104 19508
rect 13912 19320 13964 19372
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 20352 19456 20404 19508
rect 22192 19456 22244 19508
rect 26516 19499 26568 19508
rect 26516 19465 26525 19499
rect 26525 19465 26559 19499
rect 26559 19465 26568 19499
rect 26516 19456 26568 19465
rect 27896 19499 27948 19508
rect 27896 19465 27905 19499
rect 27905 19465 27939 19499
rect 27939 19465 27948 19499
rect 27896 19456 27948 19465
rect 33048 19499 33100 19508
rect 22560 19320 22612 19372
rect 28172 19363 28224 19372
rect 15108 19252 15160 19304
rect 22008 19252 22060 19304
rect 24124 19252 24176 19304
rect 24584 19252 24636 19304
rect 28172 19329 28181 19363
rect 28181 19329 28215 19363
rect 28215 19329 28224 19363
rect 28172 19320 28224 19329
rect 29736 19320 29788 19372
rect 30288 19320 30340 19372
rect 30472 19320 30524 19372
rect 25780 19295 25832 19304
rect 19892 19227 19944 19236
rect 19892 19193 19901 19227
rect 19901 19193 19935 19227
rect 19935 19193 19944 19227
rect 19892 19184 19944 19193
rect 21180 19184 21232 19236
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 26884 19295 26936 19304
rect 26884 19261 26893 19295
rect 26893 19261 26927 19295
rect 26927 19261 26936 19295
rect 26884 19252 26936 19261
rect 14556 19116 14608 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 20536 19116 20588 19168
rect 23296 19116 23348 19168
rect 24032 19159 24084 19168
rect 24032 19125 24041 19159
rect 24041 19125 24075 19159
rect 24075 19125 24084 19159
rect 24032 19116 24084 19125
rect 24216 19159 24268 19168
rect 24216 19125 24225 19159
rect 24225 19125 24259 19159
rect 24259 19125 24268 19159
rect 24216 19116 24268 19125
rect 24492 19116 24544 19168
rect 24676 19159 24728 19168
rect 24676 19125 24685 19159
rect 24685 19125 24719 19159
rect 24719 19125 24728 19159
rect 24676 19116 24728 19125
rect 25780 19116 25832 19168
rect 29276 19252 29328 19304
rect 31116 19320 31168 19372
rect 29184 19184 29236 19236
rect 30748 19252 30800 19304
rect 33048 19465 33057 19499
rect 33057 19465 33091 19499
rect 33091 19465 33100 19499
rect 33048 19456 33100 19465
rect 33232 19456 33284 19508
rect 33416 19320 33468 19372
rect 35440 19363 35492 19372
rect 35440 19329 35449 19363
rect 35449 19329 35483 19363
rect 35483 19329 35492 19363
rect 35440 19320 35492 19329
rect 33784 19227 33836 19236
rect 27068 19159 27120 19168
rect 27068 19125 27077 19159
rect 27077 19125 27111 19159
rect 27111 19125 27120 19159
rect 27068 19116 27120 19125
rect 28632 19159 28684 19168
rect 28632 19125 28641 19159
rect 28641 19125 28675 19159
rect 28675 19125 28684 19159
rect 28632 19116 28684 19125
rect 30288 19116 30340 19168
rect 30748 19116 30800 19168
rect 30932 19116 30984 19168
rect 33784 19193 33793 19227
rect 33793 19193 33827 19227
rect 33827 19193 33836 19227
rect 33784 19184 33836 19193
rect 35992 19252 36044 19304
rect 36084 19184 36136 19236
rect 33692 19116 33744 19168
rect 34060 19116 34112 19168
rect 36912 19116 36964 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 14556 18955 14608 18964
rect 14556 18921 14565 18955
rect 14565 18921 14599 18955
rect 14599 18921 14608 18955
rect 14556 18912 14608 18921
rect 16028 18912 16080 18964
rect 22284 18912 22336 18964
rect 23388 18912 23440 18964
rect 24400 18912 24452 18964
rect 24676 18912 24728 18964
rect 25688 18912 25740 18964
rect 26700 18955 26752 18964
rect 26700 18921 26709 18955
rect 26709 18921 26743 18955
rect 26743 18921 26752 18955
rect 26700 18912 26752 18921
rect 27804 18912 27856 18964
rect 28080 18912 28132 18964
rect 29184 18955 29236 18964
rect 29184 18921 29193 18955
rect 29193 18921 29227 18955
rect 29227 18921 29236 18955
rect 29184 18912 29236 18921
rect 29920 18955 29972 18964
rect 29920 18921 29929 18955
rect 29929 18921 29963 18955
rect 29963 18921 29972 18955
rect 29920 18912 29972 18921
rect 30472 18912 30524 18964
rect 30932 18912 30984 18964
rect 31668 18912 31720 18964
rect 33232 18912 33284 18964
rect 34152 18912 34204 18964
rect 35716 18912 35768 18964
rect 37188 18912 37240 18964
rect 19340 18844 19392 18896
rect 19892 18844 19944 18896
rect 29460 18844 29512 18896
rect 36176 18844 36228 18896
rect 19616 18819 19668 18828
rect 19616 18785 19625 18819
rect 19625 18785 19659 18819
rect 19659 18785 19668 18819
rect 19616 18776 19668 18785
rect 20536 18776 20588 18828
rect 21548 18776 21600 18828
rect 23848 18776 23900 18828
rect 25136 18819 25188 18828
rect 25136 18785 25145 18819
rect 25145 18785 25179 18819
rect 25179 18785 25188 18819
rect 25136 18776 25188 18785
rect 26516 18819 26568 18828
rect 26516 18785 26525 18819
rect 26525 18785 26559 18819
rect 26559 18785 26568 18819
rect 26516 18776 26568 18785
rect 27712 18776 27764 18828
rect 34060 18776 34112 18828
rect 35900 18776 35952 18828
rect 19984 18708 20036 18760
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 23664 18751 23716 18760
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 25228 18751 25280 18760
rect 23664 18708 23716 18717
rect 25228 18717 25237 18751
rect 25237 18717 25271 18751
rect 25271 18717 25280 18751
rect 25228 18708 25280 18717
rect 22468 18640 22520 18692
rect 26148 18708 26200 18760
rect 27620 18708 27672 18760
rect 31024 18751 31076 18760
rect 27896 18640 27948 18692
rect 31024 18717 31033 18751
rect 31033 18717 31067 18751
rect 31067 18717 31076 18751
rect 31024 18708 31076 18717
rect 33784 18708 33836 18760
rect 36084 18708 36136 18760
rect 31208 18640 31260 18692
rect 34428 18640 34480 18692
rect 19248 18615 19300 18624
rect 19248 18581 19257 18615
rect 19257 18581 19291 18615
rect 19291 18581 19300 18615
rect 19248 18572 19300 18581
rect 22100 18572 22152 18624
rect 32772 18615 32824 18624
rect 32772 18581 32781 18615
rect 32781 18581 32815 18615
rect 32815 18581 32824 18615
rect 32772 18572 32824 18581
rect 35624 18615 35676 18624
rect 35624 18581 35633 18615
rect 35633 18581 35667 18615
rect 35667 18581 35676 18615
rect 35624 18572 35676 18581
rect 37096 18572 37148 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 19340 18411 19392 18420
rect 19340 18377 19349 18411
rect 19349 18377 19383 18411
rect 19383 18377 19392 18411
rect 19340 18368 19392 18377
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 21180 18411 21232 18420
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 22008 18411 22060 18420
rect 22008 18377 22017 18411
rect 22017 18377 22051 18411
rect 22051 18377 22060 18411
rect 22008 18368 22060 18377
rect 22284 18368 22336 18420
rect 23572 18368 23624 18420
rect 25228 18368 25280 18420
rect 26240 18368 26292 18420
rect 27712 18368 27764 18420
rect 27896 18368 27948 18420
rect 29184 18368 29236 18420
rect 29460 18411 29512 18420
rect 29460 18377 29469 18411
rect 29469 18377 29503 18411
rect 29503 18377 29512 18411
rect 29460 18368 29512 18377
rect 30932 18368 30984 18420
rect 31024 18368 31076 18420
rect 33784 18411 33836 18420
rect 33784 18377 33793 18411
rect 33793 18377 33827 18411
rect 33827 18377 33836 18411
rect 33784 18368 33836 18377
rect 34060 18411 34112 18420
rect 34060 18377 34069 18411
rect 34069 18377 34103 18411
rect 34103 18377 34112 18411
rect 34060 18368 34112 18377
rect 34152 18368 34204 18420
rect 35716 18411 35768 18420
rect 35716 18377 35725 18411
rect 35725 18377 35759 18411
rect 35759 18377 35768 18411
rect 35716 18368 35768 18377
rect 35900 18368 35952 18420
rect 36176 18368 36228 18420
rect 24216 18300 24268 18352
rect 26516 18300 26568 18352
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 22560 18275 22612 18284
rect 22560 18241 22569 18275
rect 22569 18241 22603 18275
rect 22603 18241 22612 18275
rect 22560 18232 22612 18241
rect 28632 18232 28684 18284
rect 30472 18232 30524 18284
rect 32404 18232 32456 18284
rect 19892 18164 19944 18216
rect 22376 18207 22428 18216
rect 22376 18173 22385 18207
rect 22385 18173 22419 18207
rect 22419 18173 22428 18207
rect 22376 18164 22428 18173
rect 23848 18207 23900 18216
rect 23848 18173 23857 18207
rect 23857 18173 23891 18207
rect 23891 18173 23900 18207
rect 23848 18164 23900 18173
rect 25688 18164 25740 18216
rect 32772 18164 32824 18216
rect 20076 18139 20128 18148
rect 20076 18105 20110 18139
rect 20110 18105 20128 18139
rect 20076 18096 20128 18105
rect 23664 18096 23716 18148
rect 24400 18139 24452 18148
rect 24400 18105 24409 18139
rect 24409 18105 24443 18139
rect 24443 18105 24452 18139
rect 24400 18096 24452 18105
rect 33416 18096 33468 18148
rect 34152 18096 34204 18148
rect 34704 18096 34756 18148
rect 18604 18071 18656 18080
rect 18604 18037 18613 18071
rect 18613 18037 18647 18071
rect 18647 18037 18656 18071
rect 18604 18028 18656 18037
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 25228 18071 25280 18080
rect 25228 18037 25237 18071
rect 25237 18037 25271 18071
rect 25271 18037 25280 18071
rect 25228 18028 25280 18037
rect 32680 18071 32732 18080
rect 32680 18037 32689 18071
rect 32689 18037 32723 18071
rect 32723 18037 32732 18071
rect 32680 18028 32732 18037
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 22284 17867 22336 17876
rect 22284 17833 22293 17867
rect 22293 17833 22327 17867
rect 22327 17833 22336 17867
rect 22284 17824 22336 17833
rect 22376 17824 22428 17876
rect 23388 17824 23440 17876
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 27896 17867 27948 17876
rect 27896 17833 27905 17867
rect 27905 17833 27939 17867
rect 27939 17833 27948 17867
rect 27896 17824 27948 17833
rect 34244 17824 34296 17876
rect 18972 17756 19024 17808
rect 21364 17756 21416 17808
rect 25228 17756 25280 17808
rect 26240 17756 26292 17808
rect 26700 17756 26752 17808
rect 22560 17688 22612 17740
rect 23112 17731 23164 17740
rect 23112 17697 23121 17731
rect 23121 17697 23155 17731
rect 23155 17697 23164 17731
rect 23112 17688 23164 17697
rect 24308 17688 24360 17740
rect 27068 17688 27120 17740
rect 32496 17731 32548 17740
rect 32496 17697 32505 17731
rect 32505 17697 32539 17731
rect 32539 17697 32548 17731
rect 32496 17688 32548 17697
rect 32864 17688 32916 17740
rect 33324 17688 33376 17740
rect 36544 17688 36596 17740
rect 19616 17620 19668 17672
rect 19984 17620 20036 17672
rect 20904 17663 20956 17672
rect 19248 17527 19300 17536
rect 19248 17493 19257 17527
rect 19257 17493 19291 17527
rect 19291 17493 19300 17527
rect 19248 17484 19300 17493
rect 19892 17484 19944 17536
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 30380 17620 30432 17672
rect 32680 17663 32732 17672
rect 32680 17629 32689 17663
rect 32689 17629 32723 17663
rect 32723 17629 32732 17663
rect 32680 17620 32732 17629
rect 34888 17663 34940 17672
rect 34888 17629 34897 17663
rect 34897 17629 34931 17663
rect 34931 17629 34940 17663
rect 34888 17620 34940 17629
rect 29920 17552 29972 17604
rect 24860 17484 24912 17536
rect 29736 17527 29788 17536
rect 29736 17493 29745 17527
rect 29745 17493 29779 17527
rect 29779 17493 29788 17527
rect 29736 17484 29788 17493
rect 31668 17527 31720 17536
rect 31668 17493 31677 17527
rect 31677 17493 31711 17527
rect 31711 17493 31720 17527
rect 31668 17484 31720 17493
rect 32128 17527 32180 17536
rect 32128 17493 32137 17527
rect 32137 17493 32171 17527
rect 32171 17493 32180 17527
rect 32128 17484 32180 17493
rect 34336 17527 34388 17536
rect 34336 17493 34345 17527
rect 34345 17493 34379 17527
rect 34379 17493 34388 17527
rect 34336 17484 34388 17493
rect 35348 17484 35400 17536
rect 35992 17484 36044 17536
rect 36084 17527 36136 17536
rect 36084 17493 36093 17527
rect 36093 17493 36127 17527
rect 36127 17493 36136 17527
rect 36084 17484 36136 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 21088 17323 21140 17332
rect 21088 17289 21097 17323
rect 21097 17289 21131 17323
rect 21131 17289 21140 17323
rect 21088 17280 21140 17289
rect 25228 17323 25280 17332
rect 25228 17289 25237 17323
rect 25237 17289 25271 17323
rect 25271 17289 25280 17323
rect 25228 17280 25280 17289
rect 26700 17323 26752 17332
rect 26700 17289 26709 17323
rect 26709 17289 26743 17323
rect 26743 17289 26752 17323
rect 26700 17280 26752 17289
rect 28724 17323 28776 17332
rect 28724 17289 28733 17323
rect 28733 17289 28767 17323
rect 28767 17289 28776 17323
rect 28724 17280 28776 17289
rect 34244 17280 34296 17332
rect 34612 17280 34664 17332
rect 36544 17323 36596 17332
rect 36544 17289 36553 17323
rect 36553 17289 36587 17323
rect 36587 17289 36596 17323
rect 36544 17280 36596 17289
rect 23112 17212 23164 17264
rect 30472 17212 30524 17264
rect 35164 17212 35216 17264
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 29736 17144 29788 17196
rect 34336 17144 34388 17196
rect 20352 17076 20404 17128
rect 22284 17119 22336 17128
rect 22284 17085 22293 17119
rect 22293 17085 22327 17119
rect 22327 17085 22336 17119
rect 22284 17076 22336 17085
rect 23848 17119 23900 17128
rect 23848 17085 23857 17119
rect 23857 17085 23891 17119
rect 23891 17085 23900 17119
rect 23848 17076 23900 17085
rect 25964 17076 26016 17128
rect 28172 17119 28224 17128
rect 28172 17085 28181 17119
rect 28181 17085 28215 17119
rect 28215 17085 28224 17119
rect 28172 17076 28224 17085
rect 28908 17076 28960 17128
rect 19616 17008 19668 17060
rect 19892 17008 19944 17060
rect 21732 17051 21784 17060
rect 21732 17017 21741 17051
rect 21741 17017 21775 17051
rect 21775 17017 21784 17051
rect 21732 17008 21784 17017
rect 24860 17008 24912 17060
rect 25504 17008 25556 17060
rect 28724 17008 28776 17060
rect 18604 16983 18656 16992
rect 18604 16949 18613 16983
rect 18613 16949 18647 16983
rect 18647 16949 18656 16983
rect 18604 16940 18656 16949
rect 35992 17187 36044 17196
rect 35992 17153 36001 17187
rect 36001 17153 36035 17187
rect 36035 17153 36044 17187
rect 35992 17144 36044 17153
rect 31392 17051 31444 17060
rect 31392 17017 31401 17051
rect 31401 17017 31435 17051
rect 31435 17017 31444 17051
rect 31392 17008 31444 17017
rect 31668 17008 31720 17060
rect 31852 17051 31904 17060
rect 31852 17017 31886 17051
rect 31886 17017 31904 17051
rect 31852 17008 31904 17017
rect 32864 17008 32916 17060
rect 34428 17008 34480 17060
rect 20260 16940 20312 16992
rect 21364 16983 21416 16992
rect 21364 16949 21373 16983
rect 21373 16949 21407 16983
rect 21407 16949 21416 16983
rect 21364 16940 21416 16949
rect 27068 16940 27120 16992
rect 29000 16983 29052 16992
rect 29000 16949 29009 16983
rect 29009 16949 29043 16983
rect 29043 16949 29052 16983
rect 29000 16940 29052 16949
rect 29920 16940 29972 16992
rect 31116 16983 31168 16992
rect 31116 16949 31125 16983
rect 31125 16949 31159 16983
rect 31159 16949 31168 16983
rect 31116 16940 31168 16949
rect 32680 16940 32732 16992
rect 33324 16940 33376 16992
rect 35440 16983 35492 16992
rect 35440 16949 35449 16983
rect 35449 16949 35483 16983
rect 35483 16949 35492 16983
rect 35440 16940 35492 16949
rect 35900 16940 35952 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 22560 16779 22612 16788
rect 22560 16745 22569 16779
rect 22569 16745 22603 16779
rect 22603 16745 22612 16779
rect 22560 16736 22612 16745
rect 23112 16779 23164 16788
rect 23112 16745 23121 16779
rect 23121 16745 23155 16779
rect 23155 16745 23164 16779
rect 23112 16736 23164 16745
rect 23848 16736 23900 16788
rect 24308 16779 24360 16788
rect 24308 16745 24317 16779
rect 24317 16745 24351 16779
rect 24351 16745 24360 16779
rect 24308 16736 24360 16745
rect 24492 16736 24544 16788
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25504 16779 25556 16788
rect 25504 16745 25513 16779
rect 25513 16745 25547 16779
rect 25547 16745 25556 16779
rect 25504 16736 25556 16745
rect 25964 16736 26016 16788
rect 27068 16779 27120 16788
rect 27068 16745 27077 16779
rect 27077 16745 27111 16779
rect 27111 16745 27120 16779
rect 27068 16736 27120 16745
rect 27436 16779 27488 16788
rect 27436 16745 27445 16779
rect 27445 16745 27479 16779
rect 27479 16745 27488 16779
rect 27436 16736 27488 16745
rect 29736 16779 29788 16788
rect 29736 16745 29745 16779
rect 29745 16745 29779 16779
rect 29779 16745 29788 16779
rect 29736 16736 29788 16745
rect 32128 16736 32180 16788
rect 32496 16736 32548 16788
rect 33048 16736 33100 16788
rect 33140 16736 33192 16788
rect 34244 16736 34296 16788
rect 34796 16736 34848 16788
rect 19892 16668 19944 16720
rect 25228 16668 25280 16720
rect 28172 16668 28224 16720
rect 35992 16736 36044 16788
rect 35716 16711 35768 16720
rect 35716 16677 35728 16711
rect 35728 16677 35768 16711
rect 35716 16668 35768 16677
rect 19616 16643 19668 16652
rect 19616 16609 19625 16643
rect 19625 16609 19659 16643
rect 19659 16609 19668 16643
rect 19616 16600 19668 16609
rect 21732 16600 21784 16652
rect 27528 16600 27580 16652
rect 29000 16600 29052 16652
rect 30564 16643 30616 16652
rect 30564 16609 30573 16643
rect 30573 16609 30607 16643
rect 30607 16609 30616 16643
rect 30564 16600 30616 16609
rect 32036 16600 32088 16652
rect 33140 16600 33192 16652
rect 33416 16600 33468 16652
rect 35256 16600 35308 16652
rect 35992 16600 36044 16652
rect 19340 16532 19392 16584
rect 19984 16532 20036 16584
rect 24400 16532 24452 16584
rect 33232 16575 33284 16584
rect 33232 16541 33244 16575
rect 33244 16541 33278 16575
rect 33278 16541 33284 16575
rect 33232 16532 33284 16541
rect 20812 16396 20864 16448
rect 33232 16396 33284 16448
rect 35440 16396 35492 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 19340 16235 19392 16244
rect 19340 16201 19349 16235
rect 19349 16201 19383 16235
rect 19383 16201 19392 16235
rect 19340 16192 19392 16201
rect 19616 16235 19668 16244
rect 19616 16201 19625 16235
rect 19625 16201 19659 16235
rect 19659 16201 19668 16235
rect 19616 16192 19668 16201
rect 21364 16235 21416 16244
rect 21364 16201 21373 16235
rect 21373 16201 21407 16235
rect 21407 16201 21416 16235
rect 21364 16192 21416 16201
rect 24400 16192 24452 16244
rect 24768 16192 24820 16244
rect 25228 16235 25280 16244
rect 25228 16201 25237 16235
rect 25237 16201 25271 16235
rect 25271 16201 25280 16235
rect 25228 16192 25280 16201
rect 28172 16192 28224 16244
rect 32496 16192 32548 16244
rect 32956 16192 33008 16244
rect 33416 16192 33468 16244
rect 35348 16235 35400 16244
rect 35348 16201 35357 16235
rect 35357 16201 35391 16235
rect 35391 16201 35400 16235
rect 35348 16192 35400 16201
rect 20996 16056 21048 16108
rect 22192 16056 22244 16108
rect 32036 16099 32088 16108
rect 32036 16065 32045 16099
rect 32045 16065 32079 16099
rect 32079 16065 32088 16099
rect 32036 16056 32088 16065
rect 32220 16056 32272 16108
rect 33232 16056 33284 16108
rect 19892 15988 19944 16040
rect 20260 16031 20312 16040
rect 20260 15997 20294 16031
rect 20294 15997 20312 16031
rect 20260 15988 20312 15997
rect 24860 15988 24912 16040
rect 27068 15988 27120 16040
rect 29000 15988 29052 16040
rect 29552 16031 29604 16040
rect 29552 15997 29561 16031
rect 29561 15997 29595 16031
rect 29595 15997 29604 16031
rect 29552 15988 29604 15997
rect 32588 15988 32640 16040
rect 34336 15988 34388 16040
rect 35440 16031 35492 16040
rect 35440 15997 35449 16031
rect 35449 15997 35483 16031
rect 35483 15997 35492 16031
rect 35440 15988 35492 15997
rect 20812 15920 20864 15972
rect 18604 15852 18656 15904
rect 19984 15852 20036 15904
rect 29736 15920 29788 15972
rect 21732 15895 21784 15904
rect 21732 15861 21741 15895
rect 21741 15861 21775 15895
rect 21775 15861 21784 15895
rect 21732 15852 21784 15861
rect 22192 15852 22244 15904
rect 24308 15852 24360 15904
rect 25412 15852 25464 15904
rect 25688 15895 25740 15904
rect 25688 15861 25697 15895
rect 25697 15861 25731 15895
rect 25731 15861 25740 15895
rect 25688 15852 25740 15861
rect 26792 15895 26844 15904
rect 26792 15861 26801 15895
rect 26801 15861 26835 15895
rect 26835 15861 26844 15895
rect 26792 15852 26844 15861
rect 30932 15895 30984 15904
rect 30932 15861 30941 15895
rect 30941 15861 30975 15895
rect 30975 15861 30984 15895
rect 30932 15852 30984 15861
rect 31208 15852 31260 15904
rect 32496 15895 32548 15904
rect 32496 15861 32511 15895
rect 32511 15861 32545 15895
rect 32545 15861 32548 15895
rect 36820 15895 36872 15904
rect 32496 15852 32548 15861
rect 36820 15861 36829 15895
rect 36829 15861 36863 15895
rect 36863 15861 36872 15895
rect 36820 15852 36872 15861
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 20260 15648 20312 15700
rect 21732 15648 21784 15700
rect 24308 15648 24360 15700
rect 24860 15691 24912 15700
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 25688 15648 25740 15700
rect 26700 15648 26752 15700
rect 27620 15691 27672 15700
rect 27620 15657 27629 15691
rect 27629 15657 27663 15691
rect 27663 15657 27672 15691
rect 28724 15691 28776 15700
rect 27620 15648 27672 15657
rect 28724 15657 28733 15691
rect 28733 15657 28767 15691
rect 28767 15657 28776 15691
rect 28724 15648 28776 15657
rect 29736 15648 29788 15700
rect 30380 15648 30432 15700
rect 31024 15648 31076 15700
rect 32036 15648 32088 15700
rect 35716 15648 35768 15700
rect 19340 15580 19392 15632
rect 20904 15580 20956 15632
rect 22008 15580 22060 15632
rect 25964 15623 26016 15632
rect 25964 15589 25973 15623
rect 25973 15589 26007 15623
rect 26007 15589 26016 15623
rect 25964 15580 26016 15589
rect 27068 15580 27120 15632
rect 28632 15623 28684 15632
rect 28632 15589 28641 15623
rect 28641 15589 28675 15623
rect 28675 15589 28684 15623
rect 28632 15580 28684 15589
rect 30472 15580 30524 15632
rect 32404 15580 32456 15632
rect 35900 15648 35952 15700
rect 24676 15512 24728 15564
rect 25872 15512 25924 15564
rect 34244 15512 34296 15564
rect 20812 15444 20864 15496
rect 24952 15444 25004 15496
rect 25412 15444 25464 15496
rect 26148 15444 26200 15496
rect 27712 15444 27764 15496
rect 29000 15444 29052 15496
rect 30932 15487 30984 15496
rect 30932 15453 30941 15487
rect 30941 15453 30975 15487
rect 30975 15453 30984 15487
rect 30932 15444 30984 15453
rect 33876 15444 33928 15496
rect 34336 15444 34388 15496
rect 28632 15376 28684 15428
rect 29552 15376 29604 15428
rect 31116 15376 31168 15428
rect 28816 15308 28868 15360
rect 30288 15351 30340 15360
rect 30288 15317 30297 15351
rect 30297 15317 30331 15351
rect 30331 15317 30340 15351
rect 30288 15308 30340 15317
rect 32588 15308 32640 15360
rect 34244 15308 34296 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 20904 15147 20956 15156
rect 20904 15113 20913 15147
rect 20913 15113 20947 15147
rect 20947 15113 20956 15147
rect 20904 15104 20956 15113
rect 24952 15147 25004 15156
rect 24952 15113 24961 15147
rect 24961 15113 24995 15147
rect 24995 15113 25004 15147
rect 24952 15104 25004 15113
rect 27712 15104 27764 15156
rect 28448 15147 28500 15156
rect 28448 15113 28457 15147
rect 28457 15113 28491 15147
rect 28491 15113 28500 15147
rect 28448 15104 28500 15113
rect 28724 15147 28776 15156
rect 28724 15113 28733 15147
rect 28733 15113 28767 15147
rect 28767 15113 28776 15147
rect 28724 15104 28776 15113
rect 29000 15104 29052 15156
rect 30380 15147 30432 15156
rect 30380 15113 30389 15147
rect 30389 15113 30423 15147
rect 30423 15113 30432 15147
rect 30380 15104 30432 15113
rect 30932 15104 30984 15156
rect 20812 15036 20864 15088
rect 22100 14764 22152 14816
rect 25320 14968 25372 15020
rect 32404 15104 32456 15156
rect 33140 15104 33192 15156
rect 34244 15147 34296 15156
rect 34244 15113 34253 15147
rect 34253 15113 34287 15147
rect 34287 15113 34296 15147
rect 34244 15104 34296 15113
rect 34428 15104 34480 15156
rect 25412 14943 25464 14952
rect 25412 14909 25421 14943
rect 25421 14909 25455 14943
rect 25455 14909 25464 14943
rect 25412 14900 25464 14909
rect 25964 14900 26016 14952
rect 28448 14900 28500 14952
rect 29000 14900 29052 14952
rect 31116 14900 31168 14952
rect 33048 14968 33100 15020
rect 34244 14968 34296 15020
rect 25596 14832 25648 14884
rect 23480 14807 23532 14816
rect 23480 14773 23489 14807
rect 23489 14773 23523 14807
rect 23523 14773 23532 14807
rect 23480 14764 23532 14773
rect 24216 14807 24268 14816
rect 24216 14773 24225 14807
rect 24225 14773 24259 14807
rect 24259 14773 24268 14807
rect 24216 14764 24268 14773
rect 26240 14764 26292 14816
rect 26792 14807 26844 14816
rect 26792 14773 26801 14807
rect 26801 14773 26835 14807
rect 26835 14773 26844 14807
rect 26792 14764 26844 14773
rect 27068 14807 27120 14816
rect 27068 14773 27077 14807
rect 27077 14773 27111 14807
rect 27111 14773 27120 14807
rect 27068 14764 27120 14773
rect 27620 14764 27672 14816
rect 34704 14832 34756 14884
rect 35164 14832 35216 14884
rect 31484 14764 31536 14816
rect 33876 14807 33928 14816
rect 33876 14773 33885 14807
rect 33885 14773 33919 14807
rect 33919 14773 33928 14807
rect 33876 14764 33928 14773
rect 35532 14764 35584 14816
rect 35992 14764 36044 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 23296 14603 23348 14612
rect 23296 14569 23305 14603
rect 23305 14569 23339 14603
rect 23339 14569 23348 14603
rect 23296 14560 23348 14569
rect 24216 14560 24268 14612
rect 25596 14603 25648 14612
rect 25596 14569 25605 14603
rect 25605 14569 25639 14603
rect 25639 14569 25648 14603
rect 25596 14560 25648 14569
rect 26700 14603 26752 14612
rect 26700 14569 26709 14603
rect 26709 14569 26743 14603
rect 26743 14569 26752 14603
rect 26700 14560 26752 14569
rect 27528 14560 27580 14612
rect 28632 14560 28684 14612
rect 29000 14560 29052 14612
rect 29920 14603 29972 14612
rect 29920 14569 29929 14603
rect 29929 14569 29963 14603
rect 29963 14569 29972 14603
rect 29920 14560 29972 14569
rect 30472 14560 30524 14612
rect 32864 14560 32916 14612
rect 34244 14560 34296 14612
rect 35164 14560 35216 14612
rect 25320 14492 25372 14544
rect 26424 14492 26476 14544
rect 28816 14492 28868 14544
rect 23112 14467 23164 14476
rect 23112 14433 23121 14467
rect 23121 14433 23155 14467
rect 23155 14433 23164 14467
rect 23112 14424 23164 14433
rect 23664 14424 23716 14476
rect 24308 14424 24360 14476
rect 27160 14424 27212 14476
rect 29092 14424 29144 14476
rect 32772 14492 32824 14544
rect 31300 14424 31352 14476
rect 32588 14467 32640 14476
rect 32588 14433 32597 14467
rect 32597 14433 32631 14467
rect 32631 14433 32640 14467
rect 32588 14424 32640 14433
rect 27528 14399 27580 14408
rect 27528 14365 27537 14399
rect 27537 14365 27571 14399
rect 27571 14365 27580 14399
rect 27528 14356 27580 14365
rect 27712 14399 27764 14408
rect 27712 14365 27721 14399
rect 27721 14365 27755 14399
rect 27755 14365 27764 14399
rect 27712 14356 27764 14365
rect 32956 14356 33008 14408
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 24124 14220 24176 14272
rect 24400 14220 24452 14272
rect 27896 14220 27948 14272
rect 30380 14263 30432 14272
rect 30380 14229 30389 14263
rect 30389 14229 30423 14263
rect 30423 14229 30432 14263
rect 30380 14220 30432 14229
rect 31484 14220 31536 14272
rect 33508 14220 33560 14272
rect 33876 14220 33928 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 24308 14016 24360 14068
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 25596 14016 25648 14068
rect 25872 14059 25924 14068
rect 21364 13923 21416 13932
rect 21364 13889 21373 13923
rect 21373 13889 21407 13923
rect 21407 13889 21416 13923
rect 21364 13880 21416 13889
rect 25872 14025 25881 14059
rect 25881 14025 25915 14059
rect 25915 14025 25924 14059
rect 25872 14016 25924 14025
rect 27528 14016 27580 14068
rect 27712 14016 27764 14068
rect 29092 14059 29144 14068
rect 29092 14025 29101 14059
rect 29101 14025 29135 14059
rect 29135 14025 29144 14059
rect 29092 14016 29144 14025
rect 29184 14016 29236 14068
rect 31300 14059 31352 14068
rect 27896 13948 27948 14000
rect 28540 13991 28592 14000
rect 28540 13957 28549 13991
rect 28549 13957 28583 13991
rect 28583 13957 28592 13991
rect 28540 13948 28592 13957
rect 23112 13855 23164 13864
rect 23112 13821 23121 13855
rect 23121 13821 23155 13855
rect 23155 13821 23164 13855
rect 23664 13855 23716 13864
rect 23112 13812 23164 13821
rect 21272 13787 21324 13796
rect 21272 13753 21281 13787
rect 21281 13753 21315 13787
rect 21315 13753 21324 13787
rect 21640 13787 21692 13796
rect 21272 13744 21324 13753
rect 21640 13753 21652 13787
rect 21652 13753 21692 13787
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 27804 13880 27856 13932
rect 28632 13880 28684 13932
rect 27436 13855 27488 13864
rect 21640 13744 21692 13753
rect 23480 13744 23532 13796
rect 27436 13821 27445 13855
rect 27445 13821 27479 13855
rect 27479 13821 27488 13855
rect 27436 13812 27488 13821
rect 31300 14025 31309 14059
rect 31309 14025 31343 14059
rect 31343 14025 31352 14059
rect 31300 14016 31352 14025
rect 31484 14059 31536 14068
rect 31484 14025 31493 14059
rect 31493 14025 31527 14059
rect 31527 14025 31536 14059
rect 31484 14016 31536 14025
rect 32772 14016 32824 14068
rect 32956 14059 33008 14068
rect 32956 14025 32965 14059
rect 32965 14025 32999 14059
rect 32999 14025 33008 14059
rect 32956 14016 33008 14025
rect 31760 13948 31812 14000
rect 30380 13923 30432 13932
rect 30380 13889 30389 13923
rect 30389 13889 30423 13923
rect 30423 13889 30432 13923
rect 30380 13880 30432 13889
rect 30288 13855 30340 13864
rect 30288 13821 30297 13855
rect 30297 13821 30331 13855
rect 30331 13821 30340 13855
rect 30288 13812 30340 13821
rect 31116 13812 31168 13864
rect 31668 13855 31720 13864
rect 31668 13821 31677 13855
rect 31677 13821 31711 13855
rect 31711 13821 31720 13855
rect 31668 13812 31720 13821
rect 24124 13744 24176 13796
rect 23020 13676 23072 13728
rect 26240 13719 26292 13728
rect 26240 13685 26249 13719
rect 26249 13685 26283 13719
rect 26283 13685 26292 13719
rect 26240 13676 26292 13685
rect 29828 13676 29880 13728
rect 32588 13676 32640 13728
rect 34428 13676 34480 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 21640 13515 21692 13524
rect 21640 13481 21649 13515
rect 21649 13481 21683 13515
rect 21683 13481 21692 13515
rect 21640 13472 21692 13481
rect 22008 13472 22060 13524
rect 24124 13515 24176 13524
rect 24124 13481 24133 13515
rect 24133 13481 24167 13515
rect 24167 13481 24176 13515
rect 24124 13472 24176 13481
rect 24216 13472 24268 13524
rect 24860 13472 24912 13524
rect 27160 13515 27212 13524
rect 27160 13481 27169 13515
rect 27169 13481 27203 13515
rect 27203 13481 27212 13515
rect 27160 13472 27212 13481
rect 28632 13515 28684 13524
rect 28632 13481 28641 13515
rect 28641 13481 28675 13515
rect 28675 13481 28684 13515
rect 28632 13472 28684 13481
rect 29000 13515 29052 13524
rect 29000 13481 29009 13515
rect 29009 13481 29043 13515
rect 29043 13481 29052 13515
rect 29000 13472 29052 13481
rect 30288 13472 30340 13524
rect 31024 13472 31076 13524
rect 31760 13472 31812 13524
rect 32956 13472 33008 13524
rect 35808 13515 35860 13524
rect 35808 13481 35817 13515
rect 35817 13481 35851 13515
rect 35851 13481 35860 13515
rect 35808 13472 35860 13481
rect 26240 13404 26292 13456
rect 20904 13336 20956 13388
rect 23020 13379 23072 13388
rect 23020 13345 23054 13379
rect 23054 13345 23072 13379
rect 23020 13336 23072 13345
rect 25136 13336 25188 13388
rect 25320 13379 25372 13388
rect 25320 13345 25329 13379
rect 25329 13345 25363 13379
rect 25363 13345 25372 13379
rect 25320 13336 25372 13345
rect 28172 13336 28224 13388
rect 29828 13379 29880 13388
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 33692 13336 33744 13388
rect 36544 13336 36596 13388
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22100 13268 22152 13320
rect 21180 13175 21232 13184
rect 21180 13141 21189 13175
rect 21189 13141 21223 13175
rect 21223 13141 21232 13175
rect 21180 13132 21232 13141
rect 22192 13132 22244 13184
rect 25412 13268 25464 13320
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 27896 13311 27948 13320
rect 27896 13277 27905 13311
rect 27905 13277 27939 13311
rect 27939 13277 27948 13311
rect 27896 13268 27948 13277
rect 29184 13268 29236 13320
rect 29736 13268 29788 13320
rect 30012 13311 30064 13320
rect 30012 13277 30021 13311
rect 30021 13277 30055 13311
rect 30055 13277 30064 13311
rect 30012 13268 30064 13277
rect 33508 13268 33560 13320
rect 35716 13268 35768 13320
rect 36452 13311 36504 13320
rect 30656 13200 30708 13252
rect 31668 13200 31720 13252
rect 36452 13277 36461 13311
rect 36461 13277 36495 13311
rect 36495 13277 36504 13311
rect 36452 13268 36504 13277
rect 37556 13200 37608 13252
rect 27252 13132 27304 13184
rect 29460 13175 29512 13184
rect 29460 13141 29469 13175
rect 29469 13141 29503 13175
rect 29503 13141 29512 13175
rect 29460 13132 29512 13141
rect 34704 13132 34756 13184
rect 35348 13175 35400 13184
rect 35348 13141 35357 13175
rect 35357 13141 35391 13175
rect 35391 13141 35400 13175
rect 35348 13132 35400 13141
rect 36268 13132 36320 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 21732 12928 21784 12980
rect 22008 12928 22060 12980
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 23480 12928 23532 12980
rect 24768 12971 24820 12980
rect 24768 12937 24777 12971
rect 24777 12937 24811 12971
rect 24811 12937 24820 12971
rect 24768 12928 24820 12937
rect 25136 12971 25188 12980
rect 25136 12937 25145 12971
rect 25145 12937 25179 12971
rect 25179 12937 25188 12971
rect 25136 12928 25188 12937
rect 27436 12928 27488 12980
rect 27804 12971 27856 12980
rect 27804 12937 27813 12971
rect 27813 12937 27847 12971
rect 27847 12937 27856 12971
rect 27804 12928 27856 12937
rect 28172 12971 28224 12980
rect 28172 12937 28181 12971
rect 28181 12937 28215 12971
rect 28215 12937 28224 12971
rect 28172 12928 28224 12937
rect 29368 12928 29420 12980
rect 29828 12928 29880 12980
rect 29920 12928 29972 12980
rect 31024 12928 31076 12980
rect 34704 12971 34756 12980
rect 20904 12903 20956 12912
rect 20904 12869 20913 12903
rect 20913 12869 20947 12903
rect 20947 12869 20956 12903
rect 20904 12860 20956 12869
rect 21272 12903 21324 12912
rect 21272 12869 21281 12903
rect 21281 12869 21315 12903
rect 21315 12869 21324 12903
rect 21272 12860 21324 12869
rect 21364 12835 21416 12844
rect 21364 12801 21373 12835
rect 21373 12801 21407 12835
rect 21407 12801 21416 12835
rect 21364 12792 21416 12801
rect 24676 12792 24728 12844
rect 26148 12860 26200 12912
rect 24860 12792 24912 12844
rect 22192 12724 22244 12776
rect 23664 12724 23716 12776
rect 25228 12724 25280 12776
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 27528 12792 27580 12844
rect 27712 12792 27764 12844
rect 29460 12860 29512 12912
rect 29920 12767 29972 12776
rect 29920 12733 29929 12767
rect 29929 12733 29963 12767
rect 29963 12733 29972 12767
rect 29920 12724 29972 12733
rect 30288 12724 30340 12776
rect 33048 12860 33100 12912
rect 34704 12937 34713 12971
rect 34713 12937 34747 12971
rect 34747 12937 34756 12971
rect 34704 12928 34756 12937
rect 36452 12928 36504 12980
rect 36820 12928 36872 12980
rect 37556 12971 37608 12980
rect 37556 12937 37565 12971
rect 37565 12937 37599 12971
rect 37599 12937 37608 12971
rect 37556 12928 37608 12937
rect 33692 12792 33744 12844
rect 36544 12903 36596 12912
rect 36544 12869 36553 12903
rect 36553 12869 36587 12903
rect 36587 12869 36596 12903
rect 36544 12860 36596 12869
rect 33416 12724 33468 12776
rect 33508 12724 33560 12776
rect 21456 12656 21508 12708
rect 24216 12656 24268 12708
rect 25320 12656 25372 12708
rect 32956 12699 33008 12708
rect 32956 12665 32965 12699
rect 32965 12665 32999 12699
rect 32999 12665 33008 12699
rect 32956 12656 33008 12665
rect 35348 12656 35400 12708
rect 24032 12631 24084 12640
rect 24032 12597 24041 12631
rect 24041 12597 24075 12631
rect 24075 12597 24084 12631
rect 24032 12588 24084 12597
rect 25872 12588 25924 12640
rect 26976 12588 27028 12640
rect 31300 12588 31352 12640
rect 35992 12588 36044 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 21456 12427 21508 12436
rect 21456 12393 21465 12427
rect 21465 12393 21499 12427
rect 21499 12393 21508 12427
rect 21456 12384 21508 12393
rect 23848 12384 23900 12436
rect 24032 12427 24084 12436
rect 24032 12393 24041 12427
rect 24041 12393 24075 12427
rect 24075 12393 24084 12427
rect 24032 12384 24084 12393
rect 24216 12427 24268 12436
rect 24216 12393 24225 12427
rect 24225 12393 24259 12427
rect 24259 12393 24268 12427
rect 24216 12384 24268 12393
rect 25228 12427 25280 12436
rect 25228 12393 25237 12427
rect 25237 12393 25271 12427
rect 25271 12393 25280 12427
rect 25228 12384 25280 12393
rect 27712 12384 27764 12436
rect 29184 12427 29236 12436
rect 29184 12393 29193 12427
rect 29193 12393 29227 12427
rect 29227 12393 29236 12427
rect 29184 12384 29236 12393
rect 29552 12427 29604 12436
rect 29552 12393 29561 12427
rect 29561 12393 29595 12427
rect 29595 12393 29604 12427
rect 29552 12384 29604 12393
rect 30012 12384 30064 12436
rect 31116 12427 31168 12436
rect 31116 12393 31125 12427
rect 31125 12393 31159 12427
rect 31159 12393 31168 12427
rect 31116 12384 31168 12393
rect 34244 12384 34296 12436
rect 34704 12384 34756 12436
rect 36820 12427 36872 12436
rect 36820 12393 36829 12427
rect 36829 12393 36863 12427
rect 36863 12393 36872 12427
rect 36820 12384 36872 12393
rect 27344 12316 27396 12368
rect 27896 12316 27948 12368
rect 35992 12316 36044 12368
rect 22100 12248 22152 12300
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 27620 12291 27672 12300
rect 27620 12257 27654 12291
rect 27654 12257 27672 12291
rect 27620 12248 27672 12257
rect 30012 12291 30064 12300
rect 30012 12257 30046 12291
rect 30046 12257 30064 12291
rect 30012 12248 30064 12257
rect 32404 12248 32456 12300
rect 24492 12180 24544 12232
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 26700 12180 26752 12232
rect 24308 12112 24360 12164
rect 22192 12044 22244 12096
rect 26976 12044 27028 12096
rect 31024 12180 31076 12232
rect 31944 12180 31996 12232
rect 33232 12223 33284 12232
rect 33232 12189 33244 12223
rect 33244 12189 33278 12223
rect 33278 12189 33284 12223
rect 34244 12248 34296 12300
rect 33232 12180 33284 12189
rect 33416 12180 33468 12232
rect 34152 12180 34204 12232
rect 36268 12248 36320 12300
rect 35256 12180 35308 12232
rect 32036 12044 32088 12096
rect 32496 12087 32548 12096
rect 32496 12053 32505 12087
rect 32505 12053 32539 12087
rect 32539 12053 32548 12087
rect 32496 12044 32548 12053
rect 32588 12044 32640 12096
rect 34796 12044 34848 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 22100 11883 22152 11892
rect 22100 11849 22109 11883
rect 22109 11849 22143 11883
rect 22143 11849 22152 11883
rect 23388 11883 23440 11892
rect 22100 11840 22152 11849
rect 23388 11849 23397 11883
rect 23397 11849 23431 11883
rect 23431 11849 23440 11883
rect 23388 11840 23440 11849
rect 23664 11883 23716 11892
rect 23664 11849 23673 11883
rect 23673 11849 23707 11883
rect 23707 11849 23716 11883
rect 23664 11840 23716 11849
rect 24584 11840 24636 11892
rect 27620 11840 27672 11892
rect 29552 11840 29604 11892
rect 32404 11883 32456 11892
rect 32404 11849 32413 11883
rect 32413 11849 32447 11883
rect 32447 11849 32456 11883
rect 32404 11840 32456 11849
rect 32036 11772 32088 11824
rect 33508 11840 33560 11892
rect 33692 11840 33744 11892
rect 34152 11883 34204 11892
rect 34152 11849 34161 11883
rect 34161 11849 34195 11883
rect 34195 11849 34204 11883
rect 34152 11840 34204 11849
rect 35992 11883 36044 11892
rect 35992 11849 36001 11883
rect 36001 11849 36035 11883
rect 36035 11849 36044 11883
rect 35992 11840 36044 11849
rect 36268 11883 36320 11892
rect 36268 11849 36277 11883
rect 36277 11849 36311 11883
rect 36311 11849 36320 11883
rect 36268 11840 36320 11849
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 34796 11772 34848 11824
rect 23848 11636 23900 11688
rect 26700 11679 26752 11688
rect 26700 11645 26709 11679
rect 26709 11645 26743 11679
rect 26743 11645 26752 11679
rect 26700 11636 26752 11645
rect 29276 11679 29328 11688
rect 29276 11645 29285 11679
rect 29285 11645 29319 11679
rect 29319 11645 29328 11679
rect 29276 11636 29328 11645
rect 33968 11704 34020 11756
rect 34152 11704 34204 11756
rect 31116 11636 31168 11688
rect 33232 11636 33284 11688
rect 35256 11679 35308 11688
rect 35256 11645 35265 11679
rect 35265 11645 35299 11679
rect 35299 11645 35308 11679
rect 35256 11636 35308 11645
rect 36452 11679 36504 11688
rect 36452 11645 36461 11679
rect 36461 11645 36495 11679
rect 36495 11645 36504 11679
rect 36452 11636 36504 11645
rect 23388 11568 23440 11620
rect 26884 11568 26936 11620
rect 31668 11568 31720 11620
rect 32404 11568 32456 11620
rect 32496 11568 32548 11620
rect 22192 11500 22244 11552
rect 24492 11500 24544 11552
rect 24676 11543 24728 11552
rect 24676 11509 24685 11543
rect 24685 11509 24719 11543
rect 24719 11509 24728 11543
rect 24676 11500 24728 11509
rect 27620 11500 27672 11552
rect 30012 11500 30064 11552
rect 31760 11500 31812 11552
rect 35716 11568 35768 11620
rect 36636 11543 36688 11552
rect 36636 11509 36645 11543
rect 36645 11509 36679 11543
rect 36679 11509 36688 11543
rect 36636 11500 36688 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 23388 11296 23440 11348
rect 24308 11339 24360 11348
rect 24308 11305 24317 11339
rect 24317 11305 24351 11339
rect 24351 11305 24360 11339
rect 24308 11296 24360 11305
rect 24584 11296 24636 11348
rect 30380 11296 30432 11348
rect 31944 11339 31996 11348
rect 31944 11305 31953 11339
rect 31953 11305 31987 11339
rect 31987 11305 31996 11339
rect 31944 11296 31996 11305
rect 32496 11296 32548 11348
rect 34428 11296 34480 11348
rect 36452 11339 36504 11348
rect 36452 11305 36461 11339
rect 36461 11305 36495 11339
rect 36495 11305 36504 11339
rect 36452 11296 36504 11305
rect 24216 11228 24268 11280
rect 22284 11160 22336 11212
rect 24768 11203 24820 11212
rect 24768 11169 24777 11203
rect 24777 11169 24811 11203
rect 24811 11169 24820 11203
rect 24768 11160 24820 11169
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 27712 11228 27764 11280
rect 29552 11271 29604 11280
rect 29552 11237 29586 11271
rect 29586 11237 29604 11271
rect 29552 11228 29604 11237
rect 33140 11228 33192 11280
rect 36084 11271 36136 11280
rect 36084 11237 36093 11271
rect 36093 11237 36127 11271
rect 36127 11237 36136 11271
rect 36084 11228 36136 11237
rect 26700 11160 26752 11212
rect 32680 11160 32732 11212
rect 34612 11160 34664 11212
rect 25044 10956 25096 11008
rect 28724 11092 28776 11144
rect 29276 11135 29328 11144
rect 29276 11101 29285 11135
rect 29285 11101 29319 11135
rect 29319 11101 29328 11135
rect 29276 11092 29328 11101
rect 31484 11092 31536 11144
rect 36176 11160 36228 11212
rect 25412 10956 25464 11008
rect 26884 10956 26936 11008
rect 27436 10956 27488 11008
rect 34520 11067 34572 11076
rect 34520 11033 34529 11067
rect 34529 11033 34563 11067
rect 34563 11033 34572 11067
rect 34520 11024 34572 11033
rect 35992 10956 36044 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 22284 10795 22336 10804
rect 22284 10761 22293 10795
rect 22293 10761 22327 10795
rect 22327 10761 22336 10795
rect 22284 10752 22336 10761
rect 25412 10795 25464 10804
rect 25412 10761 25421 10795
rect 25421 10761 25455 10795
rect 25455 10761 25464 10795
rect 25412 10752 25464 10761
rect 27344 10752 27396 10804
rect 27712 10752 27764 10804
rect 29552 10752 29604 10804
rect 31760 10795 31812 10804
rect 31760 10761 31769 10795
rect 31769 10761 31803 10795
rect 31803 10761 31812 10795
rect 31760 10752 31812 10761
rect 32956 10752 33008 10804
rect 34428 10752 34480 10804
rect 29368 10616 29420 10668
rect 32496 10659 32548 10668
rect 32496 10625 32505 10659
rect 32505 10625 32539 10659
rect 32539 10625 32548 10659
rect 32496 10616 32548 10625
rect 33048 10659 33100 10668
rect 33048 10625 33057 10659
rect 33057 10625 33091 10659
rect 33091 10625 33100 10659
rect 33048 10616 33100 10625
rect 22192 10548 22244 10600
rect 22744 10548 22796 10600
rect 23756 10548 23808 10600
rect 25872 10591 25924 10600
rect 25872 10557 25881 10591
rect 25881 10557 25915 10591
rect 25915 10557 25924 10591
rect 25872 10548 25924 10557
rect 30656 10591 30708 10600
rect 30656 10557 30665 10591
rect 30665 10557 30699 10591
rect 30699 10557 30708 10591
rect 30656 10548 30708 10557
rect 24492 10480 24544 10532
rect 26148 10523 26200 10532
rect 26148 10489 26182 10523
rect 26182 10489 26200 10523
rect 26148 10480 26200 10489
rect 27528 10480 27580 10532
rect 31208 10548 31260 10600
rect 31760 10548 31812 10600
rect 33140 10548 33192 10600
rect 35992 10548 36044 10600
rect 32680 10480 32732 10532
rect 33416 10523 33468 10532
rect 33416 10489 33425 10523
rect 33425 10489 33459 10523
rect 33459 10489 33468 10523
rect 33416 10480 33468 10489
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 27252 10455 27304 10464
rect 27252 10421 27261 10455
rect 27261 10421 27295 10455
rect 27295 10421 27304 10455
rect 27252 10412 27304 10421
rect 28724 10412 28776 10464
rect 30840 10412 30892 10464
rect 31024 10455 31076 10464
rect 31024 10421 31033 10455
rect 31033 10421 31067 10455
rect 31067 10421 31076 10455
rect 31024 10412 31076 10421
rect 32404 10455 32456 10464
rect 32404 10421 32413 10455
rect 32413 10421 32447 10455
rect 32447 10421 32456 10455
rect 33692 10455 33744 10464
rect 32404 10412 32456 10421
rect 33692 10421 33701 10455
rect 33701 10421 33735 10455
rect 33735 10421 33744 10455
rect 33692 10412 33744 10421
rect 36176 10480 36228 10532
rect 37096 10455 37148 10464
rect 37096 10421 37105 10455
rect 37105 10421 37139 10455
rect 37139 10421 37148 10455
rect 37096 10412 37148 10421
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 22284 10208 22336 10260
rect 24768 10251 24820 10260
rect 24768 10217 24777 10251
rect 24777 10217 24811 10251
rect 24811 10217 24820 10251
rect 24768 10208 24820 10217
rect 26976 10251 27028 10260
rect 26976 10217 26985 10251
rect 26985 10217 27019 10251
rect 27019 10217 27028 10251
rect 26976 10208 27028 10217
rect 27528 10208 27580 10260
rect 30656 10208 30708 10260
rect 30840 10208 30892 10260
rect 31484 10251 31536 10260
rect 31484 10217 31493 10251
rect 31493 10217 31527 10251
rect 31527 10217 31536 10251
rect 31484 10208 31536 10217
rect 32404 10251 32456 10260
rect 32404 10217 32413 10251
rect 32413 10217 32447 10251
rect 32447 10217 32456 10251
rect 32404 10208 32456 10217
rect 32588 10208 32640 10260
rect 33692 10208 33744 10260
rect 34244 10208 34296 10260
rect 34612 10251 34664 10260
rect 34612 10217 34621 10251
rect 34621 10217 34655 10251
rect 34655 10217 34664 10251
rect 34612 10208 34664 10217
rect 35532 10208 35584 10260
rect 35716 10208 35768 10260
rect 36084 10251 36136 10260
rect 36084 10217 36093 10251
rect 36093 10217 36127 10251
rect 36127 10217 36136 10251
rect 36084 10208 36136 10217
rect 31024 10140 31076 10192
rect 32496 10140 32548 10192
rect 35624 10140 35676 10192
rect 22744 10115 22796 10124
rect 22744 10081 22753 10115
rect 22753 10081 22787 10115
rect 22787 10081 22796 10115
rect 22744 10072 22796 10081
rect 22836 10072 22888 10124
rect 25044 10072 25096 10124
rect 27344 10072 27396 10124
rect 27436 10047 27488 10056
rect 27436 10013 27445 10047
rect 27445 10013 27479 10047
rect 27479 10013 27488 10047
rect 27436 10004 27488 10013
rect 33968 10115 34020 10124
rect 33968 10081 33977 10115
rect 33977 10081 34011 10115
rect 34011 10081 34020 10115
rect 33968 10072 34020 10081
rect 34612 10072 34664 10124
rect 36268 10072 36320 10124
rect 36544 10115 36596 10124
rect 36544 10081 36553 10115
rect 36553 10081 36587 10115
rect 36587 10081 36596 10115
rect 36544 10072 36596 10081
rect 27620 10004 27672 10056
rect 33416 10004 33468 10056
rect 35532 9936 35584 9988
rect 25320 9868 25372 9920
rect 25872 9911 25924 9920
rect 25872 9877 25881 9911
rect 25881 9877 25915 9911
rect 25915 9877 25924 9911
rect 25872 9868 25924 9877
rect 31116 9911 31168 9920
rect 31116 9877 31125 9911
rect 31125 9877 31159 9911
rect 31159 9877 31168 9911
rect 31116 9868 31168 9877
rect 35900 9868 35952 9920
rect 36728 9911 36780 9920
rect 36728 9877 36737 9911
rect 36737 9877 36771 9911
rect 36771 9877 36780 9911
rect 36728 9868 36780 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 22836 9707 22888 9716
rect 22836 9673 22845 9707
rect 22845 9673 22879 9707
rect 22879 9673 22888 9707
rect 22836 9664 22888 9673
rect 26148 9707 26200 9716
rect 26148 9673 26157 9707
rect 26157 9673 26191 9707
rect 26191 9673 26200 9707
rect 26148 9664 26200 9673
rect 27436 9664 27488 9716
rect 32496 9707 32548 9716
rect 32496 9673 32505 9707
rect 32505 9673 32539 9707
rect 32539 9673 32548 9707
rect 32496 9664 32548 9673
rect 33968 9707 34020 9716
rect 33968 9673 33977 9707
rect 33977 9673 34011 9707
rect 34011 9673 34020 9707
rect 33968 9664 34020 9673
rect 22744 9596 22796 9648
rect 27620 9596 27672 9648
rect 28264 9528 28316 9580
rect 32588 9596 32640 9648
rect 33048 9596 33100 9648
rect 33876 9596 33928 9648
rect 34152 9664 34204 9716
rect 34612 9664 34664 9716
rect 35256 9664 35308 9716
rect 34520 9596 34572 9648
rect 23756 9503 23808 9512
rect 23756 9469 23765 9503
rect 23765 9469 23799 9503
rect 23799 9469 23808 9503
rect 23756 9460 23808 9469
rect 27620 9460 27672 9512
rect 31116 9460 31168 9512
rect 32956 9528 33008 9580
rect 34612 9528 34664 9580
rect 35900 9664 35952 9716
rect 36544 9707 36596 9716
rect 36544 9673 36553 9707
rect 36553 9673 36587 9707
rect 36587 9673 36596 9707
rect 36544 9664 36596 9673
rect 36268 9639 36320 9648
rect 36268 9605 36277 9639
rect 36277 9605 36311 9639
rect 36311 9605 36320 9639
rect 36268 9596 36320 9605
rect 37188 9596 37240 9648
rect 33232 9503 33284 9512
rect 33232 9469 33241 9503
rect 33241 9469 33275 9503
rect 33275 9469 33284 9503
rect 33232 9460 33284 9469
rect 33968 9460 34020 9512
rect 24584 9392 24636 9444
rect 26700 9392 26752 9444
rect 31576 9392 31628 9444
rect 35256 9392 35308 9444
rect 24492 9324 24544 9376
rect 27344 9367 27396 9376
rect 27344 9333 27353 9367
rect 27353 9333 27387 9367
rect 27387 9333 27396 9367
rect 27344 9324 27396 9333
rect 27436 9324 27488 9376
rect 31208 9324 31260 9376
rect 32956 9324 33008 9376
rect 34612 9367 34664 9376
rect 34612 9333 34621 9367
rect 34621 9333 34655 9367
rect 34655 9333 34664 9367
rect 34612 9324 34664 9333
rect 35532 9367 35584 9376
rect 35532 9333 35541 9367
rect 35541 9333 35575 9367
rect 35575 9333 35584 9367
rect 35532 9324 35584 9333
rect 36912 9367 36964 9376
rect 36912 9333 36921 9367
rect 36921 9333 36955 9367
rect 36955 9333 36964 9367
rect 36912 9324 36964 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 24676 9120 24728 9172
rect 27436 9163 27488 9172
rect 27436 9129 27445 9163
rect 27445 9129 27479 9163
rect 27479 9129 27488 9163
rect 27436 9120 27488 9129
rect 31116 9120 31168 9172
rect 31208 9120 31260 9172
rect 33232 9163 33284 9172
rect 33232 9129 33241 9163
rect 33241 9129 33275 9163
rect 33275 9129 33284 9163
rect 33232 9120 33284 9129
rect 34336 9163 34388 9172
rect 34336 9129 34345 9163
rect 34345 9129 34379 9163
rect 34379 9129 34388 9163
rect 34336 9120 34388 9129
rect 37096 9120 37148 9172
rect 24492 9095 24544 9104
rect 24492 9061 24501 9095
rect 24501 9061 24535 9095
rect 24535 9061 24544 9095
rect 24492 9052 24544 9061
rect 24584 9095 24636 9104
rect 24584 9061 24593 9095
rect 24593 9061 24627 9095
rect 24627 9061 24636 9095
rect 24584 9052 24636 9061
rect 32680 9052 32732 9104
rect 32956 9095 33008 9104
rect 32956 9061 32965 9095
rect 32965 9061 32999 9095
rect 32999 9061 33008 9095
rect 32956 9052 33008 9061
rect 23756 8984 23808 9036
rect 25320 8984 25372 9036
rect 27160 8984 27212 9036
rect 28816 8984 28868 9036
rect 29644 9027 29696 9036
rect 29644 8993 29653 9027
rect 29653 8993 29687 9027
rect 29687 8993 29696 9027
rect 29644 8984 29696 8993
rect 24216 8916 24268 8968
rect 28172 8959 28224 8968
rect 28172 8925 28181 8959
rect 28181 8925 28215 8959
rect 28215 8925 28224 8959
rect 28172 8916 28224 8925
rect 28264 8959 28316 8968
rect 28264 8925 28273 8959
rect 28273 8925 28307 8959
rect 28307 8925 28316 8959
rect 28264 8916 28316 8925
rect 29000 8916 29052 8968
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 29920 8959 29972 8968
rect 29920 8925 29929 8959
rect 29929 8925 29963 8959
rect 29963 8925 29972 8959
rect 29920 8916 29972 8925
rect 32036 8984 32088 9036
rect 33324 8984 33376 9036
rect 35992 9052 36044 9104
rect 35532 8984 35584 9036
rect 36820 8984 36872 9036
rect 33692 8959 33744 8968
rect 33692 8925 33701 8959
rect 33701 8925 33735 8959
rect 33735 8925 33744 8959
rect 33692 8916 33744 8925
rect 34336 8916 34388 8968
rect 30840 8848 30892 8900
rect 27712 8823 27764 8832
rect 27712 8789 27721 8823
rect 27721 8789 27755 8823
rect 27755 8789 27764 8823
rect 27712 8780 27764 8789
rect 28264 8780 28316 8832
rect 29920 8780 29972 8832
rect 30288 8823 30340 8832
rect 30288 8789 30297 8823
rect 30297 8789 30331 8823
rect 30331 8789 30340 8823
rect 30288 8780 30340 8789
rect 32312 8823 32364 8832
rect 32312 8789 32321 8823
rect 32321 8789 32355 8823
rect 32355 8789 32364 8823
rect 32312 8780 32364 8789
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 24492 8619 24544 8628
rect 24492 8585 24501 8619
rect 24501 8585 24535 8619
rect 24535 8585 24544 8619
rect 24492 8576 24544 8585
rect 26700 8619 26752 8628
rect 26700 8585 26709 8619
rect 26709 8585 26743 8619
rect 26743 8585 26752 8619
rect 26700 8576 26752 8585
rect 27160 8619 27212 8628
rect 27160 8585 27169 8619
rect 27169 8585 27203 8619
rect 27203 8585 27212 8619
rect 27160 8576 27212 8585
rect 28172 8576 28224 8628
rect 29644 8619 29696 8628
rect 29644 8585 29653 8619
rect 29653 8585 29687 8619
rect 29687 8585 29696 8619
rect 29644 8576 29696 8585
rect 29736 8576 29788 8628
rect 32312 8576 32364 8628
rect 33692 8576 33744 8628
rect 35440 8576 35492 8628
rect 36820 8619 36872 8628
rect 36820 8585 36829 8619
rect 36829 8585 36863 8619
rect 36863 8585 36872 8619
rect 36820 8576 36872 8585
rect 24400 8508 24452 8560
rect 27620 8551 27672 8560
rect 24584 8440 24636 8492
rect 27620 8517 27629 8551
rect 27629 8517 27663 8551
rect 27663 8517 27672 8551
rect 27620 8508 27672 8517
rect 25320 8415 25372 8424
rect 25320 8381 25329 8415
rect 25329 8381 25363 8415
rect 25363 8381 25372 8415
rect 25320 8372 25372 8381
rect 27344 8440 27396 8492
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 28356 8440 28408 8492
rect 30288 8440 30340 8492
rect 31852 8440 31904 8492
rect 32588 8483 32640 8492
rect 32588 8449 32597 8483
rect 32597 8449 32631 8483
rect 32631 8449 32640 8483
rect 32588 8440 32640 8449
rect 33784 8508 33836 8560
rect 34612 8508 34664 8560
rect 27712 8372 27764 8424
rect 30288 8304 30340 8356
rect 32772 8372 32824 8424
rect 33692 8415 33744 8424
rect 33692 8381 33701 8415
rect 33701 8381 33735 8415
rect 33735 8381 33744 8415
rect 33692 8372 33744 8381
rect 35440 8415 35492 8424
rect 35440 8381 35449 8415
rect 35449 8381 35483 8415
rect 35483 8381 35492 8415
rect 35440 8372 35492 8381
rect 35992 8372 36044 8424
rect 32036 8304 32088 8356
rect 35256 8304 35308 8356
rect 30380 8236 30432 8288
rect 32128 8279 32180 8288
rect 32128 8245 32137 8279
rect 32137 8245 32171 8279
rect 32171 8245 32180 8279
rect 32128 8236 32180 8245
rect 33324 8236 33376 8288
rect 36636 8236 36688 8288
rect 37096 8279 37148 8288
rect 37096 8245 37105 8279
rect 37105 8245 37139 8279
rect 37139 8245 37148 8279
rect 37096 8236 37148 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 24216 8075 24268 8084
rect 24216 8041 24225 8075
rect 24225 8041 24259 8075
rect 24259 8041 24268 8075
rect 24216 8032 24268 8041
rect 27712 8032 27764 8084
rect 28356 8032 28408 8084
rect 30840 8075 30892 8084
rect 30840 8041 30849 8075
rect 30849 8041 30883 8075
rect 30883 8041 30892 8075
rect 30840 8032 30892 8041
rect 31852 8075 31904 8084
rect 31852 8041 31861 8075
rect 31861 8041 31895 8075
rect 31895 8041 31904 8075
rect 31852 8032 31904 8041
rect 32128 8032 32180 8084
rect 33324 8075 33376 8084
rect 33324 8041 33333 8075
rect 33333 8041 33367 8075
rect 33367 8041 33376 8075
rect 33324 8032 33376 8041
rect 33692 8075 33744 8084
rect 33692 8041 33701 8075
rect 33701 8041 33735 8075
rect 33735 8041 33744 8075
rect 33692 8032 33744 8041
rect 34428 8032 34480 8084
rect 36636 8075 36688 8084
rect 36636 8041 36645 8075
rect 36645 8041 36679 8075
rect 36679 8041 36688 8075
rect 36636 8032 36688 8041
rect 26700 7964 26752 8016
rect 29000 7939 29052 7948
rect 29000 7905 29034 7939
rect 29034 7905 29052 7939
rect 29000 7896 29052 7905
rect 32496 7939 32548 7948
rect 32496 7905 32505 7939
rect 32505 7905 32539 7939
rect 32539 7905 32548 7939
rect 32496 7896 32548 7905
rect 35440 7964 35492 8016
rect 36544 7896 36596 7948
rect 25320 7828 25372 7880
rect 26240 7828 26292 7880
rect 28724 7871 28776 7880
rect 28724 7837 28733 7871
rect 28733 7837 28767 7871
rect 28767 7837 28776 7871
rect 28724 7828 28776 7837
rect 31944 7828 31996 7880
rect 34152 7871 34204 7880
rect 32036 7760 32088 7812
rect 34152 7837 34161 7871
rect 34161 7837 34195 7871
rect 34195 7837 34204 7871
rect 34152 7828 34204 7837
rect 34336 7871 34388 7880
rect 34336 7837 34345 7871
rect 34345 7837 34379 7871
rect 34379 7837 34388 7871
rect 34336 7828 34388 7837
rect 27436 7692 27488 7744
rect 30104 7735 30156 7744
rect 30104 7701 30113 7735
rect 30113 7701 30147 7735
rect 30147 7701 30156 7735
rect 30104 7692 30156 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 26240 7531 26292 7540
rect 26240 7497 26249 7531
rect 26249 7497 26283 7531
rect 26283 7497 26292 7531
rect 26240 7488 26292 7497
rect 26700 7488 26752 7540
rect 28172 7488 28224 7540
rect 29000 7488 29052 7540
rect 32496 7488 32548 7540
rect 33232 7488 33284 7540
rect 34428 7488 34480 7540
rect 37096 7488 37148 7540
rect 30380 7420 30432 7472
rect 30932 7420 30984 7472
rect 28816 7352 28868 7404
rect 27436 7284 27488 7336
rect 28724 7284 28776 7336
rect 29276 7327 29328 7336
rect 29276 7293 29285 7327
rect 29285 7293 29319 7327
rect 29319 7293 29328 7327
rect 29276 7284 29328 7293
rect 27252 7216 27304 7268
rect 32588 7420 32640 7472
rect 31484 7327 31536 7336
rect 31484 7293 31493 7327
rect 31493 7293 31527 7327
rect 31527 7293 31536 7327
rect 31484 7284 31536 7293
rect 34888 7327 34940 7336
rect 34888 7293 34897 7327
rect 34897 7293 34931 7327
rect 34931 7293 34940 7327
rect 34888 7284 34940 7293
rect 35440 7284 35492 7336
rect 34152 7148 34204 7200
rect 34428 7148 34480 7200
rect 34612 7191 34664 7200
rect 34612 7157 34621 7191
rect 34621 7157 34655 7191
rect 34655 7157 34664 7191
rect 34612 7148 34664 7157
rect 35900 7148 35952 7200
rect 36544 7191 36596 7200
rect 36544 7157 36553 7191
rect 36553 7157 36587 7191
rect 36587 7157 36596 7191
rect 36544 7148 36596 7157
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 27436 6944 27488 6996
rect 31944 6987 31996 6996
rect 31944 6953 31953 6987
rect 31953 6953 31987 6987
rect 31987 6953 31996 6987
rect 31944 6944 31996 6953
rect 32128 6944 32180 6996
rect 34336 6944 34388 6996
rect 34612 6944 34664 6996
rect 27344 6808 27396 6860
rect 28172 6876 28224 6928
rect 29092 6876 29144 6928
rect 30104 6876 30156 6928
rect 29276 6808 29328 6860
rect 29552 6808 29604 6860
rect 32772 6851 32824 6860
rect 32772 6817 32806 6851
rect 32806 6817 32824 6851
rect 32772 6808 32824 6817
rect 35072 6876 35124 6928
rect 27252 6783 27304 6792
rect 27252 6749 27261 6783
rect 27261 6749 27295 6783
rect 27295 6749 27304 6783
rect 27252 6740 27304 6749
rect 31484 6740 31536 6792
rect 32496 6783 32548 6792
rect 32496 6749 32505 6783
rect 32505 6749 32539 6783
rect 32539 6749 32548 6783
rect 32496 6740 32548 6749
rect 28816 6672 28868 6724
rect 30380 6604 30432 6656
rect 33692 6604 33744 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 27344 6443 27396 6452
rect 27344 6409 27353 6443
rect 27353 6409 27387 6443
rect 27387 6409 27396 6443
rect 27344 6400 27396 6409
rect 29092 6443 29144 6452
rect 29092 6409 29101 6443
rect 29101 6409 29135 6443
rect 29135 6409 29144 6443
rect 29092 6400 29144 6409
rect 30932 6443 30984 6452
rect 30932 6409 30941 6443
rect 30941 6409 30975 6443
rect 30975 6409 30984 6443
rect 30932 6400 30984 6409
rect 32772 6400 32824 6452
rect 36544 6400 36596 6452
rect 37096 6400 37148 6452
rect 27252 6196 27304 6248
rect 29552 6239 29604 6248
rect 29552 6205 29561 6239
rect 29561 6205 29595 6239
rect 29595 6205 29604 6239
rect 29552 6196 29604 6205
rect 29828 6239 29880 6248
rect 29828 6205 29862 6239
rect 29862 6205 29880 6239
rect 29828 6196 29880 6205
rect 30380 6196 30432 6248
rect 31760 6239 31812 6248
rect 31760 6205 31769 6239
rect 31769 6205 31803 6239
rect 31803 6205 31812 6239
rect 31760 6196 31812 6205
rect 32588 6196 32640 6248
rect 34796 6196 34848 6248
rect 35440 6196 35492 6248
rect 35900 6196 35952 6248
rect 33692 6060 33744 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 28908 5856 28960 5908
rect 29092 5856 29144 5908
rect 29828 5899 29880 5908
rect 29828 5865 29837 5899
rect 29837 5865 29871 5899
rect 29871 5865 29880 5899
rect 29828 5856 29880 5865
rect 32772 5856 32824 5908
rect 33232 5899 33284 5908
rect 33232 5865 33241 5899
rect 33241 5865 33275 5899
rect 33275 5865 33284 5899
rect 33232 5856 33284 5865
rect 34520 5856 34572 5908
rect 35532 5856 35584 5908
rect 36544 5856 36596 5908
rect 29000 5788 29052 5840
rect 29552 5788 29604 5840
rect 31760 5788 31812 5840
rect 32496 5788 32548 5840
rect 34796 5831 34848 5840
rect 34796 5797 34805 5831
rect 34805 5797 34839 5831
rect 34839 5797 34848 5831
rect 34796 5788 34848 5797
rect 35440 5788 35492 5840
rect 33600 5763 33652 5772
rect 33600 5729 33609 5763
rect 33609 5729 33643 5763
rect 33643 5729 33652 5763
rect 33600 5720 33652 5729
rect 34612 5720 34664 5772
rect 28356 5652 28408 5704
rect 33692 5695 33744 5704
rect 33692 5661 33701 5695
rect 33701 5661 33735 5695
rect 33735 5661 33744 5695
rect 33692 5652 33744 5661
rect 33784 5695 33836 5704
rect 33784 5661 33793 5695
rect 33793 5661 33827 5695
rect 33827 5661 33836 5695
rect 33784 5652 33836 5661
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 28356 5312 28408 5364
rect 28908 5355 28960 5364
rect 28908 5321 28917 5355
rect 28917 5321 28951 5355
rect 28951 5321 28960 5355
rect 28908 5312 28960 5321
rect 29092 5312 29144 5364
rect 33692 5312 33744 5364
rect 33784 5312 33836 5364
rect 35532 5355 35584 5364
rect 35532 5321 35541 5355
rect 35541 5321 35575 5355
rect 35575 5321 35584 5355
rect 35532 5312 35584 5321
rect 33600 5287 33652 5296
rect 33600 5253 33609 5287
rect 33609 5253 33643 5287
rect 33643 5253 33652 5287
rect 33600 5244 33652 5253
rect 35440 5244 35492 5296
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 33876 2635 33928 2644
rect 33876 2601 33885 2635
rect 33885 2601 33919 2635
rect 33919 2601 33928 2635
rect 33876 2592 33928 2601
rect 36636 2456 36688 2508
rect 33508 2363 33560 2372
rect 33508 2329 33517 2363
rect 33517 2329 33551 2363
rect 33551 2329 33560 2363
rect 33508 2320 33560 2329
rect 9956 2252 10008 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
<< metal2 >>
rect 570 39520 626 40000
rect 1674 39520 1730 40000
rect 2778 39520 2834 40000
rect 3882 39520 3938 40000
rect 4986 39520 5042 40000
rect 6090 39520 6146 40000
rect 7194 39520 7250 40000
rect 8298 39520 8354 40000
rect 9402 39520 9458 40000
rect 10506 39520 10562 40000
rect 11610 39520 11666 40000
rect 12714 39520 12770 40000
rect 13910 39520 13966 40000
rect 15014 39520 15070 40000
rect 16118 39520 16174 40000
rect 17222 39520 17278 40000
rect 18326 39520 18382 40000
rect 19430 39520 19486 40000
rect 20534 39520 20590 40000
rect 21638 39520 21694 40000
rect 22742 39520 22798 40000
rect 23846 39520 23902 40000
rect 24950 39520 25006 40000
rect 26054 39520 26110 40000
rect 27250 39520 27306 40000
rect 28354 39520 28410 40000
rect 29458 39520 29514 40000
rect 30562 39520 30618 40000
rect 31666 39520 31722 40000
rect 32770 39520 32826 40000
rect 33874 39520 33930 40000
rect 34978 39520 35034 40000
rect 36082 39520 36138 40000
rect 37186 39520 37242 40000
rect 38290 39520 38346 40000
rect 39394 39520 39450 40000
rect 584 34746 612 39520
rect 1688 35290 1716 39520
rect 1676 35284 1728 35290
rect 1676 35226 1728 35232
rect 2042 35184 2098 35193
rect 1400 35148 1452 35154
rect 2042 35119 2098 35128
rect 1400 35090 1452 35096
rect 572 34740 624 34746
rect 572 34682 624 34688
rect 1412 34134 1440 35090
rect 2056 34746 2084 35119
rect 2044 34740 2096 34746
rect 2044 34682 2096 34688
rect 2056 34542 2084 34682
rect 2688 34672 2740 34678
rect 2792 34626 2820 39520
rect 3896 34746 3924 39520
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4710 35456 4766 35465
rect 4710 35391 4766 35400
rect 4724 35154 4752 35391
rect 5000 35290 5028 39520
rect 6104 35834 6132 39520
rect 7208 36922 7236 39520
rect 7196 36916 7248 36922
rect 7196 36858 7248 36864
rect 7472 36576 7524 36582
rect 7470 36544 7472 36553
rect 7524 36544 7526 36553
rect 7470 36479 7526 36488
rect 6828 36236 6880 36242
rect 6828 36178 6880 36184
rect 6840 35834 6868 36178
rect 7380 36032 7432 36038
rect 7380 35974 7432 35980
rect 6092 35828 6144 35834
rect 6092 35770 6144 35776
rect 6828 35828 6880 35834
rect 6828 35770 6880 35776
rect 7102 35728 7158 35737
rect 7102 35663 7158 35672
rect 7116 35630 7144 35663
rect 7104 35624 7156 35630
rect 7104 35566 7156 35572
rect 6092 35488 6144 35494
rect 6092 35430 6144 35436
rect 6104 35329 6132 35430
rect 6090 35320 6146 35329
rect 4988 35284 5040 35290
rect 7116 35290 7144 35566
rect 7288 35488 7340 35494
rect 7288 35430 7340 35436
rect 6090 35255 6146 35264
rect 7104 35284 7156 35290
rect 4988 35226 5040 35232
rect 7104 35226 7156 35232
rect 4712 35148 4764 35154
rect 4712 35090 4764 35096
rect 5172 35148 5224 35154
rect 5172 35090 5224 35096
rect 4618 35048 4674 35057
rect 4618 34983 4674 34992
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4632 34746 4660 34983
rect 3884 34740 3936 34746
rect 3884 34682 3936 34688
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 2740 34620 2820 34626
rect 2688 34614 2820 34620
rect 2700 34598 2820 34614
rect 3146 34640 3202 34649
rect 4724 34610 4752 35090
rect 3146 34575 3148 34584
rect 3200 34575 3202 34584
rect 4712 34604 4764 34610
rect 3148 34546 3200 34552
rect 4712 34546 4764 34552
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 5184 34406 5212 35090
rect 5908 34944 5960 34950
rect 5908 34886 5960 34892
rect 6644 34944 6696 34950
rect 6644 34886 6696 34892
rect 5448 34672 5500 34678
rect 5448 34614 5500 34620
rect 5172 34400 5224 34406
rect 5172 34342 5224 34348
rect 1400 34128 1452 34134
rect 2872 34128 2924 34134
rect 1400 34070 1452 34076
rect 2870 34096 2872 34105
rect 2924 34096 2926 34105
rect 5184 34066 5212 34342
rect 2870 34031 2926 34040
rect 5172 34060 5224 34066
rect 5172 34002 5224 34008
rect 4712 33992 4764 33998
rect 4712 33934 4764 33940
rect 3516 33924 3568 33930
rect 3516 33866 3568 33872
rect 2964 33856 3016 33862
rect 2964 33798 3016 33804
rect 2976 33454 3004 33798
rect 3528 33522 3556 33866
rect 4068 33856 4120 33862
rect 4068 33798 4120 33804
rect 3516 33516 3568 33522
rect 3516 33458 3568 33464
rect 4080 33454 4108 33798
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 2964 33448 3016 33454
rect 2964 33390 3016 33396
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 1768 33312 1820 33318
rect 1768 33254 1820 33260
rect 2872 33312 2924 33318
rect 2872 33254 2924 33260
rect 1780 32910 1808 33254
rect 2884 33114 2912 33254
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 1860 32972 1912 32978
rect 1860 32914 1912 32920
rect 1768 32904 1820 32910
rect 1768 32846 1820 32852
rect 1400 32768 1452 32774
rect 1400 32710 1452 32716
rect 1412 32366 1440 32710
rect 1872 32570 1900 32914
rect 2976 32842 3004 33390
rect 3332 33312 3384 33318
rect 3332 33254 3384 33260
rect 3344 32978 3372 33254
rect 3792 33108 3844 33114
rect 3792 33050 3844 33056
rect 3332 32972 3384 32978
rect 3332 32914 3384 32920
rect 2964 32836 3016 32842
rect 2964 32778 3016 32784
rect 1860 32564 1912 32570
rect 1860 32506 1912 32512
rect 2976 32502 3004 32778
rect 3344 32570 3372 32914
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 3700 32768 3752 32774
rect 3700 32710 3752 32716
rect 3332 32564 3384 32570
rect 3332 32506 3384 32512
rect 2964 32496 3016 32502
rect 2964 32438 3016 32444
rect 3528 32434 3556 32710
rect 3516 32428 3568 32434
rect 3516 32370 3568 32376
rect 3712 32366 3740 32710
rect 3804 32366 3832 33050
rect 4080 32910 4108 33390
rect 4724 33386 4752 33934
rect 4712 33380 4764 33386
rect 4712 33322 4764 33328
rect 4724 33114 4752 33322
rect 4712 33108 4764 33114
rect 4712 33050 4764 33056
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 5460 32552 5488 34614
rect 5920 34542 5948 34886
rect 6092 34604 6144 34610
rect 6092 34546 6144 34552
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5632 34400 5684 34406
rect 5632 34342 5684 34348
rect 5644 34202 5672 34342
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 5724 34196 5776 34202
rect 5724 34138 5776 34144
rect 5540 33992 5592 33998
rect 5540 33934 5592 33940
rect 5552 33114 5580 33934
rect 5540 33108 5592 33114
rect 5540 33050 5592 33056
rect 5552 32722 5580 33050
rect 5552 32694 5672 32722
rect 5540 32564 5592 32570
rect 5460 32524 5540 32552
rect 5540 32506 5592 32512
rect 3976 32428 4028 32434
rect 3976 32370 4028 32376
rect 5172 32428 5224 32434
rect 5172 32370 5224 32376
rect 1400 32360 1452 32366
rect 1400 32302 1452 32308
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3792 32360 3844 32366
rect 3792 32302 3844 32308
rect 1412 31822 1440 32302
rect 2780 32292 2832 32298
rect 2780 32234 2832 32240
rect 2792 32026 2820 32234
rect 3252 32026 3280 32302
rect 3700 32224 3752 32230
rect 3700 32166 3752 32172
rect 2780 32020 2832 32026
rect 2780 31962 2832 31968
rect 3240 32020 3292 32026
rect 3240 31962 3292 31968
rect 3712 31958 3740 32166
rect 3424 31952 3476 31958
rect 3424 31894 3476 31900
rect 3700 31952 3752 31958
rect 3700 31894 3752 31900
rect 2504 31884 2556 31890
rect 2504 31826 2556 31832
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31346 1440 31758
rect 2516 31414 2544 31826
rect 3436 31482 3464 31894
rect 3700 31680 3752 31686
rect 3700 31622 3752 31628
rect 3424 31476 3476 31482
rect 3424 31418 3476 31424
rect 2504 31408 2556 31414
rect 2504 31350 2556 31356
rect 1400 31340 1452 31346
rect 1400 31282 1452 31288
rect 1412 30870 1440 31282
rect 1676 31204 1728 31210
rect 1676 31146 1728 31152
rect 1400 30864 1452 30870
rect 1400 30806 1452 30812
rect 1412 30394 1440 30806
rect 1688 30705 1716 31146
rect 2516 30938 2544 31350
rect 3712 31210 3740 31622
rect 3988 31346 4016 32370
rect 4068 32224 4120 32230
rect 4068 32166 4120 32172
rect 4528 32224 4580 32230
rect 4528 32166 4580 32172
rect 4080 31929 4108 32166
rect 4540 32026 4568 32166
rect 5184 32026 5212 32370
rect 5552 32366 5580 32506
rect 5540 32360 5592 32366
rect 5540 32302 5592 32308
rect 5540 32224 5592 32230
rect 5460 32172 5540 32178
rect 5460 32166 5592 32172
rect 5460 32150 5580 32166
rect 4528 32020 4580 32026
rect 4528 31962 4580 31968
rect 5172 32020 5224 32026
rect 5172 31962 5224 31968
rect 4066 31920 4122 31929
rect 4066 31855 4122 31864
rect 4712 31884 4764 31890
rect 4712 31826 4764 31832
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4724 31482 4752 31826
rect 5184 31822 5212 31962
rect 5172 31816 5224 31822
rect 5172 31758 5224 31764
rect 4896 31748 4948 31754
rect 4896 31690 4948 31696
rect 4712 31476 4764 31482
rect 4712 31418 4764 31424
rect 3976 31340 4028 31346
rect 3976 31282 4028 31288
rect 2964 31204 3016 31210
rect 2964 31146 3016 31152
rect 3700 31204 3752 31210
rect 3700 31146 3752 31152
rect 2504 30932 2556 30938
rect 2504 30874 2556 30880
rect 2780 30932 2832 30938
rect 2780 30874 2832 30880
rect 1674 30696 1730 30705
rect 2792 30648 2820 30874
rect 1674 30631 1676 30640
rect 1728 30631 1730 30640
rect 1676 30602 1728 30608
rect 2700 30620 2820 30648
rect 1400 30388 1452 30394
rect 1400 30330 1452 30336
rect 2320 30320 2372 30326
rect 2320 30262 2372 30268
rect 2332 29850 2360 30262
rect 2700 29850 2728 30620
rect 2976 30394 3004 31146
rect 3608 31136 3660 31142
rect 3608 31078 3660 31084
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 3620 30802 3648 31078
rect 4080 30938 4108 31078
rect 4068 30932 4120 30938
rect 4068 30874 4120 30880
rect 4908 30802 4936 31690
rect 5264 31204 5316 31210
rect 5264 31146 5316 31152
rect 5080 31136 5132 31142
rect 5276 31090 5304 31146
rect 5132 31084 5304 31090
rect 5080 31078 5304 31084
rect 5356 31136 5408 31142
rect 5356 31078 5408 31084
rect 5092 31062 5304 31078
rect 3608 30796 3660 30802
rect 3608 30738 3660 30744
rect 3976 30796 4028 30802
rect 3976 30738 4028 30744
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 3056 30592 3108 30598
rect 3056 30534 3108 30540
rect 2964 30388 3016 30394
rect 2964 30330 3016 30336
rect 3068 30190 3096 30534
rect 3988 30394 4016 30738
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4908 30394 4936 30738
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4896 30388 4948 30394
rect 4896 30330 4948 30336
rect 3056 30184 3108 30190
rect 3056 30126 3108 30132
rect 2320 29844 2372 29850
rect 2320 29786 2372 29792
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 3068 29782 3096 30126
rect 4068 30116 4120 30122
rect 4068 30058 4120 30064
rect 3056 29776 3108 29782
rect 3056 29718 3108 29724
rect 2780 29708 2832 29714
rect 2780 29650 2832 29656
rect 3884 29708 3936 29714
rect 3884 29650 3936 29656
rect 2504 29640 2556 29646
rect 2504 29582 2556 29588
rect 2516 29306 2544 29582
rect 2504 29300 2556 29306
rect 2504 29242 2556 29248
rect 2044 29096 2096 29102
rect 2044 29038 2096 29044
rect 1860 28688 1912 28694
rect 1860 28630 1912 28636
rect 1872 28218 1900 28630
rect 2056 28422 2084 29038
rect 2516 28694 2544 29242
rect 2792 29034 2820 29650
rect 2780 29028 2832 29034
rect 2780 28970 2832 28976
rect 2792 28762 2820 28970
rect 3896 28762 3924 29650
rect 4080 29306 4108 30058
rect 4620 29776 4672 29782
rect 4620 29718 4672 29724
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4632 29306 4660 29718
rect 5092 29306 5120 31062
rect 5368 30954 5396 31078
rect 5276 30926 5396 30954
rect 5460 30938 5488 32150
rect 5644 32042 5672 32694
rect 5552 32014 5672 32042
rect 5448 30932 5500 30938
rect 5276 30598 5304 30926
rect 5448 30874 5500 30880
rect 5448 30796 5500 30802
rect 5448 30738 5500 30744
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 5460 30682 5488 30738
rect 5552 30682 5580 32014
rect 5630 31920 5686 31929
rect 5630 31855 5632 31864
rect 5684 31855 5686 31864
rect 5632 31826 5684 31832
rect 5644 31482 5672 31826
rect 5736 31770 5764 34138
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 5828 33658 5856 34002
rect 5920 33998 5948 34478
rect 6104 34202 6132 34546
rect 6276 34400 6328 34406
rect 6276 34342 6328 34348
rect 6092 34196 6144 34202
rect 6092 34138 6144 34144
rect 5908 33992 5960 33998
rect 5908 33934 5960 33940
rect 5816 33652 5868 33658
rect 5816 33594 5868 33600
rect 5920 33454 5948 33934
rect 6288 33658 6316 34342
rect 6656 34134 6684 34886
rect 7300 34610 7328 35430
rect 7288 34604 7340 34610
rect 7288 34546 7340 34552
rect 7196 34400 7248 34406
rect 7196 34342 7248 34348
rect 6644 34128 6696 34134
rect 6644 34070 6696 34076
rect 6276 33652 6328 33658
rect 6276 33594 6328 33600
rect 6656 33590 6684 34070
rect 7208 33862 7236 34342
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 6644 33584 6696 33590
rect 6644 33526 6696 33532
rect 5908 33448 5960 33454
rect 5908 33390 5960 33396
rect 5920 33046 5948 33390
rect 6656 33386 6684 33526
rect 6828 33448 6880 33454
rect 6828 33390 6880 33396
rect 6644 33380 6696 33386
rect 6644 33322 6696 33328
rect 6840 33114 6868 33390
rect 7208 33318 7236 33798
rect 7392 33522 7420 35974
rect 7746 35864 7802 35873
rect 8312 35834 8340 39520
rect 9416 35873 9444 39520
rect 9402 35864 9458 35873
rect 7746 35799 7748 35808
rect 7800 35799 7802 35808
rect 8300 35828 8352 35834
rect 7748 35770 7800 35776
rect 9402 35799 9458 35808
rect 9586 35864 9642 35873
rect 9586 35799 9642 35808
rect 8300 35770 8352 35776
rect 8850 35592 8906 35601
rect 8850 35527 8852 35536
rect 8904 35527 8906 35536
rect 8852 35498 8904 35504
rect 9600 35465 9628 35799
rect 10520 35737 10548 39520
rect 10506 35728 10562 35737
rect 10506 35663 10562 35672
rect 10690 35728 10746 35737
rect 10690 35663 10746 35672
rect 9586 35456 9642 35465
rect 9586 35391 9642 35400
rect 10704 35222 10732 35663
rect 9496 35216 9548 35222
rect 9496 35158 9548 35164
rect 10692 35216 10744 35222
rect 10692 35158 10744 35164
rect 9128 35148 9180 35154
rect 9128 35090 9180 35096
rect 7472 34944 7524 34950
rect 7472 34886 7524 34892
rect 8300 34944 8352 34950
rect 8300 34886 8352 34892
rect 7484 34542 7512 34886
rect 7472 34536 7524 34542
rect 7472 34478 7524 34484
rect 7380 33516 7432 33522
rect 7380 33458 7432 33464
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 7208 33114 7236 33254
rect 6828 33108 6880 33114
rect 6828 33050 6880 33056
rect 7196 33108 7248 33114
rect 7196 33050 7248 33056
rect 5908 33040 5960 33046
rect 5908 32982 5960 32988
rect 7288 32972 7340 32978
rect 7288 32914 7340 32920
rect 6276 32904 6328 32910
rect 6276 32846 6328 32852
rect 6288 32570 6316 32846
rect 7300 32570 7328 32914
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 8208 32904 8260 32910
rect 8312 32892 8340 34886
rect 9140 34785 9168 35090
rect 9126 34776 9182 34785
rect 9508 34746 9536 35158
rect 9864 35148 9916 35154
rect 9864 35090 9916 35096
rect 9680 34944 9732 34950
rect 9680 34886 9732 34892
rect 9126 34711 9128 34720
rect 9180 34711 9182 34720
rect 9496 34740 9548 34746
rect 9128 34682 9180 34688
rect 9496 34682 9548 34688
rect 8852 34672 8904 34678
rect 8852 34614 8904 34620
rect 8392 34536 8444 34542
rect 8392 34478 8444 34484
rect 8404 33454 8432 34478
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8392 33448 8444 33454
rect 8392 33390 8444 33396
rect 8404 33114 8432 33390
rect 8680 33114 8708 33798
rect 8864 33454 8892 34614
rect 9312 34468 9364 34474
rect 9312 34410 9364 34416
rect 8852 33448 8904 33454
rect 8852 33390 8904 33396
rect 8392 33108 8444 33114
rect 8392 33050 8444 33056
rect 8668 33108 8720 33114
rect 8668 33050 8720 33056
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 8260 32864 8340 32892
rect 8208 32846 8260 32852
rect 6276 32564 6328 32570
rect 6276 32506 6328 32512
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 6288 32026 6316 32506
rect 7196 32224 7248 32230
rect 7196 32166 7248 32172
rect 7208 32026 7236 32166
rect 7300 32026 7328 32506
rect 7392 32434 7420 32846
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7852 32570 7880 32710
rect 7840 32564 7892 32570
rect 7840 32506 7892 32512
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 6276 32020 6328 32026
rect 6276 31962 6328 31968
rect 7196 32020 7248 32026
rect 7196 31962 7248 31968
rect 7288 32020 7340 32026
rect 7288 31962 7340 31968
rect 5736 31742 5948 31770
rect 5920 31686 5948 31742
rect 5724 31680 5776 31686
rect 5724 31622 5776 31628
rect 5908 31680 5960 31686
rect 5908 31622 5960 31628
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5736 31346 5764 31622
rect 7208 31482 7236 31962
rect 7392 31958 7420 32370
rect 7852 32366 7880 32506
rect 7840 32360 7892 32366
rect 7840 32302 7892 32308
rect 8404 32230 8432 32914
rect 8484 32496 8536 32502
rect 8484 32438 8536 32444
rect 8496 32298 8524 32438
rect 8680 32434 8708 33050
rect 8668 32428 8720 32434
rect 8668 32370 8720 32376
rect 8484 32292 8536 32298
rect 8484 32234 8536 32240
rect 8392 32224 8444 32230
rect 8392 32166 8444 32172
rect 8404 32026 8432 32166
rect 8392 32020 8444 32026
rect 8392 31962 8444 31968
rect 7380 31952 7432 31958
rect 7380 31894 7432 31900
rect 8496 31890 8524 32234
rect 8484 31884 8536 31890
rect 8484 31826 8536 31832
rect 8496 31482 8524 31826
rect 9324 31822 9352 34410
rect 9588 34400 9640 34406
rect 9586 34368 9588 34377
rect 9640 34368 9642 34377
rect 9586 34303 9642 34312
rect 9588 34196 9640 34202
rect 9692 34184 9720 34886
rect 9876 34746 9904 35090
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 10324 34944 10376 34950
rect 10324 34886 10376 34892
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 10140 34604 10192 34610
rect 10140 34546 10192 34552
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9640 34156 9720 34184
rect 9588 34138 9640 34144
rect 9784 34082 9812 34478
rect 10152 34134 10180 34546
rect 10336 34474 10364 34886
rect 10324 34468 10376 34474
rect 10324 34410 10376 34416
rect 11152 34400 11204 34406
rect 11152 34342 11204 34348
rect 11242 34368 11298 34377
rect 9600 34054 9812 34082
rect 10140 34128 10192 34134
rect 10140 34070 10192 34076
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 9416 33046 9444 33934
rect 9404 33040 9456 33046
rect 9404 32982 9456 32988
rect 9416 31890 9444 32982
rect 9600 32842 9628 34054
rect 10152 33658 10180 34070
rect 11060 33856 11112 33862
rect 11060 33798 11112 33804
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 10784 33584 10836 33590
rect 10782 33552 10784 33561
rect 10836 33552 10838 33561
rect 11072 33522 11100 33798
rect 10782 33487 10838 33496
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 11072 33402 11100 33458
rect 11164 33454 11192 34342
rect 11242 34303 11298 34312
rect 11256 33454 11284 34303
rect 11532 34066 11560 35022
rect 11624 34785 11652 39520
rect 12728 35737 12756 39520
rect 12714 35728 12770 35737
rect 12714 35663 12770 35672
rect 12256 35488 12308 35494
rect 12256 35430 12308 35436
rect 11796 35148 11848 35154
rect 11796 35090 11848 35096
rect 11610 34776 11666 34785
rect 11808 34746 11836 35090
rect 11610 34711 11666 34720
rect 11796 34740 11848 34746
rect 11796 34682 11848 34688
rect 11610 34096 11666 34105
rect 11520 34060 11572 34066
rect 11610 34031 11666 34040
rect 11796 34060 11848 34066
rect 11520 34002 11572 34008
rect 10980 33374 11100 33402
rect 11152 33448 11204 33454
rect 11152 33390 11204 33396
rect 11244 33448 11296 33454
rect 11244 33390 11296 33396
rect 10980 33114 11008 33374
rect 11256 33114 11284 33390
rect 10968 33108 11020 33114
rect 10968 33050 11020 33056
rect 11244 33108 11296 33114
rect 11244 33050 11296 33056
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9588 32836 9640 32842
rect 9588 32778 9640 32784
rect 9692 32366 9720 32914
rect 11624 32842 11652 34031
rect 11796 34002 11848 34008
rect 11808 33522 11836 34002
rect 11796 33516 11848 33522
rect 11796 33458 11848 33464
rect 12164 33312 12216 33318
rect 12164 33254 12216 33260
rect 12176 33114 12204 33254
rect 12164 33108 12216 33114
rect 12164 33050 12216 33056
rect 11612 32836 11664 32842
rect 11612 32778 11664 32784
rect 9864 32768 9916 32774
rect 9864 32710 9916 32716
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 9876 32609 9904 32710
rect 9862 32600 9918 32609
rect 9862 32535 9918 32544
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 11060 31952 11112 31958
rect 11060 31894 11112 31900
rect 9404 31884 9456 31890
rect 9404 31826 9456 31832
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 9416 31482 9444 31826
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 7196 31476 7248 31482
rect 7196 31418 7248 31424
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8576 31476 8628 31482
rect 8576 31418 8628 31424
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 5724 31340 5776 31346
rect 5724 31282 5776 31288
rect 6276 30864 6328 30870
rect 6276 30806 6328 30812
rect 5264 30592 5316 30598
rect 5264 30534 5316 30540
rect 5276 30394 5304 30534
rect 5264 30388 5316 30394
rect 5264 30330 5316 30336
rect 5368 30190 5396 30670
rect 5460 30654 5580 30682
rect 5552 30258 5580 30654
rect 5906 30696 5962 30705
rect 5906 30631 5962 30640
rect 5920 30326 5948 30631
rect 5908 30320 5960 30326
rect 5908 30262 5960 30268
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 6000 30252 6052 30258
rect 6000 30194 6052 30200
rect 5356 30184 5408 30190
rect 5356 30126 5408 30132
rect 5368 29714 5396 30126
rect 6012 29850 6040 30194
rect 6288 30054 6316 30806
rect 7010 30696 7066 30705
rect 7010 30631 7012 30640
rect 7064 30631 7066 30640
rect 7012 30602 7064 30608
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 6460 30184 6512 30190
rect 6460 30126 6512 30132
rect 6276 30048 6328 30054
rect 6276 29990 6328 29996
rect 6288 29850 6316 29990
rect 6000 29844 6052 29850
rect 6000 29786 6052 29792
rect 6276 29844 6328 29850
rect 6276 29786 6328 29792
rect 5356 29708 5408 29714
rect 5356 29650 5408 29656
rect 4068 29300 4120 29306
rect 4620 29300 4672 29306
rect 4120 29260 4200 29288
rect 4068 29242 4120 29248
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 3884 28756 3936 28762
rect 3884 28698 3936 28704
rect 4172 28694 4200 29260
rect 4620 29242 4672 29248
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 4632 28762 4660 29242
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 2504 28688 2556 28694
rect 2504 28630 2556 28636
rect 4160 28688 4212 28694
rect 4160 28630 4212 28636
rect 2044 28416 2096 28422
rect 2044 28358 2096 28364
rect 1860 28212 1912 28218
rect 1860 28154 1912 28160
rect 2056 27878 2084 28358
rect 2044 27872 2096 27878
rect 2044 27814 2096 27820
rect 2056 27606 2084 27814
rect 2516 27674 2544 28630
rect 4172 28506 4200 28630
rect 4080 28478 4200 28506
rect 4080 28218 4108 28478
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 5368 28218 5396 29650
rect 5632 29572 5684 29578
rect 5632 29514 5684 29520
rect 5644 29170 5672 29514
rect 6012 29170 6040 29786
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 6000 29164 6052 29170
rect 6000 29106 6052 29112
rect 6288 29102 6316 29786
rect 6472 29646 6500 30126
rect 6748 30122 6776 30534
rect 7024 30190 7052 30602
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 7012 30184 7064 30190
rect 7012 30126 7064 30132
rect 6736 30116 6788 30122
rect 6736 30058 6788 30064
rect 8392 30048 8444 30054
rect 8392 29990 8444 29996
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6460 29640 6512 29646
rect 6460 29582 6512 29588
rect 6472 29170 6500 29582
rect 6564 29306 6592 29650
rect 7748 29640 7800 29646
rect 7748 29582 7800 29588
rect 6552 29300 6604 29306
rect 6552 29242 6604 29248
rect 7760 29170 7788 29582
rect 6460 29164 6512 29170
rect 6460 29106 6512 29112
rect 7748 29164 7800 29170
rect 7748 29106 7800 29112
rect 5816 29096 5868 29102
rect 5816 29038 5868 29044
rect 6276 29096 6328 29102
rect 6276 29038 6328 29044
rect 5828 28762 5856 29038
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8312 28762 8340 28970
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 7288 28620 7340 28626
rect 7288 28562 7340 28568
rect 7300 28218 7328 28562
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 4068 28212 4120 28218
rect 4068 28154 4120 28160
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 7288 28212 7340 28218
rect 7288 28154 7340 28160
rect 7564 28008 7616 28014
rect 7564 27950 7616 27956
rect 7288 27940 7340 27946
rect 7288 27882 7340 27888
rect 2504 27668 2556 27674
rect 2504 27610 2556 27616
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 1676 27532 1728 27538
rect 1676 27474 1728 27480
rect 1688 26858 1716 27474
rect 2056 27130 2084 27542
rect 7300 27538 7328 27882
rect 7576 27878 7604 27950
rect 7852 27946 7880 28358
rect 8312 28218 8340 28698
rect 8404 28626 8432 29990
rect 8496 29646 8524 30534
rect 8588 30190 8616 31418
rect 9600 31346 9628 31758
rect 11072 31498 11100 31894
rect 11532 31890 11560 32710
rect 12176 32570 12204 33050
rect 12268 33046 12296 35430
rect 12532 35284 12584 35290
rect 12532 35226 12584 35232
rect 12440 34740 12492 34746
rect 12440 34682 12492 34688
rect 12348 34604 12400 34610
rect 12348 34546 12400 34552
rect 12256 33040 12308 33046
rect 12256 32982 12308 32988
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 12268 32502 12296 32982
rect 12360 32910 12388 34546
rect 12452 34202 12480 34682
rect 12544 34542 12572 35226
rect 12808 34944 12860 34950
rect 13820 34944 13872 34950
rect 12808 34886 12860 34892
rect 13634 34912 13690 34921
rect 12820 34542 12848 34886
rect 13820 34886 13872 34892
rect 13634 34847 13690 34856
rect 12532 34536 12584 34542
rect 12532 34478 12584 34484
rect 12808 34536 12860 34542
rect 12808 34478 12860 34484
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12992 34196 13044 34202
rect 12992 34138 13044 34144
rect 12622 33960 12678 33969
rect 12622 33895 12678 33904
rect 12348 32904 12400 32910
rect 12348 32846 12400 32852
rect 12532 32904 12584 32910
rect 12532 32846 12584 32852
rect 12544 32570 12572 32846
rect 12636 32842 12664 33895
rect 12806 33552 12862 33561
rect 13004 33522 13032 34138
rect 12806 33487 12862 33496
rect 12992 33516 13044 33522
rect 12820 33454 12848 33487
rect 12992 33458 13044 33464
rect 12808 33448 12860 33454
rect 12808 33390 12860 33396
rect 12820 33114 12848 33390
rect 12900 33380 12952 33386
rect 12900 33322 12952 33328
rect 12912 33289 12940 33322
rect 12898 33280 12954 33289
rect 12898 33215 12954 33224
rect 13648 33114 13676 34847
rect 12808 33108 12860 33114
rect 12808 33050 12860 33056
rect 13636 33108 13688 33114
rect 13636 33050 13688 33056
rect 13268 32972 13320 32978
rect 13268 32914 13320 32920
rect 12624 32836 12676 32842
rect 12624 32778 12676 32784
rect 13280 32609 13308 32914
rect 13266 32600 13322 32609
rect 12532 32564 12584 32570
rect 13266 32535 13268 32544
rect 12532 32506 12584 32512
rect 13320 32535 13322 32544
rect 13268 32506 13320 32512
rect 12256 32496 12308 32502
rect 12256 32438 12308 32444
rect 11520 31884 11572 31890
rect 11520 31826 11572 31832
rect 10980 31482 11100 31498
rect 10968 31476 11100 31482
rect 11020 31470 11100 31476
rect 10968 31418 11020 31424
rect 11532 31414 11560 31826
rect 12348 31680 12400 31686
rect 12348 31622 12400 31628
rect 11886 31512 11942 31521
rect 11886 31447 11888 31456
rect 11940 31447 11942 31456
rect 11888 31418 11940 31424
rect 11520 31408 11572 31414
rect 11520 31350 11572 31356
rect 9220 31340 9272 31346
rect 9220 31282 9272 31288
rect 9588 31340 9640 31346
rect 9588 31282 9640 31288
rect 8668 31272 8720 31278
rect 8668 31214 8720 31220
rect 8680 30802 8708 31214
rect 8668 30796 8720 30802
rect 8668 30738 8720 30744
rect 8576 30184 8628 30190
rect 8576 30126 8628 30132
rect 8588 29850 8616 30126
rect 8576 29844 8628 29850
rect 8576 29786 8628 29792
rect 8680 29714 8708 30738
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9140 28626 9168 28902
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 7840 27940 7892 27946
rect 7840 27882 7892 27888
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 7748 27872 7800 27878
rect 7748 27814 7800 27820
rect 8206 27840 8262 27849
rect 6644 27532 6696 27538
rect 6644 27474 6696 27480
rect 7288 27532 7340 27538
rect 7288 27474 7340 27480
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 6656 27130 6684 27474
rect 2044 27124 2096 27130
rect 2044 27066 2096 27072
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 2700 26858 2820 26874
rect 1676 26852 1728 26858
rect 1676 26794 1728 26800
rect 2688 26852 2820 26858
rect 2740 26846 2820 26852
rect 2688 26794 2740 26800
rect 2792 20097 2820 26846
rect 7300 26790 7328 27474
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 7300 26586 7328 26726
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7576 26518 7604 27814
rect 7760 27130 7788 27814
rect 8206 27775 8262 27784
rect 8220 27130 8248 27775
rect 8312 27674 8340 28154
rect 8680 28082 8708 28494
rect 9232 28082 9260 31282
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 9864 31204 9916 31210
rect 9864 31146 9916 31152
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9600 29084 9628 31078
rect 9784 30734 9812 31078
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9876 30394 9904 31146
rect 11164 30977 11192 31214
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11150 30968 11206 30977
rect 11150 30903 11206 30912
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9864 30388 9916 30394
rect 9864 30330 9916 30336
rect 9876 29782 9904 30330
rect 9864 29776 9916 29782
rect 9864 29718 9916 29724
rect 9772 29708 9824 29714
rect 9772 29650 9824 29656
rect 9680 29096 9732 29102
rect 9600 29056 9680 29084
rect 9680 29038 9732 29044
rect 9784 28558 9812 29650
rect 9876 29238 9904 29718
rect 9968 29306 9996 30738
rect 10692 30728 10744 30734
rect 10692 30670 10744 30676
rect 10704 30054 10732 30670
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10782 30424 10838 30433
rect 10782 30359 10838 30368
rect 10796 30326 10824 30359
rect 10784 30320 10836 30326
rect 10784 30262 10836 30268
rect 11072 30190 11100 30534
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 10232 30048 10284 30054
rect 10232 29990 10284 29996
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 9864 29232 9916 29238
rect 9864 29174 9916 29180
rect 10244 28762 10272 29990
rect 10704 29850 10732 29990
rect 10692 29844 10744 29850
rect 10692 29786 10744 29792
rect 11060 29640 11112 29646
rect 11060 29582 11112 29588
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10232 28620 10284 28626
rect 10232 28562 10284 28568
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 8668 28076 8720 28082
rect 8668 28018 8720 28024
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 9232 27878 9260 28018
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 7748 27124 7800 27130
rect 7748 27066 7800 27072
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 7760 26926 7788 27066
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 7748 26920 7800 26926
rect 7748 26862 7800 26868
rect 7840 26784 7892 26790
rect 7840 26726 7892 26732
rect 6920 26512 6972 26518
rect 6920 26454 6972 26460
rect 7564 26512 7616 26518
rect 7564 26454 7616 26460
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 6932 26042 6960 26454
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 7024 25838 7052 26386
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7024 25362 7052 25774
rect 7104 25764 7156 25770
rect 7104 25706 7156 25712
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 7024 24954 7052 25298
rect 7116 25158 7144 25706
rect 7196 25356 7248 25362
rect 7196 25298 7248 25304
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 7208 24410 7236 25298
rect 7380 24744 7432 24750
rect 7380 24686 7432 24692
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 7392 24138 7420 24686
rect 7656 24676 7708 24682
rect 7656 24618 7708 24624
rect 7668 24585 7696 24618
rect 7654 24576 7710 24585
rect 7654 24511 7710 24520
rect 7852 24410 7880 26726
rect 8864 26586 8892 26930
rect 8852 26580 8904 26586
rect 8852 26522 8904 26528
rect 8208 26512 8260 26518
rect 8208 26454 8260 26460
rect 8220 26024 8248 26454
rect 8300 26036 8352 26042
rect 8220 25996 8300 26024
rect 8300 25978 8352 25984
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7932 24336 7984 24342
rect 7932 24278 7984 24284
rect 7380 24132 7432 24138
rect 7380 24074 7432 24080
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 7944 23866 7972 24278
rect 8220 24274 8248 25094
rect 9232 24857 9260 27814
rect 9508 27674 9536 28494
rect 10244 27878 10272 28562
rect 10428 28490 10456 28902
rect 10612 28762 10640 29106
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 10600 28756 10652 28762
rect 10600 28698 10652 28704
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10980 28218 11008 28902
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 10232 27872 10284 27878
rect 10230 27840 10232 27849
rect 10284 27840 10286 27849
rect 10230 27775 10286 27784
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 10138 27568 10194 27577
rect 9956 27532 10008 27538
rect 11072 27538 11100 29582
rect 11348 29306 11376 31078
rect 11532 30938 11560 31350
rect 11900 31278 11928 31418
rect 11888 31272 11940 31278
rect 11888 31214 11940 31220
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11428 30252 11480 30258
rect 11428 30194 11480 30200
rect 11440 29850 11468 30194
rect 11428 29844 11480 29850
rect 11428 29786 11480 29792
rect 11440 29306 11468 29786
rect 11336 29300 11388 29306
rect 11336 29242 11388 29248
rect 11428 29300 11480 29306
rect 11428 29242 11480 29248
rect 11348 28082 11376 29242
rect 12360 28694 12388 31622
rect 13544 31272 13596 31278
rect 13544 31214 13596 31220
rect 13084 31136 13136 31142
rect 12714 31104 12770 31113
rect 13084 31078 13136 31084
rect 12714 31039 12770 31048
rect 12728 30938 12756 31039
rect 13096 30938 13124 31078
rect 13556 30938 13584 31214
rect 12716 30932 12768 30938
rect 12716 30874 12768 30880
rect 13084 30932 13136 30938
rect 13084 30874 13136 30880
rect 13544 30932 13596 30938
rect 13544 30874 13596 30880
rect 12728 30433 12756 30874
rect 12900 30660 12952 30666
rect 12900 30602 12952 30608
rect 12714 30424 12770 30433
rect 12714 30359 12770 30368
rect 12440 30116 12492 30122
rect 12440 30058 12492 30064
rect 12452 29238 12480 30058
rect 12728 30054 12756 30359
rect 12912 30190 12940 30602
rect 13096 30258 13124 30874
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13740 30433 13768 30738
rect 13726 30424 13782 30433
rect 13726 30359 13728 30368
rect 13780 30359 13782 30368
rect 13728 30330 13780 30336
rect 13084 30252 13136 30258
rect 13084 30194 13136 30200
rect 12900 30184 12952 30190
rect 12900 30126 12952 30132
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 12440 29232 12492 29238
rect 12440 29174 12492 29180
rect 12348 28688 12400 28694
rect 12348 28630 12400 28636
rect 12360 28218 12388 28630
rect 12348 28212 12400 28218
rect 12348 28154 12400 28160
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11152 27872 11204 27878
rect 11152 27814 11204 27820
rect 11164 27674 11192 27814
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 11060 27532 11112 27538
rect 10138 27503 10194 27512
rect 9956 27474 10008 27480
rect 9968 27130 9996 27474
rect 10152 27402 10180 27503
rect 10980 27492 11060 27520
rect 10140 27396 10192 27402
rect 10140 27338 10192 27344
rect 9956 27124 10008 27130
rect 9956 27066 10008 27072
rect 10980 26926 11008 27492
rect 11060 27474 11112 27480
rect 11348 26994 11376 28018
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 12348 27668 12400 27674
rect 12348 27610 12400 27616
rect 11796 27532 11848 27538
rect 11796 27474 11848 27480
rect 11808 27130 11836 27474
rect 12268 27130 12296 27610
rect 12360 27538 12388 27610
rect 12452 27538 12480 29174
rect 12636 28626 12664 29990
rect 12912 29782 12940 30126
rect 12900 29776 12952 29782
rect 12900 29718 12952 29724
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12728 29102 12756 29446
rect 12912 29306 12940 29718
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 13832 29186 13860 34886
rect 13924 31482 13952 39520
rect 14004 36032 14056 36038
rect 14004 35974 14056 35980
rect 14016 35630 14044 35974
rect 15028 35714 15056 39520
rect 15660 36236 15712 36242
rect 15660 36178 15712 36184
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 14844 35686 15056 35714
rect 14004 35624 14056 35630
rect 14004 35566 14056 35572
rect 14016 35290 14044 35566
rect 14004 35284 14056 35290
rect 14004 35226 14056 35232
rect 14740 35284 14792 35290
rect 14740 35226 14792 35232
rect 14016 34202 14044 35226
rect 14188 35148 14240 35154
rect 14188 35090 14240 35096
rect 14648 35148 14700 35154
rect 14648 35090 14700 35096
rect 14200 34785 14228 35090
rect 14186 34776 14242 34785
rect 14660 34746 14688 35090
rect 14186 34711 14188 34720
rect 14240 34711 14242 34720
rect 14648 34740 14700 34746
rect 14188 34682 14240 34688
rect 14648 34682 14700 34688
rect 14280 34672 14332 34678
rect 14280 34614 14332 34620
rect 14292 34474 14320 34614
rect 14280 34468 14332 34474
rect 14280 34410 14332 34416
rect 14004 34196 14056 34202
rect 14004 34138 14056 34144
rect 14292 33862 14320 34410
rect 14660 34202 14688 34682
rect 14752 34610 14780 35226
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 14752 33998 14780 34546
rect 14740 33992 14792 33998
rect 14740 33934 14792 33940
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 14096 32904 14148 32910
rect 14094 32872 14096 32881
rect 14148 32872 14150 32881
rect 14094 32807 14150 32816
rect 14108 32434 14136 32807
rect 14200 32570 14228 33254
rect 14292 32910 14320 33798
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 14188 32564 14240 32570
rect 14188 32506 14240 32512
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14200 32366 14228 32506
rect 14188 32360 14240 32366
rect 14188 32302 14240 32308
rect 14292 32026 14320 32846
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14844 31521 14872 35686
rect 14924 34060 14976 34066
rect 14924 34002 14976 34008
rect 14936 33114 14964 34002
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 15120 33114 15148 33458
rect 14924 33108 14976 33114
rect 14924 33050 14976 33056
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 15120 32570 15148 33050
rect 15108 32564 15160 32570
rect 15108 32506 15160 32512
rect 14922 32464 14978 32473
rect 15212 32450 15240 35974
rect 15672 35766 15700 36178
rect 15752 36168 15804 36174
rect 15752 36110 15804 36116
rect 15936 36168 15988 36174
rect 15936 36110 15988 36116
rect 15764 35834 15792 36110
rect 15752 35828 15804 35834
rect 15752 35770 15804 35776
rect 15660 35760 15712 35766
rect 15658 35728 15660 35737
rect 15712 35728 15714 35737
rect 15658 35663 15714 35672
rect 15384 35624 15436 35630
rect 15384 35566 15436 35572
rect 15396 35494 15424 35566
rect 15384 35488 15436 35494
rect 15384 35430 15436 35436
rect 15292 35284 15344 35290
rect 15292 35226 15344 35232
rect 15304 35193 15332 35226
rect 15290 35184 15346 35193
rect 15290 35119 15346 35128
rect 15396 34066 15424 35430
rect 15764 35170 15792 35770
rect 15948 35630 15976 36110
rect 15936 35624 15988 35630
rect 15936 35566 15988 35572
rect 15844 35556 15896 35562
rect 15844 35498 15896 35504
rect 15672 35142 15792 35170
rect 15384 34060 15436 34066
rect 15384 34002 15436 34008
rect 15672 33561 15700 35142
rect 15856 35086 15884 35498
rect 15752 35080 15804 35086
rect 15752 35022 15804 35028
rect 15844 35080 15896 35086
rect 15844 35022 15896 35028
rect 15764 34921 15792 35022
rect 15750 34912 15806 34921
rect 15750 34847 15806 34856
rect 15764 34678 15792 34847
rect 15856 34746 15884 35022
rect 16132 34785 16160 39520
rect 17236 35714 17264 39520
rect 16960 35686 17264 35714
rect 18340 35714 18368 39520
rect 18340 35686 18552 35714
rect 16854 35048 16910 35057
rect 16854 34983 16856 34992
rect 16908 34983 16910 34992
rect 16856 34954 16908 34960
rect 16118 34776 16174 34785
rect 15844 34740 15896 34746
rect 16118 34711 16174 34720
rect 15844 34682 15896 34688
rect 15752 34672 15804 34678
rect 15752 34614 15804 34620
rect 16212 33856 16264 33862
rect 16212 33798 16264 33804
rect 16672 33856 16724 33862
rect 16672 33798 16724 33804
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 15948 33561 15976 33594
rect 15658 33552 15714 33561
rect 15658 33487 15714 33496
rect 15934 33552 15990 33561
rect 15934 33487 15936 33496
rect 15988 33487 15990 33496
rect 15936 33458 15988 33464
rect 15568 33448 15620 33454
rect 15568 33390 15620 33396
rect 15292 33312 15344 33318
rect 15292 33254 15344 33260
rect 15304 32978 15332 33254
rect 15580 32978 15608 33390
rect 16026 33280 16082 33289
rect 16026 33215 16082 33224
rect 16040 32978 16068 33215
rect 15292 32972 15344 32978
rect 15292 32914 15344 32920
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 16028 32972 16080 32978
rect 16028 32914 16080 32920
rect 14922 32399 14924 32408
rect 14976 32399 14978 32408
rect 15120 32422 15240 32450
rect 14924 32370 14976 32376
rect 14936 31958 14964 32370
rect 15120 32366 15148 32422
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 15304 32314 15332 32914
rect 15580 32570 15608 32914
rect 15752 32904 15804 32910
rect 15752 32846 15804 32852
rect 15568 32564 15620 32570
rect 15620 32524 15700 32552
rect 15568 32506 15620 32512
rect 15120 32026 15148 32302
rect 15304 32286 15608 32314
rect 15580 32026 15608 32286
rect 15108 32020 15160 32026
rect 15108 31962 15160 31968
rect 15568 32020 15620 32026
rect 15568 31962 15620 31968
rect 14924 31952 14976 31958
rect 14924 31894 14976 31900
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 14830 31512 14886 31521
rect 13912 31476 13964 31482
rect 14830 31447 14886 31456
rect 13912 31418 13964 31424
rect 14372 31272 14424 31278
rect 14372 31214 14424 31220
rect 14384 30977 14412 31214
rect 14370 30968 14426 30977
rect 14370 30903 14372 30912
rect 14424 30903 14426 30912
rect 14372 30874 14424 30880
rect 14556 30796 14608 30802
rect 14556 30738 14608 30744
rect 14280 30592 14332 30598
rect 14280 30534 14332 30540
rect 14292 30190 14320 30534
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14280 30184 14332 30190
rect 14280 30126 14332 30132
rect 14200 29714 14228 30126
rect 14292 29850 14320 30126
rect 14280 29844 14332 29850
rect 14280 29786 14332 29792
rect 14188 29708 14240 29714
rect 14188 29650 14240 29656
rect 14004 29504 14056 29510
rect 14004 29446 14056 29452
rect 13740 29170 13860 29186
rect 13728 29164 13860 29170
rect 13780 29158 13860 29164
rect 13728 29106 13780 29112
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12728 27577 12756 29038
rect 13740 29034 13860 29050
rect 13740 29028 13872 29034
rect 13740 29022 13820 29028
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 12992 28416 13044 28422
rect 12992 28358 13044 28364
rect 12820 28014 12848 28358
rect 13004 28082 13032 28358
rect 13464 28218 13492 28562
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12808 28008 12860 28014
rect 12808 27950 12860 27956
rect 12820 27674 12848 27950
rect 12808 27668 12860 27674
rect 12808 27610 12860 27616
rect 12714 27568 12770 27577
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12440 27532 12492 27538
rect 12714 27503 12770 27512
rect 12440 27474 12492 27480
rect 12348 27328 12400 27334
rect 12348 27270 12400 27276
rect 12900 27328 12952 27334
rect 13004 27316 13032 28018
rect 13452 27532 13504 27538
rect 13452 27474 13504 27480
rect 12952 27288 13032 27316
rect 12900 27270 12952 27276
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 12256 27124 12308 27130
rect 12256 27066 12308 27072
rect 12360 26994 12388 27270
rect 12912 27062 12940 27270
rect 13464 27130 13492 27474
rect 13740 27402 13768 29022
rect 13820 28970 13872 28976
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 12900 27056 12952 27062
rect 12900 26998 12952 27004
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10980 26382 11008 26862
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 11072 26518 11100 26726
rect 11348 26586 11376 26930
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 26790 11836 26862
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 11796 26784 11848 26790
rect 11796 26726 11848 26732
rect 12360 26738 12388 26794
rect 12532 26784 12584 26790
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11060 26512 11112 26518
rect 11060 26454 11112 26460
rect 11808 26450 11836 26726
rect 12360 26710 12480 26738
rect 12532 26726 12584 26732
rect 12348 26512 12400 26518
rect 12348 26454 12400 26460
rect 11796 26444 11848 26450
rect 11796 26386 11848 26392
rect 10968 26376 11020 26382
rect 10414 26344 10470 26353
rect 10968 26318 11020 26324
rect 10414 26279 10470 26288
rect 10428 25838 10456 26279
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 9692 24954 9720 25774
rect 10692 25764 10744 25770
rect 10692 25706 10744 25712
rect 10704 25498 10732 25706
rect 10980 25498 11008 26318
rect 11808 26042 11836 26386
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 12360 25922 12388 26454
rect 12452 26042 12480 26710
rect 12544 26353 12572 26726
rect 12530 26344 12586 26353
rect 12530 26279 12532 26288
rect 12584 26279 12586 26288
rect 12532 26250 12584 26256
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12360 25894 12480 25922
rect 12912 25906 12940 26998
rect 14016 26790 14044 29446
rect 14292 29170 14320 29786
rect 14568 29510 14596 30738
rect 15016 29708 15068 29714
rect 15016 29650 15068 29656
rect 14556 29504 14608 29510
rect 14556 29446 14608 29452
rect 15028 29170 15056 29650
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 14280 29164 14332 29170
rect 14280 29106 14332 29112
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 14292 28694 14320 29106
rect 14464 28960 14516 28966
rect 14464 28902 14516 28908
rect 14476 28762 14504 28902
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14280 28688 14332 28694
rect 14280 28630 14332 28636
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14660 28218 14688 28494
rect 15028 28422 15056 29106
rect 15212 28694 15240 29174
rect 15304 28762 15332 31758
rect 15476 31272 15528 31278
rect 15476 31214 15528 31220
rect 15488 31113 15516 31214
rect 15474 31104 15530 31113
rect 15474 31039 15530 31048
rect 15580 30954 15608 31962
rect 15488 30926 15608 30954
rect 15384 29708 15436 29714
rect 15384 29650 15436 29656
rect 15396 29102 15424 29650
rect 15488 29646 15516 30926
rect 15568 30864 15620 30870
rect 15568 30806 15620 30812
rect 15580 30054 15608 30806
rect 15672 30122 15700 32524
rect 15764 32502 15792 32846
rect 15752 32496 15804 32502
rect 15752 32438 15804 32444
rect 16040 31958 16068 32914
rect 16224 32910 16252 33798
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 16224 32570 16252 32846
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 16684 32473 16712 33798
rect 16762 32872 16818 32881
rect 16762 32807 16818 32816
rect 16776 32774 16804 32807
rect 16764 32768 16816 32774
rect 16764 32710 16816 32716
rect 16670 32464 16726 32473
rect 16670 32399 16726 32408
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16028 31952 16080 31958
rect 16028 31894 16080 31900
rect 16486 31648 16542 31657
rect 16486 31583 16542 31592
rect 16500 31482 16528 31583
rect 16488 31476 16540 31482
rect 16488 31418 16540 31424
rect 16500 30258 16528 31418
rect 16592 31414 16620 32302
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 15660 30116 15712 30122
rect 15660 30058 15712 30064
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15476 29640 15528 29646
rect 15476 29582 15528 29588
rect 15384 29096 15436 29102
rect 15384 29038 15436 29044
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15200 28688 15252 28694
rect 15200 28630 15252 28636
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 15304 28218 15332 28698
rect 15580 28558 15608 29990
rect 15672 29850 15700 30058
rect 16592 30054 16620 30534
rect 16776 30190 16804 32710
rect 16960 30433 16988 35686
rect 17958 35320 18014 35329
rect 17958 35255 18014 35264
rect 17224 35148 17276 35154
rect 17224 35090 17276 35096
rect 17040 35012 17092 35018
rect 17040 34954 17092 34960
rect 17052 33862 17080 34954
rect 17236 34746 17264 35090
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 17328 33862 17356 35022
rect 17972 34921 18000 35255
rect 18052 34944 18104 34950
rect 17958 34912 18014 34921
rect 18052 34886 18104 34892
rect 17958 34847 18014 34856
rect 17960 34604 18012 34610
rect 17880 34564 17960 34592
rect 17684 34536 17736 34542
rect 17684 34478 17736 34484
rect 17040 33856 17092 33862
rect 17040 33798 17092 33804
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 17052 33658 17080 33798
rect 17040 33652 17092 33658
rect 17040 33594 17092 33600
rect 17040 33312 17092 33318
rect 17038 33280 17040 33289
rect 17092 33280 17094 33289
rect 17038 33215 17094 33224
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17604 32609 17632 32846
rect 17590 32600 17646 32609
rect 17590 32535 17646 32544
rect 17696 32434 17724 34478
rect 17776 33856 17828 33862
rect 17776 33798 17828 33804
rect 17684 32428 17736 32434
rect 17684 32370 17736 32376
rect 17038 31512 17094 31521
rect 17038 31447 17040 31456
rect 17092 31447 17094 31456
rect 17040 31418 17092 31424
rect 17052 30802 17080 31418
rect 17788 30938 17816 33798
rect 17880 32026 17908 34564
rect 17960 34546 18012 34552
rect 18064 33300 18092 34886
rect 18144 34672 18196 34678
rect 18142 34640 18144 34649
rect 18196 34640 18198 34649
rect 18142 34575 18198 34584
rect 18144 34128 18196 34134
rect 18144 34070 18196 34076
rect 18156 33318 18184 34070
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18340 33386 18368 33594
rect 18328 33380 18380 33386
rect 18328 33322 18380 33328
rect 17972 33272 18092 33300
rect 18144 33312 18196 33318
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 17868 31748 17920 31754
rect 17868 31690 17920 31696
rect 17880 31482 17908 31690
rect 17868 31476 17920 31482
rect 17868 31418 17920 31424
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 17040 30796 17092 30802
rect 17040 30738 17092 30744
rect 17776 30728 17828 30734
rect 17776 30670 17828 30676
rect 16946 30424 17002 30433
rect 16946 30359 17002 30368
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16396 30048 16448 30054
rect 16580 30048 16632 30054
rect 16396 29990 16448 29996
rect 16500 29996 16580 30002
rect 16500 29990 16632 29996
rect 15660 29844 15712 29850
rect 15660 29786 15712 29792
rect 15672 29306 15700 29786
rect 15844 29640 15896 29646
rect 15842 29608 15844 29617
rect 16304 29640 16356 29646
rect 15896 29608 15898 29617
rect 16304 29582 16356 29588
rect 15842 29543 15898 29552
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 15844 28688 15896 28694
rect 15844 28630 15896 28636
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15292 27940 15344 27946
rect 15292 27882 15344 27888
rect 15304 27130 15332 27882
rect 15396 27334 15424 28358
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15580 27674 15608 27950
rect 15856 27674 15884 28630
rect 16316 28422 16344 29582
rect 16304 28416 16356 28422
rect 16304 28358 16356 28364
rect 16316 28218 16344 28358
rect 16408 28218 16436 29990
rect 16500 29974 16620 29990
rect 16500 28490 16528 29974
rect 16776 29714 16804 30126
rect 16764 29708 16816 29714
rect 16764 29650 16816 29656
rect 17328 29306 17356 30194
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17512 29850 17540 29990
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17788 29306 17816 30670
rect 16580 29300 16632 29306
rect 16580 29242 16632 29248
rect 17316 29300 17368 29306
rect 17316 29242 17368 29248
rect 17776 29300 17828 29306
rect 17776 29242 17828 29248
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16304 28212 16356 28218
rect 16304 28154 16356 28160
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 16592 28098 16620 29242
rect 17328 29102 17356 29242
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16500 28082 16620 28098
rect 16488 28076 16620 28082
rect 16540 28070 16620 28076
rect 16488 28018 16540 28024
rect 16868 28014 16896 28494
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 15568 27668 15620 27674
rect 15568 27610 15620 27616
rect 15844 27668 15896 27674
rect 15844 27610 15896 27616
rect 17038 27568 17094 27577
rect 16488 27532 16540 27538
rect 17038 27503 17094 27512
rect 16488 27474 16540 27480
rect 15384 27328 15436 27334
rect 15384 27270 15436 27276
rect 15292 27124 15344 27130
rect 15292 27066 15344 27072
rect 15292 26920 15344 26926
rect 15396 26908 15424 27270
rect 16500 27130 16528 27474
rect 16672 27328 16724 27334
rect 16672 27270 16724 27276
rect 16488 27124 16540 27130
rect 16488 27066 16540 27072
rect 15344 26880 15424 26908
rect 15292 26862 15344 26868
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 11520 25696 11572 25702
rect 11520 25638 11572 25644
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 10060 24954 10088 25298
rect 10704 25294 10732 25434
rect 11532 25362 11560 25638
rect 11520 25356 11572 25362
rect 11520 25298 11572 25304
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 9680 24948 9732 24954
rect 9680 24890 9732 24896
rect 10048 24948 10100 24954
rect 10048 24890 10100 24896
rect 8482 24848 8538 24857
rect 8482 24783 8538 24792
rect 9218 24848 9274 24857
rect 9218 24783 9274 24792
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8220 23866 8248 24210
rect 8496 24206 8524 24783
rect 10152 24750 10180 25094
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 8760 24608 8812 24614
rect 8760 24550 8812 24556
rect 8772 24342 8800 24550
rect 8760 24336 8812 24342
rect 8760 24278 8812 24284
rect 10152 24206 10180 24686
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10244 24410 10272 24618
rect 10704 24426 10732 25230
rect 11060 25152 11112 25158
rect 10980 25112 11060 25140
rect 10232 24404 10284 24410
rect 10704 24398 10824 24426
rect 10232 24346 10284 24352
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 8484 24200 8536 24206
rect 8484 24142 8536 24148
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 8496 23866 8524 24142
rect 7932 23860 7984 23866
rect 7932 23802 7984 23808
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8484 23860 8536 23866
rect 8484 23802 8536 23808
rect 10428 23798 10456 24142
rect 10704 23866 10732 24210
rect 10796 23866 10824 24398
rect 10980 24342 11008 25112
rect 11060 25094 11112 25100
rect 12452 24954 12480 25894
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12544 25498 12572 25638
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12544 25158 12572 25434
rect 12912 25158 12940 25842
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12912 24886 12940 25094
rect 12900 24880 12952 24886
rect 11886 24848 11942 24857
rect 11886 24783 11888 24792
rect 11940 24783 11942 24792
rect 12898 24848 12900 24857
rect 12952 24848 12954 24857
rect 12898 24783 12954 24792
rect 11888 24754 11940 24760
rect 12912 24757 12940 24783
rect 11520 24608 11572 24614
rect 11518 24576 11520 24585
rect 12164 24608 12216 24614
rect 11572 24576 11574 24585
rect 12164 24550 12216 24556
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 11518 24511 11574 24520
rect 11532 24342 11560 24511
rect 12176 24410 12204 24550
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12544 24342 12572 24550
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 12532 24336 12584 24342
rect 12532 24278 12584 24284
rect 13648 24274 13676 25094
rect 13740 24818 13768 25230
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13636 24268 13688 24274
rect 13636 24210 13688 24216
rect 13280 23866 13308 24210
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 10416 23792 10468 23798
rect 10416 23734 10468 23740
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 10428 23322 10456 23734
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 11072 23186 11100 23598
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 10520 22778 10548 23122
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 11808 22098 11836 23734
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12360 23338 12388 23598
rect 12714 23488 12770 23497
rect 12714 23423 12770 23432
rect 12360 23322 12480 23338
rect 12360 23316 12492 23322
rect 12360 23310 12440 23316
rect 12440 23258 12492 23264
rect 12728 23186 12756 23423
rect 12716 23180 12768 23186
rect 12716 23122 12768 23128
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 12728 22794 12756 23122
rect 12990 22944 13046 22953
rect 12990 22879 13046 22888
rect 12636 22778 12756 22794
rect 13004 22778 13032 22879
rect 12624 22772 12756 22778
rect 12676 22766 12756 22772
rect 12992 22772 13044 22778
rect 12624 22714 12676 22720
rect 12992 22714 13044 22720
rect 12636 22234 12664 22714
rect 13280 22642 13308 23122
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 12808 22092 12860 22098
rect 12808 22034 12860 22040
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 11808 21690 11836 22034
rect 12820 22001 12848 22034
rect 12806 21992 12862 22001
rect 12806 21927 12862 21936
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 12820 21146 12848 21927
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12912 21570 12940 21830
rect 13004 21690 13032 22034
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 12912 21542 13032 21570
rect 13004 21486 13032 21542
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 13004 20942 13032 21422
rect 13084 21072 13136 21078
rect 13084 21014 13136 21020
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 13004 20602 13032 20878
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 13096 20534 13124 21014
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13648 20398 13676 22918
rect 13820 22432 13872 22438
rect 13740 22380 13820 22386
rect 13740 22374 13872 22380
rect 13740 22358 13860 22374
rect 13740 22098 13768 22358
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 14016 22001 14044 26726
rect 14752 26489 14780 26726
rect 14738 26480 14794 26489
rect 14738 26415 14794 26424
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 14096 25424 14148 25430
rect 14096 25366 14148 25372
rect 14108 24614 14136 25366
rect 15120 25362 15148 26182
rect 15304 25838 15332 26862
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 15948 26586 15976 26726
rect 15936 26580 15988 26586
rect 15936 26522 15988 26528
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 15304 25294 15332 25774
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14108 24410 14136 24550
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14476 24070 14504 25230
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 15016 25152 15068 25158
rect 15016 25094 15068 25100
rect 14752 24750 14780 25094
rect 15028 24954 15056 25094
rect 15016 24948 15068 24954
rect 15016 24890 15068 24896
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22438 14320 22918
rect 14384 22642 14412 23462
rect 14476 23050 14504 24006
rect 14752 23594 14780 24686
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15120 24342 15148 24618
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 24410 15700 24550
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 15120 23866 15148 24278
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 14740 23588 14792 23594
rect 14740 23530 14792 23536
rect 15212 23338 15240 24142
rect 15672 23866 15700 24346
rect 15764 24206 15792 26318
rect 15856 25702 15884 26386
rect 15948 25838 15976 26522
rect 16684 26382 16712 27270
rect 17052 26450 17080 27503
rect 17040 26444 17092 26450
rect 17040 26386 17092 26392
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 17052 26042 17080 26386
rect 17224 26308 17276 26314
rect 17224 26250 17276 26256
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 15936 25832 15988 25838
rect 15936 25774 15988 25780
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15856 25362 15884 25638
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 15948 24886 15976 25094
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 16394 24576 16450 24585
rect 16394 24511 16450 24520
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 16408 23866 16436 24511
rect 16488 24404 16540 24410
rect 16592 24392 16620 25094
rect 16540 24364 16620 24392
rect 16488 24346 16540 24352
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 15672 23662 15700 23802
rect 16684 23746 16712 25230
rect 16948 24132 17000 24138
rect 16948 24074 17000 24080
rect 16500 23718 16712 23746
rect 16500 23662 16528 23718
rect 15660 23656 15712 23662
rect 15290 23624 15346 23633
rect 15660 23598 15712 23604
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 15290 23559 15346 23568
rect 15120 23322 15240 23338
rect 15304 23322 15332 23559
rect 16500 23497 16528 23598
rect 16960 23594 16988 24074
rect 16948 23588 17000 23594
rect 16948 23530 17000 23536
rect 16580 23520 16632 23526
rect 16486 23488 16542 23497
rect 16580 23462 16632 23468
rect 16486 23423 16542 23432
rect 15108 23316 15240 23322
rect 15160 23310 15240 23316
rect 15292 23316 15344 23322
rect 15108 23258 15160 23264
rect 15292 23258 15344 23264
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 15016 23044 15068 23050
rect 15016 22986 15068 22992
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14660 22234 14688 22578
rect 15028 22234 15056 22986
rect 15120 22642 15148 23258
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15396 22778 15424 23054
rect 15672 22778 15700 23122
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15672 22234 15700 22714
rect 16040 22642 16068 22986
rect 16396 22976 16448 22982
rect 16394 22944 16396 22953
rect 16592 22964 16620 23462
rect 16448 22944 16620 22964
rect 16450 22936 16620 22944
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16394 22879 16450 22888
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15844 22500 15896 22506
rect 15844 22442 15896 22448
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 14002 21992 14058 22001
rect 14660 21962 14688 22170
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14002 21927 14058 21936
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14292 21486 14320 21898
rect 14752 21690 14780 22034
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15120 21690 15148 21966
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14200 20398 14228 21082
rect 14752 21078 14780 21626
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 14740 21072 14792 21078
rect 14740 21014 14792 21020
rect 15304 20602 15332 21354
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15672 21146 15700 21286
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15856 20602 15884 22442
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 15936 22092 15988 22098
rect 15936 22034 15988 22040
rect 15948 21554 15976 22034
rect 16316 21894 16344 22374
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16316 21690 16344 21830
rect 16684 21690 16712 22918
rect 16960 21690 16988 23530
rect 17236 23050 17264 26250
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17420 24750 17448 25094
rect 17972 24834 18000 33272
rect 18144 33254 18196 33260
rect 18156 33130 18184 33254
rect 18064 33102 18184 33130
rect 18064 31754 18092 33102
rect 18236 32972 18288 32978
rect 18236 32914 18288 32920
rect 18144 32768 18196 32774
rect 18144 32710 18196 32716
rect 18156 32366 18184 32710
rect 18144 32360 18196 32366
rect 18144 32302 18196 32308
rect 18144 32224 18196 32230
rect 18248 32178 18276 32914
rect 18196 32172 18276 32178
rect 18144 32166 18276 32172
rect 18156 32150 18276 32166
rect 18144 31884 18196 31890
rect 18144 31826 18196 31832
rect 18052 31748 18104 31754
rect 18052 31690 18104 31696
rect 18156 31210 18184 31826
rect 18144 31204 18196 31210
rect 18144 31146 18196 31152
rect 18156 30274 18184 31146
rect 18248 30818 18276 32150
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 18248 30790 18368 30818
rect 18340 30734 18368 30790
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18156 30258 18276 30274
rect 18156 30252 18288 30258
rect 18156 30246 18236 30252
rect 18156 29782 18184 30246
rect 18236 30194 18288 30200
rect 18432 30190 18460 31826
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 18144 29776 18196 29782
rect 18144 29718 18196 29724
rect 18432 29306 18460 30126
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 18524 27130 18552 35686
rect 19156 35148 19208 35154
rect 19156 35090 19208 35096
rect 18696 35012 18748 35018
rect 18696 34954 18748 34960
rect 18708 34610 18736 34954
rect 18970 34912 19026 34921
rect 18970 34847 19026 34856
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18880 32360 18932 32366
rect 18880 32302 18932 32308
rect 18892 32026 18920 32302
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 18604 31748 18656 31754
rect 18604 31690 18656 31696
rect 18616 31482 18644 31690
rect 18892 31521 18920 31962
rect 18878 31512 18934 31521
rect 18604 31476 18656 31482
rect 18878 31447 18934 31456
rect 18604 31418 18656 31424
rect 18788 30796 18840 30802
rect 18788 30738 18840 30744
rect 18800 30258 18828 30738
rect 18880 30592 18932 30598
rect 18880 30534 18932 30540
rect 18892 30394 18920 30534
rect 18880 30388 18932 30394
rect 18880 30330 18932 30336
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18800 29850 18828 30194
rect 18788 29844 18840 29850
rect 18788 29786 18840 29792
rect 18892 29617 18920 30330
rect 18878 29608 18934 29617
rect 18878 29543 18934 29552
rect 18892 29102 18920 29543
rect 18880 29096 18932 29102
rect 18880 29038 18932 29044
rect 18984 27402 19012 34847
rect 19168 34785 19196 35090
rect 19154 34776 19210 34785
rect 19154 34711 19156 34720
rect 19208 34711 19210 34720
rect 19156 34682 19208 34688
rect 19156 34604 19208 34610
rect 19156 34546 19208 34552
rect 19168 33862 19196 34546
rect 19156 33856 19208 33862
rect 19156 33798 19208 33804
rect 19168 32298 19196 33798
rect 19444 33674 19472 39520
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 20258 36000 20314 36009
rect 20258 35935 20314 35944
rect 20168 35760 20220 35766
rect 20168 35702 20220 35708
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 20076 34604 20128 34610
rect 20076 34546 20128 34552
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 20088 34241 20116 34546
rect 20180 34474 20208 35702
rect 20272 35290 20300 35935
rect 20260 35284 20312 35290
rect 20260 35226 20312 35232
rect 20272 34542 20300 35226
rect 20548 34785 20576 39520
rect 21178 35864 21234 35873
rect 21178 35799 21234 35808
rect 20904 35488 20956 35494
rect 20904 35430 20956 35436
rect 21088 35488 21140 35494
rect 21088 35430 21140 35436
rect 20916 35290 20944 35430
rect 20994 35320 21050 35329
rect 20904 35284 20956 35290
rect 20994 35255 21050 35264
rect 20904 35226 20956 35232
rect 21008 35154 21036 35255
rect 20996 35148 21048 35154
rect 20996 35090 21048 35096
rect 20904 34944 20956 34950
rect 20904 34886 20956 34892
rect 20534 34776 20590 34785
rect 20534 34711 20590 34720
rect 20536 34672 20588 34678
rect 20536 34614 20588 34620
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20168 34468 20220 34474
rect 20168 34410 20220 34416
rect 20074 34232 20130 34241
rect 20074 34167 20076 34176
rect 20128 34167 20130 34176
rect 20076 34138 20128 34144
rect 20180 34134 20208 34410
rect 20168 34128 20220 34134
rect 20168 34070 20220 34076
rect 19248 33652 19300 33658
rect 19444 33646 19932 33674
rect 19248 33594 19300 33600
rect 19260 33300 19288 33594
rect 19260 33272 19380 33300
rect 19352 33114 19380 33272
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19156 32292 19208 32298
rect 19156 32234 19208 32240
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19444 31657 19472 32166
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19430 31648 19486 31657
rect 19430 31583 19486 31592
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 19064 29572 19116 29578
rect 19064 29514 19116 29520
rect 19076 28694 19104 29514
rect 19168 29238 19196 29990
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19616 29708 19668 29714
rect 19616 29650 19668 29656
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19248 29504 19300 29510
rect 19248 29446 19300 29452
rect 19156 29232 19208 29238
rect 19156 29174 19208 29180
rect 19168 29034 19196 29174
rect 19260 29170 19288 29446
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19248 28756 19300 28762
rect 19352 28744 19380 29582
rect 19628 29306 19656 29650
rect 19616 29300 19668 29306
rect 19616 29242 19668 29248
rect 19628 29050 19656 29242
rect 19300 28716 19380 28744
rect 19444 29022 19656 29050
rect 19248 28698 19300 28704
rect 19064 28688 19116 28694
rect 19064 28630 19116 28636
rect 19444 28082 19472 29022
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19524 28688 19576 28694
rect 19524 28630 19576 28636
rect 19536 28218 19564 28630
rect 19708 28552 19760 28558
rect 19708 28494 19760 28500
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19720 28218 19748 28494
rect 19524 28212 19576 28218
rect 19524 28154 19576 28160
rect 19708 28212 19760 28218
rect 19708 28154 19760 28160
rect 19812 28150 19840 28494
rect 19800 28144 19852 28150
rect 19800 28086 19852 28092
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19904 27577 19932 33646
rect 20168 33448 20220 33454
rect 20168 33390 20220 33396
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 19996 32366 20024 33254
rect 20180 32774 20208 33390
rect 20168 32768 20220 32774
rect 20168 32710 20220 32716
rect 20180 32609 20208 32710
rect 20166 32600 20222 32609
rect 20166 32535 20168 32544
rect 20220 32535 20222 32544
rect 20168 32506 20220 32512
rect 20548 32450 20576 34614
rect 20916 34542 20944 34886
rect 21008 34746 21036 35090
rect 20996 34740 21048 34746
rect 20996 34682 21048 34688
rect 21100 34592 21128 35430
rect 21192 34785 21220 35799
rect 21178 34776 21234 34785
rect 21178 34711 21234 34720
rect 21008 34564 21128 34592
rect 20904 34536 20956 34542
rect 20904 34478 20956 34484
rect 20916 33998 20944 34478
rect 21008 34066 21036 34564
rect 20996 34060 21048 34066
rect 20996 34002 21048 34008
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20904 33992 20956 33998
rect 20904 33934 20956 33940
rect 20640 33454 20668 33934
rect 21008 33658 21036 34002
rect 20996 33652 21048 33658
rect 20996 33594 21048 33600
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 20628 32972 20680 32978
rect 20628 32914 20680 32920
rect 20640 32570 20668 32914
rect 21088 32768 21140 32774
rect 21088 32710 21140 32716
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20548 32422 20668 32450
rect 21100 32434 21128 32710
rect 19984 32360 20036 32366
rect 19984 32302 20036 32308
rect 20640 30841 20668 32422
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 20904 32360 20956 32366
rect 20904 32302 20956 32308
rect 20812 32224 20864 32230
rect 20812 32166 20864 32172
rect 20824 32026 20852 32166
rect 20812 32020 20864 32026
rect 20812 31962 20864 31968
rect 20824 31482 20852 31962
rect 20916 31822 20944 32302
rect 21100 31958 21128 32370
rect 21088 31952 21140 31958
rect 21088 31894 21140 31900
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 20824 31278 20852 31418
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20916 30938 20944 31758
rect 20904 30932 20956 30938
rect 20904 30874 20956 30880
rect 20626 30832 20682 30841
rect 20626 30767 20682 30776
rect 20916 30274 20944 30874
rect 20824 30246 20944 30274
rect 20824 30190 20852 30246
rect 20812 30184 20864 30190
rect 20812 30126 20864 30132
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20536 30048 20588 30054
rect 20536 29990 20588 29996
rect 20088 29170 20116 29990
rect 20548 29850 20576 29990
rect 20536 29844 20588 29850
rect 20536 29786 20588 29792
rect 20548 29646 20576 29786
rect 20824 29714 20852 30126
rect 21192 29866 21220 34711
rect 21652 34082 21680 39520
rect 22756 36258 22784 39520
rect 22664 36230 22784 36258
rect 22836 36304 22888 36310
rect 22836 36246 22888 36252
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 21732 36032 21784 36038
rect 22284 36032 22336 36038
rect 21732 35974 21784 35980
rect 22282 36000 22284 36009
rect 22336 36000 22338 36009
rect 21744 35630 21772 35974
rect 22282 35935 22338 35944
rect 22480 35834 22508 36110
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 21732 35624 21784 35630
rect 21732 35566 21784 35572
rect 21744 34542 21772 35566
rect 22020 35290 22048 35634
rect 22008 35284 22060 35290
rect 22008 35226 22060 35232
rect 22480 35222 22508 35770
rect 22664 35329 22692 36230
rect 22848 35834 22876 36246
rect 22928 36168 22980 36174
rect 22928 36110 22980 36116
rect 22836 35828 22888 35834
rect 22836 35770 22888 35776
rect 22650 35320 22706 35329
rect 22848 35290 22876 35770
rect 22940 35766 22968 36110
rect 22928 35760 22980 35766
rect 22928 35702 22980 35708
rect 22650 35255 22706 35264
rect 22836 35284 22888 35290
rect 22836 35226 22888 35232
rect 22468 35216 22520 35222
rect 22468 35158 22520 35164
rect 22480 34746 22508 35158
rect 22468 34740 22520 34746
rect 22468 34682 22520 34688
rect 21732 34536 21784 34542
rect 21732 34478 21784 34484
rect 22284 34468 22336 34474
rect 22284 34410 22336 34416
rect 22296 34202 22324 34410
rect 22284 34196 22336 34202
rect 22284 34138 22336 34144
rect 21100 29838 21220 29866
rect 21284 34054 21680 34082
rect 22744 34060 22796 34066
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20536 29640 20588 29646
rect 20536 29582 20588 29588
rect 20824 29306 20852 29650
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 20088 28762 20116 29106
rect 20352 29096 20404 29102
rect 20352 29038 20404 29044
rect 20720 29096 20772 29102
rect 20720 29038 20772 29044
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 20364 28422 20392 29038
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20548 28506 20576 28902
rect 20732 28558 20760 29038
rect 20824 28762 20852 29242
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 20720 28552 20772 28558
rect 20548 28478 20668 28506
rect 20720 28494 20772 28500
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20640 28370 20668 28478
rect 20548 28234 20576 28358
rect 20640 28342 20760 28370
rect 19984 28212 20036 28218
rect 20548 28206 20668 28234
rect 19984 28154 20036 28160
rect 19890 27568 19946 27577
rect 19340 27532 19392 27538
rect 19890 27503 19946 27512
rect 19340 27474 19392 27480
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 18972 27396 19024 27402
rect 18972 27338 19024 27344
rect 19076 27130 19104 27406
rect 19352 27130 19380 27474
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19076 26586 19104 27066
rect 19904 26858 19932 27406
rect 19892 26852 19944 26858
rect 19892 26794 19944 26800
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19996 26586 20024 28154
rect 19064 26580 19116 26586
rect 19064 26522 19116 26528
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 19156 26512 19208 26518
rect 19156 26454 19208 26460
rect 20166 26480 20222 26489
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 17880 24818 18000 24834
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17868 24812 18000 24818
rect 17920 24806 18000 24812
rect 17868 24754 17920 24760
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17328 23866 17356 24142
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17420 23730 17448 24686
rect 17512 24206 17540 24754
rect 18156 24682 18184 25298
rect 18340 24954 18368 25774
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18616 24993 18644 25094
rect 18602 24984 18658 24993
rect 18328 24948 18380 24954
rect 18602 24919 18658 24928
rect 18328 24890 18380 24896
rect 18708 24857 18736 25094
rect 18694 24848 18750 24857
rect 18694 24783 18750 24792
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 24410 17816 24550
rect 17776 24404 17828 24410
rect 17776 24346 17828 24352
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17328 22778 17356 23054
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 17328 22234 17356 22714
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15948 21146 15976 21490
rect 16684 21486 16712 21626
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 17328 21350 17356 21966
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 2778 20088 2834 20097
rect 13924 20058 13952 20334
rect 2778 20023 2834 20032
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 13924 19378 13952 19994
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 19378 14596 19790
rect 15304 19394 15332 20538
rect 15948 20466 15976 21082
rect 17328 21010 17356 21286
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16224 20602 16252 20878
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 16040 19990 16068 20266
rect 16224 19990 16252 20538
rect 17328 20534 17356 20946
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16684 20058 16712 20198
rect 16960 20058 16988 20402
rect 17420 20398 17448 23666
rect 17512 23662 17540 24142
rect 17788 23866 17816 24210
rect 18616 24206 18644 24686
rect 18708 24614 18736 24783
rect 18696 24608 18748 24614
rect 18694 24576 18696 24585
rect 18748 24576 18750 24585
rect 18694 24511 18750 24520
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17500 23656 17552 23662
rect 18052 23656 18104 23662
rect 17500 23598 17552 23604
rect 18050 23624 18052 23633
rect 18104 23624 18106 23633
rect 18050 23559 18106 23568
rect 18616 23186 18644 24142
rect 18800 23798 18828 25638
rect 18984 24818 19012 25910
rect 19168 25498 19196 26454
rect 20166 26415 20222 26424
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19720 25770 19748 26318
rect 19708 25764 19760 25770
rect 19708 25706 19760 25712
rect 19248 25696 19300 25702
rect 19300 25644 19380 25650
rect 19248 25638 19380 25644
rect 19260 25622 19380 25638
rect 19156 25492 19208 25498
rect 19156 25434 19208 25440
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18984 24410 19012 24754
rect 18972 24404 19024 24410
rect 18972 24346 19024 24352
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18788 23792 18840 23798
rect 18788 23734 18840 23740
rect 18892 23322 18920 24210
rect 19352 23866 19380 25622
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19616 25356 19668 25362
rect 19616 25298 19668 25304
rect 19628 24682 19656 25298
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19812 24954 19840 25230
rect 19800 24948 19852 24954
rect 19800 24890 19852 24896
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19616 24676 19668 24682
rect 19616 24618 19668 24624
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19904 24342 19932 24686
rect 19996 24410 20024 24686
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19892 24336 19944 24342
rect 19892 24278 19944 24284
rect 19982 24304 20038 24313
rect 19982 24239 20038 24248
rect 19996 23866 20024 24239
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 19444 23254 19472 23598
rect 19996 23594 20024 23802
rect 19984 23588 20036 23594
rect 19984 23530 20036 23536
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 17604 22778 17632 23122
rect 18420 22976 18472 22982
rect 18420 22918 18472 22924
rect 17592 22772 17644 22778
rect 17592 22714 17644 22720
rect 17604 22234 17632 22714
rect 18432 22574 18460 22918
rect 19444 22778 19472 23190
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 18420 22568 18472 22574
rect 18472 22528 18552 22556
rect 18420 22510 18472 22516
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17684 22092 17736 22098
rect 17684 22034 17736 22040
rect 17696 21690 17724 22034
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17696 21146 17724 21626
rect 18064 21486 18092 22374
rect 18524 22234 18552 22528
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17420 20058 17448 20334
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 16212 19984 16264 19990
rect 16212 19926 16264 19932
rect 16040 19514 16068 19926
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 15120 19366 15332 19394
rect 14568 19174 14596 19314
rect 15120 19310 15148 19366
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18970 14596 19110
rect 16040 18970 16068 19450
rect 16224 19174 16252 19926
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 570 6760 626 6769
rect 570 6695 626 6704
rect 584 5681 612 6695
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 17512 5681 17540 20198
rect 17880 20058 17908 20470
rect 17972 20330 18000 20946
rect 18064 20602 18092 21422
rect 18892 21418 18920 21966
rect 19352 21690 19380 22170
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 18880 21412 18932 21418
rect 18880 21354 18932 21360
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17592 19984 17644 19990
rect 17592 19926 17644 19932
rect 17604 19514 17632 19926
rect 18064 19514 18092 20538
rect 18156 20398 18184 21082
rect 19444 20602 19472 21286
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 18144 20392 18196 20398
rect 19536 20369 19564 20470
rect 19904 20398 19932 21354
rect 20180 20942 20208 26415
rect 20640 25838 20668 28206
rect 20732 27010 20760 28342
rect 20824 28014 20852 28698
rect 20812 28008 20864 28014
rect 20812 27950 20864 27956
rect 20824 27674 20852 27950
rect 20812 27668 20864 27674
rect 20812 27610 20864 27616
rect 21100 27402 21128 29838
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 21192 29102 21220 29650
rect 21284 29186 21312 34054
rect 22744 34002 22796 34008
rect 22756 33658 22784 34002
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 21824 33448 21876 33454
rect 21824 33390 21876 33396
rect 21640 31884 21692 31890
rect 21640 31826 21692 31832
rect 21652 31210 21680 31826
rect 21836 31482 21864 33390
rect 21916 33380 21968 33386
rect 21916 33322 21968 33328
rect 21928 33130 21956 33322
rect 21928 33114 22140 33130
rect 21928 33108 22152 33114
rect 21928 33102 22100 33108
rect 22100 33050 22152 33056
rect 22112 32502 22140 33050
rect 22940 32978 22968 35702
rect 23860 35630 23888 39520
rect 24964 37074 24992 39520
rect 24780 37046 24992 37074
rect 24780 36242 24808 37046
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 24216 36032 24268 36038
rect 24216 35974 24268 35980
rect 23848 35624 23900 35630
rect 23754 35592 23810 35601
rect 23848 35566 23900 35572
rect 23754 35527 23810 35536
rect 23572 35488 23624 35494
rect 23572 35430 23624 35436
rect 23480 35284 23532 35290
rect 23480 35226 23532 35232
rect 23492 34134 23520 35226
rect 23584 35018 23612 35430
rect 23572 35012 23624 35018
rect 23572 34954 23624 34960
rect 23584 34241 23612 34954
rect 23570 34232 23626 34241
rect 23570 34167 23572 34176
rect 23624 34167 23626 34176
rect 23572 34138 23624 34144
rect 23480 34128 23532 34134
rect 23480 34070 23532 34076
rect 23492 33658 23520 34070
rect 23480 33652 23532 33658
rect 23480 33594 23532 33600
rect 23584 33522 23612 34138
rect 23572 33516 23624 33522
rect 23572 33458 23624 33464
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 22928 32972 22980 32978
rect 22928 32914 22980 32920
rect 22100 32496 22152 32502
rect 22100 32438 22152 32444
rect 22940 32026 22968 32914
rect 23400 32842 23428 33390
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23388 32836 23440 32842
rect 23388 32778 23440 32784
rect 23296 32360 23348 32366
rect 23296 32302 23348 32308
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 22008 31952 22060 31958
rect 22008 31894 22060 31900
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 22020 31346 22048 31894
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 21640 31204 21692 31210
rect 21640 31146 21692 31152
rect 21652 30938 21680 31146
rect 22020 30938 22048 31282
rect 23308 30938 23336 32302
rect 23388 31884 23440 31890
rect 23492 31872 23520 33254
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23584 32570 23612 32846
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23664 32224 23716 32230
rect 23664 32166 23716 32172
rect 23440 31844 23520 31872
rect 23388 31826 23440 31832
rect 23400 31482 23428 31826
rect 23388 31476 23440 31482
rect 23388 31418 23440 31424
rect 21640 30932 21692 30938
rect 21640 30874 21692 30880
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 21652 30394 21680 30874
rect 22558 30832 22614 30841
rect 22558 30767 22560 30776
rect 22612 30767 22614 30776
rect 22560 30738 22612 30744
rect 22572 30394 22600 30738
rect 23676 30734 23704 32166
rect 23664 30728 23716 30734
rect 23664 30670 23716 30676
rect 21640 30388 21692 30394
rect 21640 30330 21692 30336
rect 22560 30388 22612 30394
rect 22560 30330 22612 30336
rect 23676 30190 23704 30670
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 21548 29232 21600 29238
rect 21284 29158 21404 29186
rect 21548 29174 21600 29180
rect 21180 29096 21232 29102
rect 21180 29038 21232 29044
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 21192 27878 21220 28562
rect 21180 27872 21232 27878
rect 21180 27814 21232 27820
rect 21284 27606 21312 28970
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 20732 26982 20852 27010
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 20732 26586 20760 26794
rect 20720 26580 20772 26586
rect 20720 26522 20772 26528
rect 20720 26444 20772 26450
rect 20720 26386 20772 26392
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20640 25537 20668 25774
rect 20626 25528 20682 25537
rect 20732 25498 20760 26386
rect 20824 26042 20852 26982
rect 21008 26926 21036 27270
rect 21180 27124 21232 27130
rect 21284 27112 21312 27542
rect 21232 27084 21312 27112
rect 21180 27066 21232 27072
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 20904 26376 20956 26382
rect 21008 26330 21036 26862
rect 20956 26324 21036 26330
rect 20904 26318 21036 26324
rect 20916 26302 21036 26318
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20824 25702 20852 25978
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20626 25463 20682 25472
rect 20720 25492 20772 25498
rect 20640 25430 20668 25463
rect 20720 25434 20772 25440
rect 20628 25424 20680 25430
rect 20628 25366 20680 25372
rect 20260 25356 20312 25362
rect 20260 25298 20312 25304
rect 20272 24410 20300 25298
rect 20732 25106 20760 25434
rect 21008 25430 21036 26302
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 21100 25498 21128 25842
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 20996 25424 21048 25430
rect 20996 25366 21048 25372
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 20732 25078 20852 25106
rect 20718 24984 20774 24993
rect 20824 24954 20852 25078
rect 20718 24919 20774 24928
rect 20812 24948 20864 24954
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 20732 24342 20760 24919
rect 20812 24890 20864 24896
rect 20916 24886 20944 25298
rect 20904 24880 20956 24886
rect 20902 24848 20904 24857
rect 20956 24848 20958 24857
rect 21008 24818 21036 25366
rect 20902 24783 20958 24792
rect 20996 24812 21048 24818
rect 20916 24757 20944 24783
rect 20996 24754 21048 24760
rect 20720 24336 20772 24342
rect 20720 24278 20772 24284
rect 20732 23866 20760 24278
rect 21008 24274 21036 24754
rect 21376 24313 21404 29158
rect 21560 25838 21588 29174
rect 21836 28937 21864 29242
rect 21916 29096 21968 29102
rect 21916 29038 21968 29044
rect 21822 28928 21878 28937
rect 21822 28863 21878 28872
rect 21928 28778 21956 29038
rect 23662 28928 23718 28937
rect 23662 28863 23718 28872
rect 21928 28762 22140 28778
rect 23676 28762 23704 28863
rect 21928 28756 22152 28762
rect 21928 28750 22100 28756
rect 22100 28698 22152 28704
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23768 28150 23796 35527
rect 24032 34944 24084 34950
rect 24032 34886 24084 34892
rect 24044 34542 24072 34886
rect 24032 34536 24084 34542
rect 24032 34478 24084 34484
rect 24044 34134 24072 34478
rect 24032 34128 24084 34134
rect 24032 34070 24084 34076
rect 24124 33584 24176 33590
rect 24124 33526 24176 33532
rect 24136 33386 24164 33526
rect 24124 33380 24176 33386
rect 24124 33322 24176 33328
rect 24124 32768 24176 32774
rect 24124 32710 24176 32716
rect 24136 32366 24164 32710
rect 24228 32434 24256 35974
rect 24780 35834 24808 36178
rect 24952 36032 25004 36038
rect 24952 35974 25004 35980
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 24964 35630 24992 35974
rect 24952 35624 25004 35630
rect 24952 35566 25004 35572
rect 24964 35290 24992 35566
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 25044 35284 25096 35290
rect 25044 35226 25096 35232
rect 24950 34776 25006 34785
rect 25056 34746 25084 35226
rect 24950 34711 25006 34720
rect 25044 34740 25096 34746
rect 24676 33516 24728 33522
rect 24676 33458 24728 33464
rect 24688 33114 24716 33458
rect 24676 33108 24728 33114
rect 24676 33050 24728 33056
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24872 33017 24900 33050
rect 24858 33008 24914 33017
rect 24858 32943 24914 32952
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24124 32360 24176 32366
rect 24124 32302 24176 32308
rect 24124 32224 24176 32230
rect 24124 32166 24176 32172
rect 24136 32026 24164 32166
rect 24228 32026 24256 32370
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24216 32020 24268 32026
rect 24216 31962 24268 31968
rect 24228 31822 24256 31962
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 24216 31816 24268 31822
rect 24216 31758 24268 31764
rect 24780 31482 24808 31826
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24768 31476 24820 31482
rect 24768 31418 24820 31424
rect 24766 31240 24822 31249
rect 24688 31184 24766 31192
rect 24688 31164 24768 31184
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23860 29850 23888 29990
rect 23848 29844 23900 29850
rect 23848 29786 23900 29792
rect 23952 29102 23980 30874
rect 24124 30660 24176 30666
rect 24124 30602 24176 30608
rect 24032 30116 24084 30122
rect 24032 30058 24084 30064
rect 24044 29102 24072 30058
rect 24136 29782 24164 30602
rect 24400 30592 24452 30598
rect 24400 30534 24452 30540
rect 24412 30297 24440 30534
rect 24688 30394 24716 31164
rect 24820 31175 24822 31184
rect 24768 31146 24820 31152
rect 24768 30932 24820 30938
rect 24872 30920 24900 31622
rect 24820 30892 24900 30920
rect 24768 30874 24820 30880
rect 24676 30388 24728 30394
rect 24676 30330 24728 30336
rect 24398 30288 24454 30297
rect 24398 30223 24454 30232
rect 24400 30184 24452 30190
rect 24400 30126 24452 30132
rect 24412 29782 24440 30126
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24124 29776 24176 29782
rect 24124 29718 24176 29724
rect 24400 29776 24452 29782
rect 24400 29718 24452 29724
rect 24492 29776 24544 29782
rect 24492 29718 24544 29724
rect 24504 29238 24532 29718
rect 24596 29306 24624 29786
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24780 29345 24808 29446
rect 24766 29336 24822 29345
rect 24584 29300 24636 29306
rect 24766 29271 24822 29280
rect 24584 29242 24636 29248
rect 24216 29232 24268 29238
rect 24216 29174 24268 29180
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 24032 29096 24084 29102
rect 24032 29038 24084 29044
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23860 28218 23888 28494
rect 23848 28212 23900 28218
rect 23848 28154 23900 28160
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23860 28014 23888 28154
rect 23848 28008 23900 28014
rect 23848 27950 23900 27956
rect 21824 27940 21876 27946
rect 21824 27882 21876 27888
rect 21836 27130 21864 27882
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 22112 27470 22140 27814
rect 22836 27532 22888 27538
rect 22836 27474 22888 27480
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 22112 27062 22140 27406
rect 22100 27056 22152 27062
rect 22100 26998 22152 27004
rect 22100 26852 22152 26858
rect 22100 26794 22152 26800
rect 22112 26194 22140 26794
rect 22664 26790 22692 27406
rect 22848 26858 22876 27474
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 23124 27130 23152 27406
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 22836 26852 22888 26858
rect 22836 26794 22888 26800
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 24032 26784 24084 26790
rect 24032 26726 24084 26732
rect 22020 26166 22140 26194
rect 22020 25906 22048 26166
rect 22664 26042 22692 26726
rect 23940 26580 23992 26586
rect 23940 26522 23992 26528
rect 23846 26344 23902 26353
rect 23846 26279 23902 26288
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 21548 25832 21600 25838
rect 21548 25774 21600 25780
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 21560 25498 21588 25774
rect 23676 25537 23704 25774
rect 22006 25528 22062 25537
rect 21548 25492 21600 25498
rect 22006 25463 22062 25472
rect 23662 25528 23718 25537
rect 23662 25463 23664 25472
rect 21548 25434 21600 25440
rect 21362 24304 21418 24313
rect 20996 24268 21048 24274
rect 21362 24239 21418 24248
rect 20996 24210 21048 24216
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 21008 22778 21036 24210
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21376 23798 21404 24142
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21468 23322 21496 24142
rect 22020 23866 22048 25463
rect 23716 25463 23718 25472
rect 23664 25434 23716 25440
rect 23860 25294 23888 26279
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23848 25288 23900 25294
rect 23848 25230 23900 25236
rect 23492 24342 23520 25230
rect 23860 24954 23888 25230
rect 23848 24948 23900 24954
rect 23848 24890 23900 24896
rect 23952 24818 23980 26522
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 23492 23866 23520 24278
rect 24044 24274 24072 26726
rect 24228 26217 24256 29174
rect 24768 28960 24820 28966
rect 24768 28902 24820 28908
rect 24780 28762 24808 28902
rect 24768 28756 24820 28762
rect 24768 28698 24820 28704
rect 24492 27872 24544 27878
rect 24492 27814 24544 27820
rect 24504 27674 24532 27814
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24412 26314 24440 26726
rect 24596 26586 24624 26930
rect 24964 26586 24992 34711
rect 25044 34682 25096 34688
rect 25044 34468 25096 34474
rect 25044 34410 25096 34416
rect 25056 34202 25084 34410
rect 25044 34196 25096 34202
rect 25044 34138 25096 34144
rect 25056 33658 25084 34138
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 25056 32434 25084 32846
rect 25044 32428 25096 32434
rect 25044 32370 25096 32376
rect 25148 31958 25176 35430
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 25332 33658 25360 35022
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25320 33652 25372 33658
rect 25320 33594 25372 33600
rect 25792 33454 25820 34138
rect 25872 33856 25924 33862
rect 25872 33798 25924 33804
rect 25884 33538 25912 33798
rect 25884 33522 26004 33538
rect 25884 33516 26016 33522
rect 25884 33510 25964 33516
rect 25780 33448 25832 33454
rect 25780 33390 25832 33396
rect 25228 32972 25280 32978
rect 25228 32914 25280 32920
rect 25240 32570 25268 32914
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25332 32570 25360 32846
rect 25228 32564 25280 32570
rect 25228 32506 25280 32512
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25240 32026 25268 32506
rect 25884 32434 25912 33510
rect 25964 33458 26016 33464
rect 25872 32428 25924 32434
rect 25872 32370 25924 32376
rect 25884 32026 25912 32370
rect 25228 32020 25280 32026
rect 25228 31962 25280 31968
rect 25872 32020 25924 32026
rect 25872 31962 25924 31968
rect 25136 31952 25188 31958
rect 25136 31894 25188 31900
rect 25226 31920 25282 31929
rect 25148 31482 25176 31894
rect 25226 31855 25228 31864
rect 25280 31855 25282 31864
rect 25228 31826 25280 31832
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 25148 30802 25176 31078
rect 25516 30938 25544 31758
rect 26068 31414 26096 39520
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26252 35698 26280 35974
rect 27264 35737 27292 39520
rect 27250 35728 27306 35737
rect 26240 35692 26292 35698
rect 27250 35663 27306 35672
rect 26240 35634 26292 35640
rect 26148 35148 26200 35154
rect 26148 35090 26200 35096
rect 26160 34746 26188 35090
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 26160 34202 26188 34682
rect 26148 34196 26200 34202
rect 26148 34138 26200 34144
rect 26252 33862 26280 35634
rect 26700 35624 26752 35630
rect 26700 35566 26752 35572
rect 26516 35556 26568 35562
rect 26516 35498 26568 35504
rect 26332 35488 26384 35494
rect 26332 35430 26384 35436
rect 26344 35290 26372 35430
rect 26332 35284 26384 35290
rect 26332 35226 26384 35232
rect 26424 35080 26476 35086
rect 26424 35022 26476 35028
rect 26436 34524 26464 35022
rect 26528 34950 26556 35498
rect 26516 34944 26568 34950
rect 26516 34886 26568 34892
rect 26528 34746 26556 34886
rect 26712 34762 26740 35566
rect 29472 35193 29500 39520
rect 29458 35184 29514 35193
rect 29458 35119 29514 35128
rect 26712 34746 26832 34762
rect 26516 34740 26568 34746
rect 26516 34682 26568 34688
rect 26712 34740 26844 34746
rect 26712 34734 26792 34740
rect 26608 34536 26660 34542
rect 26436 34496 26608 34524
rect 26608 34478 26660 34484
rect 26620 33998 26648 34478
rect 26712 34134 26740 34734
rect 26792 34682 26844 34688
rect 28632 34400 28684 34406
rect 28632 34342 28684 34348
rect 26700 34128 26752 34134
rect 26700 34070 26752 34076
rect 26608 33992 26660 33998
rect 26608 33934 26660 33940
rect 26240 33856 26292 33862
rect 26240 33798 26292 33804
rect 26712 33658 26740 34070
rect 27526 33960 27582 33969
rect 27526 33895 27582 33904
rect 26792 33856 26844 33862
rect 26792 33798 26844 33804
rect 26700 33652 26752 33658
rect 26700 33594 26752 33600
rect 26804 33454 26832 33798
rect 27540 33697 27568 33895
rect 28264 33856 28316 33862
rect 28264 33798 28316 33804
rect 27526 33688 27582 33697
rect 27526 33623 27582 33632
rect 28276 33454 28304 33798
rect 26792 33448 26844 33454
rect 26792 33390 26844 33396
rect 27068 33448 27120 33454
rect 27068 33390 27120 33396
rect 28264 33448 28316 33454
rect 28264 33390 28316 33396
rect 27080 33114 27108 33390
rect 27160 33380 27212 33386
rect 27160 33322 27212 33328
rect 27068 33108 27120 33114
rect 27068 33050 27120 33056
rect 27080 32434 27108 33050
rect 27172 32978 27200 33322
rect 28644 33318 28672 34342
rect 30576 33969 30604 39520
rect 31680 34649 31708 39520
rect 32784 35057 32812 39520
rect 33888 35057 33916 39520
rect 34992 37210 35020 39520
rect 35622 39400 35678 39409
rect 35622 39335 35678 39344
rect 34808 37182 35020 37210
rect 34520 35624 34572 35630
rect 34520 35566 34572 35572
rect 32770 35048 32826 35057
rect 32770 34983 32826 34992
rect 33874 35048 33930 35057
rect 33874 34983 33930 34992
rect 31666 34640 31722 34649
rect 31666 34575 31722 34584
rect 30562 33960 30618 33969
rect 30562 33895 30618 33904
rect 30194 33552 30250 33561
rect 30194 33487 30250 33496
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 28632 33312 28684 33318
rect 28632 33254 28684 33260
rect 28368 33046 28396 33254
rect 27804 33040 27856 33046
rect 27804 32982 27856 32988
rect 28356 33040 28408 33046
rect 28356 32982 28408 32988
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 26884 32360 26936 32366
rect 26884 32302 26936 32308
rect 26240 32292 26292 32298
rect 26240 32234 26292 32240
rect 26252 31482 26280 32234
rect 26700 32224 26752 32230
rect 26700 32166 26752 32172
rect 26712 31958 26740 32166
rect 26896 32026 26924 32302
rect 26884 32020 26936 32026
rect 26884 31962 26936 31968
rect 26700 31952 26752 31958
rect 26700 31894 26752 31900
rect 26712 31482 26740 31894
rect 27172 31890 27200 32914
rect 27816 32570 27844 32982
rect 28644 32978 28672 33254
rect 29366 33008 29422 33017
rect 28632 32972 28684 32978
rect 29366 32943 29368 32952
rect 28632 32914 28684 32920
rect 29420 32943 29422 32952
rect 29368 32914 29420 32920
rect 28540 32768 28592 32774
rect 28540 32710 28592 32716
rect 27804 32564 27856 32570
rect 27804 32506 27856 32512
rect 27816 32366 27844 32506
rect 27804 32360 27856 32366
rect 27804 32302 27856 32308
rect 28552 31958 28580 32710
rect 28644 32570 28672 32914
rect 29380 32570 29408 32914
rect 29552 32768 29604 32774
rect 29552 32710 29604 32716
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 29368 32564 29420 32570
rect 29368 32506 29420 32512
rect 28540 31952 28592 31958
rect 29564 31929 29592 32710
rect 28540 31894 28592 31900
rect 29550 31920 29606 31929
rect 26792 31884 26844 31890
rect 26792 31826 26844 31832
rect 27160 31884 27212 31890
rect 29550 31855 29606 31864
rect 27160 31826 27212 31832
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 26700 31476 26752 31482
rect 26700 31418 26752 31424
rect 26056 31408 26108 31414
rect 26056 31350 26108 31356
rect 26804 31278 26832 31826
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 28460 31278 28488 31622
rect 26608 31272 26660 31278
rect 26608 31214 26660 31220
rect 26792 31272 26844 31278
rect 28448 31272 28500 31278
rect 26792 31214 26844 31220
rect 28170 31240 28226 31249
rect 25504 30932 25556 30938
rect 25504 30874 25556 30880
rect 25136 30796 25188 30802
rect 25136 30738 25188 30744
rect 26516 30796 26568 30802
rect 26516 30738 26568 30744
rect 26528 30394 26556 30738
rect 26620 30598 26648 31214
rect 28448 31214 28500 31220
rect 28170 31175 28226 31184
rect 28184 31142 28212 31175
rect 28172 31136 28224 31142
rect 28172 31078 28224 31084
rect 26608 30592 26660 30598
rect 26608 30534 26660 30540
rect 26516 30388 26568 30394
rect 26516 30330 26568 30336
rect 26148 30048 26200 30054
rect 26620 30002 26648 30534
rect 26974 30288 27030 30297
rect 26974 30223 27030 30232
rect 26988 30190 27016 30223
rect 26976 30184 27028 30190
rect 26976 30126 27028 30132
rect 26148 29990 26200 29996
rect 26160 29646 26188 29990
rect 26528 29974 26648 30002
rect 27160 30048 27212 30054
rect 27160 29990 27212 29996
rect 25136 29640 25188 29646
rect 25136 29582 25188 29588
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 25148 29034 25176 29582
rect 26148 29504 26200 29510
rect 26148 29446 26200 29452
rect 26160 29306 26188 29446
rect 26422 29336 26478 29345
rect 26148 29300 26200 29306
rect 26422 29271 26424 29280
rect 26148 29242 26200 29248
rect 26476 29271 26478 29280
rect 26424 29242 26476 29248
rect 25136 29028 25188 29034
rect 25136 28970 25188 28976
rect 25504 28960 25556 28966
rect 25504 28902 25556 28908
rect 25516 28490 25544 28902
rect 26160 28694 26188 29242
rect 26436 29034 26464 29242
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26148 28688 26200 28694
rect 26148 28630 26200 28636
rect 25596 28620 25648 28626
rect 25596 28562 25648 28568
rect 25504 28484 25556 28490
rect 25504 28426 25556 28432
rect 25412 28008 25464 28014
rect 25516 27962 25544 28426
rect 25608 28422 25636 28562
rect 25596 28416 25648 28422
rect 25596 28358 25648 28364
rect 25464 27956 25544 27962
rect 25412 27950 25544 27956
rect 25424 27934 25544 27950
rect 25412 27600 25464 27606
rect 25412 27542 25464 27548
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 25332 26858 25360 27406
rect 25424 27130 25452 27542
rect 25516 27282 25544 27934
rect 25608 27470 25636 28358
rect 25870 28112 25926 28121
rect 25870 28047 25926 28056
rect 25884 28014 25912 28047
rect 25872 28008 25924 28014
rect 25872 27950 25924 27956
rect 26160 27946 26188 28630
rect 26528 28558 26556 29974
rect 27172 29850 27200 29990
rect 27160 29844 27212 29850
rect 27160 29786 27212 29792
rect 26792 29640 26844 29646
rect 26792 29582 26844 29588
rect 26804 29306 26832 29582
rect 27068 29504 27120 29510
rect 27068 29446 27120 29452
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26884 29232 26936 29238
rect 26884 29174 26936 29180
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 26148 27940 26200 27946
rect 26148 27882 26200 27888
rect 26896 27606 26924 29174
rect 27080 29170 27108 29446
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 27252 28620 27304 28626
rect 27252 28562 27304 28568
rect 29920 28620 29972 28626
rect 29920 28562 29972 28568
rect 27264 28218 27292 28562
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 27252 28212 27304 28218
rect 27252 28154 27304 28160
rect 27908 28121 27936 28358
rect 27894 28112 27950 28121
rect 27894 28047 27950 28056
rect 29840 28014 29868 28494
rect 29932 28218 29960 28562
rect 29920 28212 29972 28218
rect 29920 28154 29972 28160
rect 29828 28008 29880 28014
rect 29828 27950 29880 27956
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 26884 27600 26936 27606
rect 26884 27542 26936 27548
rect 25596 27464 25648 27470
rect 25596 27406 25648 27412
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 25596 27328 25648 27334
rect 25516 27276 25596 27282
rect 25516 27270 25648 27276
rect 25516 27254 25636 27270
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 25424 26926 25452 27066
rect 25608 26926 25636 27254
rect 25412 26920 25464 26926
rect 25412 26862 25464 26868
rect 25596 26920 25648 26926
rect 25596 26862 25648 26868
rect 25320 26852 25372 26858
rect 25320 26794 25372 26800
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 24400 26308 24452 26314
rect 24400 26250 24452 26256
rect 24214 26208 24270 26217
rect 24214 26143 24270 26152
rect 24308 25900 24360 25906
rect 24308 25842 24360 25848
rect 24216 25424 24268 25430
rect 24216 25366 24268 25372
rect 24228 24954 24256 25366
rect 24216 24948 24268 24954
rect 24216 24890 24268 24896
rect 24320 24410 24348 25842
rect 24688 25430 24716 26386
rect 25320 26376 25372 26382
rect 25608 26353 25636 26862
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 25320 26318 25372 26324
rect 25594 26344 25650 26353
rect 24860 26240 24912 26246
rect 24860 26182 24912 26188
rect 24872 25906 24900 26182
rect 25332 26042 25360 26318
rect 25884 26314 25912 26794
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 26056 26784 26108 26790
rect 26056 26726 26108 26732
rect 25976 26450 26004 26726
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 25594 26279 25650 26288
rect 25872 26308 25924 26314
rect 25872 26250 25924 26256
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 25332 25498 25360 25978
rect 25976 25974 26004 26386
rect 26068 26382 26096 26726
rect 26528 26586 26556 27406
rect 26516 26580 26568 26586
rect 26516 26522 26568 26528
rect 26056 26376 26108 26382
rect 26240 26376 26292 26382
rect 26056 26318 26108 26324
rect 26238 26344 26240 26353
rect 26332 26376 26384 26382
rect 26292 26344 26294 26353
rect 26700 26376 26752 26382
rect 26332 26318 26384 26324
rect 26620 26324 26700 26330
rect 26620 26318 26752 26324
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 26238 26279 26294 26288
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 25964 25968 26016 25974
rect 25964 25910 26016 25916
rect 26252 25906 26280 26182
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26238 25528 26294 25537
rect 25320 25492 25372 25498
rect 26344 25514 26372 26318
rect 26620 26302 26740 26318
rect 26620 25702 26648 26302
rect 26988 26217 27016 26318
rect 26974 26208 27030 26217
rect 26974 26143 27030 26152
rect 26988 25770 27016 26143
rect 27080 25906 27108 27814
rect 29840 27606 29868 27950
rect 29828 27600 29880 27606
rect 29828 27542 29880 27548
rect 29460 27532 29512 27538
rect 29460 27474 29512 27480
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27816 27130 27844 27270
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27712 26920 27764 26926
rect 27712 26862 27764 26868
rect 29472 26908 29500 27474
rect 29552 26920 29604 26926
rect 29472 26880 29552 26908
rect 27528 26444 27580 26450
rect 27528 26386 27580 26392
rect 27540 26330 27568 26386
rect 27540 26302 27660 26330
rect 27252 26240 27304 26246
rect 27252 26182 27304 26188
rect 27068 25900 27120 25906
rect 27068 25842 27120 25848
rect 27264 25838 27292 26182
rect 27632 26042 27660 26302
rect 27620 26036 27672 26042
rect 27620 25978 27672 25984
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27252 25832 27304 25838
rect 27252 25774 27304 25780
rect 26976 25764 27028 25770
rect 26976 25706 27028 25712
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26294 25486 26372 25514
rect 26238 25463 26240 25472
rect 25320 25434 25372 25440
rect 26292 25463 26294 25472
rect 26240 25434 26292 25440
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24860 25152 24912 25158
rect 24780 25100 24860 25106
rect 26620 25129 26648 25638
rect 26988 25430 27016 25706
rect 27264 25498 27292 25774
rect 27540 25498 27568 25842
rect 27252 25492 27304 25498
rect 27252 25434 27304 25440
rect 27528 25492 27580 25498
rect 27528 25434 27580 25440
rect 26976 25424 27028 25430
rect 26976 25366 27028 25372
rect 24780 25094 24912 25100
rect 26606 25120 26662 25129
rect 24780 25078 24900 25094
rect 24780 24750 24808 25078
rect 26606 25055 26662 25064
rect 25042 24848 25098 24857
rect 25042 24783 25098 24792
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24584 24676 24636 24682
rect 24584 24618 24636 24624
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 24044 23730 24072 24210
rect 24216 24200 24268 24206
rect 24216 24142 24268 24148
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 21548 23588 21600 23594
rect 21548 23530 21600 23536
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21560 22982 21588 23530
rect 24228 22982 24256 24142
rect 24596 23866 24624 24618
rect 24584 23860 24636 23866
rect 24636 23820 24716 23848
rect 24584 23802 24636 23808
rect 24688 23186 24716 23820
rect 25056 23594 25084 24783
rect 25872 24608 25924 24614
rect 27724 24562 27752 26862
rect 29000 26444 29052 26450
rect 29000 26386 29052 26392
rect 28446 26344 28502 26353
rect 28446 26279 28502 26288
rect 28816 26308 28868 26314
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 27816 24993 27844 25094
rect 27802 24984 27858 24993
rect 27802 24919 27858 24928
rect 28184 24614 28212 25298
rect 28460 25294 28488 26279
rect 28816 26250 28868 26256
rect 28828 25922 28856 26250
rect 29012 26042 29040 26386
rect 29472 26382 29500 26880
rect 29552 26862 29604 26868
rect 29460 26376 29512 26382
rect 29460 26318 29512 26324
rect 29000 26036 29052 26042
rect 29000 25978 29052 25984
rect 28828 25894 29132 25922
rect 29472 25906 29500 26318
rect 28816 25356 28868 25362
rect 28816 25298 28868 25304
rect 29000 25356 29052 25362
rect 29000 25298 29052 25304
rect 28448 25288 28500 25294
rect 28448 25230 28500 25236
rect 28460 24954 28488 25230
rect 28722 25120 28778 25129
rect 28722 25055 28778 25064
rect 28448 24948 28500 24954
rect 28448 24890 28500 24896
rect 25872 24550 25924 24556
rect 25884 24206 25912 24550
rect 27540 24534 27752 24562
rect 28172 24608 28224 24614
rect 28172 24550 28224 24556
rect 27540 24410 27568 24534
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27436 24268 27488 24274
rect 27436 24210 27488 24216
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25148 23662 25176 24006
rect 27448 23866 27476 24210
rect 27436 23860 27488 23866
rect 27436 23802 27488 23808
rect 27540 23798 27568 24346
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 27528 23792 27580 23798
rect 27528 23734 27580 23740
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25044 23588 25096 23594
rect 25044 23530 25096 23536
rect 24860 23520 24912 23526
rect 24780 23468 24860 23474
rect 24780 23462 24912 23468
rect 24780 23446 24900 23462
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 21548 22976 21600 22982
rect 21548 22918 21600 22924
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 21560 22817 21588 22918
rect 21546 22808 21602 22817
rect 20996 22772 21048 22778
rect 21546 22743 21602 22752
rect 20996 22714 21048 22720
rect 22112 22574 22140 22918
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 20364 22234 20392 22374
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 21008 21978 21036 22034
rect 20916 21950 21036 21978
rect 20916 21350 20944 21950
rect 21272 21888 21324 21894
rect 21640 21888 21692 21894
rect 21324 21836 21404 21842
rect 21272 21830 21404 21836
rect 21640 21830 21692 21836
rect 21284 21814 21404 21830
rect 21376 21486 21404 21814
rect 21652 21486 21680 21830
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20180 20777 20208 20878
rect 20166 20768 20222 20777
rect 20166 20703 20222 20712
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19892 20392 19944 20398
rect 18144 20334 18196 20340
rect 19522 20360 19578 20369
rect 19892 20334 19944 20340
rect 19522 20295 19578 20304
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19904 19990 19932 20334
rect 19996 20262 20024 20538
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19996 20058 20024 20198
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 20088 19802 20116 20402
rect 20364 20398 20392 20878
rect 20916 20602 20944 21286
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 19996 19774 20116 19802
rect 19996 19718 20024 19774
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 19892 19236 19944 19242
rect 19892 19178 19944 19184
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19904 18902 19932 19178
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19260 18329 19288 18566
rect 19352 18426 19380 18838
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 19628 18426 19656 18770
rect 19996 18766 20024 19654
rect 20364 19514 20392 20334
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 19718 20576 20198
rect 21192 20058 21220 20946
rect 21376 20942 21404 21422
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21376 20097 21404 20742
rect 21362 20088 21418 20097
rect 21180 20052 21232 20058
rect 21362 20023 21418 20032
rect 22020 20040 22048 22374
rect 22112 22166 22140 22510
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22756 21690 22784 22374
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 23124 21690 23152 21830
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 22756 21078 22784 21626
rect 22744 21072 22796 21078
rect 22744 21014 22796 21020
rect 22756 20602 22784 21014
rect 23124 21010 23152 21626
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22190 20360 22246 20369
rect 23124 20330 23152 20946
rect 23400 20346 23428 22578
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23768 21690 23796 22034
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23768 21146 23796 21626
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23860 21026 23888 21286
rect 23768 20998 23888 21026
rect 23664 20392 23716 20398
rect 22190 20295 22246 20304
rect 23112 20324 23164 20330
rect 22020 20012 22140 20040
rect 21180 19994 21232 20000
rect 22112 19922 22140 20012
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22204 19854 22232 20295
rect 23400 20318 23612 20346
rect 23664 20334 23716 20340
rect 23112 20266 23164 20272
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23492 19938 23520 20198
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 23308 19910 23520 19938
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20548 19174 20576 19654
rect 22204 19514 22232 19790
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18834 20576 19110
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19246 18320 19302 18329
rect 19246 18255 19302 18264
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 16998 18644 18022
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 18984 17338 19012 17750
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19260 17241 19288 17478
rect 19246 17232 19302 17241
rect 19246 17167 19302 17176
rect 19246 17096 19302 17105
rect 19628 17066 19656 17614
rect 19904 17542 19932 18158
rect 19996 17678 20024 18702
rect 20074 18184 20130 18193
rect 20074 18119 20076 18128
rect 20128 18119 20130 18128
rect 20076 18090 20128 18096
rect 20350 18048 20406 18057
rect 20350 17983 20406 17992
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19904 17066 19932 17478
rect 19246 17031 19302 17040
rect 19616 17060 19668 17066
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18616 15910 18644 16934
rect 19260 16794 19288 17031
rect 19616 17002 19668 17008
rect 19892 17060 19944 17066
rect 19892 17002 19944 17008
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19904 16726 19932 17002
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19352 16250 19380 16526
rect 19628 16250 19656 16594
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 19352 15638 19380 16186
rect 19904 16046 19932 16662
rect 19996 16590 20024 17614
rect 20364 17134 20392 17983
rect 20916 17678 20944 18702
rect 21192 18426 21220 19178
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21086 18184 21142 18193
rect 21086 18119 21142 18128
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 21100 17338 21128 18119
rect 21560 18086 21588 18770
rect 22020 18426 22048 19246
rect 22296 18970 22324 19858
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22572 19378 22600 19790
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20272 16697 20300 16934
rect 20364 16794 20392 17070
rect 21376 16998 21404 17750
rect 21560 17377 21588 18022
rect 21546 17368 21602 17377
rect 21546 17303 21602 17312
rect 21730 17096 21786 17105
rect 21730 17031 21732 17040
rect 21784 17031 21786 17040
rect 21732 17002 21784 17008
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20258 16688 20314 16697
rect 20258 16623 20314 16632
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19996 15910 20024 16526
rect 20272 16046 20300 16623
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20824 16130 20852 16390
rect 21376 16250 21404 16934
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 20824 16114 21036 16130
rect 20824 16108 21048 16114
rect 20824 16102 20996 16108
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 20272 15706 20300 15982
rect 20824 15978 20852 16102
rect 20996 16050 21048 16056
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 20824 15502 20852 15914
rect 21744 15910 21772 16594
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 15706 21772 15846
rect 22112 15722 22140 18566
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22296 18057 22324 18362
rect 22374 18320 22430 18329
rect 22480 18290 22508 18634
rect 22572 18290 22600 19314
rect 23308 19174 23336 19910
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 22374 18255 22430 18264
rect 22468 18284 22520 18290
rect 22388 18222 22416 18255
rect 22468 18226 22520 18232
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22282 18048 22338 18057
rect 22282 17983 22338 17992
rect 22296 17882 22324 17983
rect 22388 17882 22416 18158
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22572 17746 22600 18226
rect 23400 17882 23428 18906
rect 23584 18850 23612 20318
rect 23676 20097 23704 20334
rect 23768 20262 23796 20998
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23662 20088 23718 20097
rect 23662 20023 23664 20032
rect 23716 20023 23718 20032
rect 23664 19994 23716 20000
rect 23768 19281 23796 20198
rect 23754 19272 23810 19281
rect 23754 19207 23810 19216
rect 23584 18822 23704 18850
rect 23676 18766 23704 18822
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23584 18426 23612 18702
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23676 18154 23704 18702
rect 23860 18222 23888 18770
rect 23848 18216 23900 18222
rect 23846 18184 23848 18193
rect 23900 18184 23902 18193
rect 23664 18148 23716 18154
rect 23846 18119 23902 18128
rect 23664 18090 23716 18096
rect 23676 17882 23704 18090
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 22282 17232 22338 17241
rect 22572 17202 22600 17682
rect 23124 17270 23152 17682
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 22282 17167 22338 17176
rect 22560 17196 22612 17202
rect 22296 17134 22324 17167
rect 22560 17138 22612 17144
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22572 16794 22600 17138
rect 23124 16794 23152 17206
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 23860 16794 23888 17070
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 22296 16697 22324 16730
rect 22282 16688 22338 16697
rect 22282 16623 22338 16632
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22204 15910 22232 16050
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 22020 15694 22140 15722
rect 22020 15638 22048 15694
rect 20904 15632 20956 15638
rect 20904 15574 20956 15580
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20824 15094 20852 15438
rect 20916 15162 20944 15574
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 22100 14816 22152 14822
rect 23480 14816 23532 14822
rect 22100 14758 22152 14764
rect 23294 14784 23350 14793
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 13938 21404 14214
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20916 12918 20944 13330
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 20904 12912 20956 12918
rect 21192 12889 21220 13126
rect 21284 12918 21312 13738
rect 21272 12912 21324 12918
rect 20904 12854 20956 12860
rect 21178 12880 21234 12889
rect 21272 12854 21324 12860
rect 21376 12850 21404 13874
rect 21640 13796 21692 13802
rect 21640 13738 21692 13744
rect 21652 13530 21680 13738
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21744 12986 21772 13262
rect 22020 12986 22048 13466
rect 22112 13326 22140 14758
rect 23480 14758 23532 14764
rect 23294 14719 23350 14728
rect 23308 14618 23336 14719
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 23124 13870 23152 14418
rect 23492 14074 23520 14758
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23676 13870 23704 14418
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 23032 13394 23060 13670
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 21178 12815 21234 12824
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 22204 12782 22232 13126
rect 23032 12986 23060 13330
rect 23492 12986 23520 13738
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 21468 12442 21496 12650
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22112 11898 22140 12242
rect 22204 12102 22232 12718
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22204 11558 22232 12038
rect 23676 11898 23704 12718
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23400 11626 23428 11834
rect 23860 11694 23888 12378
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 22204 11150 22232 11494
rect 23400 11354 23428 11562
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22204 10606 22232 11086
rect 22296 10810 22324 11154
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 22296 10266 22324 10746
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22756 10130 22784 10542
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22756 9654 22784 10066
rect 22848 9722 22876 10066
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 23768 9518 23796 10542
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 23768 9042 23796 9454
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 570 5672 626 5681
rect 570 5607 626 5616
rect 17498 5672 17554 5681
rect 17498 5607 17554 5616
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 23952 4049 23980 22374
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 24044 20058 24072 21082
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 24044 19174 24072 19790
rect 24228 19417 24256 22918
rect 24490 22536 24546 22545
rect 24490 22471 24546 22480
rect 24504 21554 24532 22471
rect 24688 21894 24716 23122
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24780 21690 24808 23446
rect 25148 23254 25176 23598
rect 26148 23588 26200 23594
rect 26148 23530 26200 23536
rect 25596 23520 25648 23526
rect 25596 23462 25648 23468
rect 25136 23248 25188 23254
rect 25136 23190 25188 23196
rect 25148 22778 25176 23190
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25148 22234 25176 22714
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24674 21584 24730 21593
rect 24492 21548 24544 21554
rect 24674 21519 24676 21528
rect 24492 21490 24544 21496
rect 24728 21519 24730 21528
rect 24676 21490 24728 21496
rect 24504 21146 24532 21490
rect 24492 21140 24544 21146
rect 24492 21082 24544 21088
rect 24688 21010 24716 21490
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 25148 20942 25176 21286
rect 25240 21146 25268 22374
rect 25504 21888 25556 21894
rect 25504 21830 25556 21836
rect 25516 21486 25544 21830
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25608 21146 25636 23462
rect 25872 22976 25924 22982
rect 25872 22918 25924 22924
rect 25686 22808 25742 22817
rect 25686 22743 25688 22752
rect 25740 22743 25742 22752
rect 25688 22714 25740 22720
rect 25228 21140 25280 21146
rect 25228 21082 25280 21088
rect 25596 21140 25648 21146
rect 25596 21082 25648 21088
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 24306 20496 24362 20505
rect 24306 20431 24308 20440
rect 24360 20431 24362 20440
rect 24308 20402 24360 20408
rect 24320 19990 24348 20402
rect 25148 20058 25176 20878
rect 25240 20602 25268 21082
rect 25608 20602 25636 21082
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 24308 19984 24360 19990
rect 24308 19926 24360 19932
rect 24400 19916 24452 19922
rect 24400 19858 24452 19864
rect 24214 19408 24270 19417
rect 24214 19343 24270 19352
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 24044 19009 24072 19110
rect 24030 19000 24086 19009
rect 24030 18935 24086 18944
rect 24136 14278 24164 19246
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 24228 18358 24256 19110
rect 24412 18970 24440 19858
rect 24490 19408 24546 19417
rect 24546 19366 24624 19394
rect 24490 19343 24546 19352
rect 24596 19310 24624 19366
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 24400 18148 24452 18154
rect 24400 18090 24452 18096
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24320 16794 24348 17682
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24320 15910 24348 16730
rect 24412 16590 24440 18090
rect 24504 16794 24532 19110
rect 24688 18970 24716 19110
rect 25700 18970 25728 22714
rect 25884 21418 25912 22918
rect 26160 22114 26188 23530
rect 28092 23322 28120 23802
rect 28080 23316 28132 23322
rect 28080 23258 28132 23264
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 26884 22568 26936 22574
rect 26882 22536 26884 22545
rect 26936 22536 26938 22545
rect 26882 22471 26938 22480
rect 27816 22438 27844 23122
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27620 22160 27672 22166
rect 26160 22098 26280 22114
rect 27620 22102 27672 22108
rect 26160 22092 26292 22098
rect 26160 22086 26240 22092
rect 26240 22034 26292 22040
rect 26516 22092 26568 22098
rect 26516 22034 26568 22040
rect 26252 22003 26280 22034
rect 26528 21690 26556 22034
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 26516 21684 26568 21690
rect 26516 21626 26568 21632
rect 26712 21593 26740 21830
rect 26698 21584 26754 21593
rect 26698 21519 26754 21528
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 25872 21412 25924 21418
rect 25872 21354 25924 21360
rect 26804 20942 26832 21422
rect 27068 21344 27120 21350
rect 27068 21286 27120 21292
rect 27080 21010 27108 21286
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 26252 20466 26280 20742
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26056 20256 26108 20262
rect 26054 20224 26056 20233
rect 26108 20224 26110 20233
rect 26054 20159 26110 20168
rect 26620 20058 26648 20402
rect 26608 20052 26660 20058
rect 26608 19994 26660 20000
rect 26514 19952 26570 19961
rect 26514 19887 26516 19896
rect 26568 19887 26570 19896
rect 26516 19858 26568 19864
rect 26240 19712 26292 19718
rect 26160 19660 26240 19666
rect 26160 19654 26292 19660
rect 26160 19638 26280 19654
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25792 19174 25820 19246
rect 25780 19168 25832 19174
rect 25778 19136 25780 19145
rect 25832 19136 25834 19145
rect 25778 19071 25834 19080
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25148 18170 25176 18770
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25240 18426 25268 18702
rect 25228 18420 25280 18426
rect 25228 18362 25280 18368
rect 25700 18222 25728 18906
rect 26160 18766 26188 19638
rect 26528 19514 26556 19858
rect 26804 19854 26832 20878
rect 27080 20466 27108 20946
rect 27632 20754 27660 22102
rect 27540 20726 27660 20754
rect 27710 20768 27766 20777
rect 27540 20466 27568 20726
rect 27710 20703 27766 20712
rect 27618 20632 27674 20641
rect 27618 20567 27620 20576
rect 27672 20567 27674 20576
rect 27620 20538 27672 20544
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26884 19304 26936 19310
rect 26882 19272 26884 19281
rect 26936 19272 26938 19281
rect 26882 19207 26938 19216
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 27080 19009 27108 19110
rect 26698 19000 26754 19009
rect 26698 18935 26700 18944
rect 26752 18935 26754 18944
rect 27066 19000 27122 19009
rect 27066 18935 27122 18944
rect 26700 18906 26752 18912
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 25688 18216 25740 18222
rect 25148 18142 25268 18170
rect 25688 18158 25740 18164
rect 25240 18086 25268 18142
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 17921 25268 18022
rect 25226 17912 25282 17921
rect 25226 17847 25282 17856
rect 25240 17814 25268 17847
rect 26252 17814 26280 18362
rect 26528 18358 26556 18770
rect 27632 18766 27660 19790
rect 27724 18834 27752 20703
rect 27816 18970 27844 22374
rect 28446 21992 28502 22001
rect 28446 21927 28502 21936
rect 28460 21690 28488 21927
rect 28632 21888 28684 21894
rect 28632 21830 28684 21836
rect 28448 21684 28500 21690
rect 28448 21626 28500 21632
rect 28460 21486 28488 21626
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27908 19922 27936 20742
rect 28000 20505 28028 21286
rect 28644 21146 28672 21830
rect 28632 21140 28684 21146
rect 28632 21082 28684 21088
rect 28736 20602 28764 25055
rect 28828 24682 28856 25298
rect 29012 24954 29040 25298
rect 29000 24948 29052 24954
rect 29000 24890 29052 24896
rect 29012 24818 29040 24890
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 28816 24676 28868 24682
rect 28816 24618 28868 24624
rect 28828 23798 28856 24618
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 28906 24032 28962 24041
rect 28906 23967 28962 23976
rect 28920 23866 28948 23967
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 28816 23792 28868 23798
rect 29012 23746 29040 24142
rect 28816 23734 28868 23740
rect 28920 23718 29040 23746
rect 28920 23526 28948 23718
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28920 23118 28948 23462
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28828 21690 28856 21966
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 28920 21486 28948 23054
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 27986 20496 28042 20505
rect 27986 20431 28042 20440
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 28172 20324 28224 20330
rect 28172 20266 28224 20272
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 28092 19990 28120 20198
rect 28080 19984 28132 19990
rect 28080 19926 28132 19932
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 27908 19514 27936 19858
rect 27896 19508 27948 19514
rect 27896 19450 27948 19456
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 27712 18828 27764 18834
rect 27712 18770 27764 18776
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27724 18426 27752 18770
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 26516 18352 26568 18358
rect 26516 18294 26568 18300
rect 25228 17808 25280 17814
rect 25228 17750 25280 17756
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 26700 17808 26752 17814
rect 26700 17750 26752 17756
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24872 17066 24900 17478
rect 25226 17368 25282 17377
rect 26712 17338 26740 17750
rect 27068 17740 27120 17746
rect 27068 17682 27120 17688
rect 25226 17303 25228 17312
rect 25280 17303 25282 17312
rect 26700 17332 26752 17338
rect 25228 17274 25280 17280
rect 26700 17274 26752 17280
rect 24860 17060 24912 17066
rect 24860 17002 24912 17008
rect 24872 16794 24900 17002
rect 24492 16788 24544 16794
rect 24492 16730 24544 16736
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24872 16640 24900 16730
rect 25240 16726 25268 17274
rect 25964 17128 26016 17134
rect 25502 17096 25558 17105
rect 25964 17070 26016 17076
rect 25502 17031 25504 17040
rect 25556 17031 25558 17040
rect 25504 17002 25556 17008
rect 25516 16794 25544 17002
rect 25976 16794 26004 17070
rect 27080 16998 27108 17682
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 27434 16960 27490 16969
rect 27080 16794 27108 16934
rect 27434 16895 27490 16904
rect 27448 16794 27476 16895
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 27068 16788 27120 16794
rect 27068 16730 27120 16736
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 24780 16612 24900 16640
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24412 16250 24440 16526
rect 24780 16250 24808 16612
rect 25240 16250 25268 16662
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24320 15706 24348 15846
rect 24872 15706 24900 15982
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25688 15904 25740 15910
rect 25688 15846 25740 15852
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24228 14618 24256 14758
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24228 14090 24256 14554
rect 24320 14482 24348 15642
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24228 14074 24348 14090
rect 24228 14068 24360 14074
rect 24228 14062 24308 14068
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24136 13530 24164 13738
rect 24228 13530 24256 14062
rect 24308 14010 24360 14016
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24030 12880 24086 12889
rect 24030 12815 24086 12824
rect 24044 12646 24072 12815
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 24044 12442 24072 12582
rect 24228 12442 24256 12650
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24228 11286 24256 11698
rect 24320 11354 24348 12106
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24228 8974 24256 11222
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24228 8090 24256 8910
rect 24412 8566 24440 14214
rect 24688 13512 24716 15506
rect 25424 15502 25452 15846
rect 25700 15706 25728 15846
rect 25688 15700 25740 15706
rect 25688 15642 25740 15648
rect 25976 15638 26004 16730
rect 27080 16046 27108 16730
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26700 15700 26752 15706
rect 26700 15642 26752 15648
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 25872 15564 25924 15570
rect 25872 15506 25924 15512
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 24964 15162 24992 15438
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25332 14550 25360 14962
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25424 14074 25452 14894
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25608 14618 25636 14826
rect 25596 14612 25648 14618
rect 25596 14554 25648 14560
rect 25608 14074 25636 14554
rect 25884 14074 25912 15506
rect 25976 14958 26004 15574
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 25134 13696 25190 13705
rect 25134 13631 25190 13640
rect 24860 13524 24912 13530
rect 24688 13484 24860 13512
rect 24860 13466 24912 13472
rect 24766 13016 24822 13025
rect 24766 12951 24768 12960
rect 24820 12951 24822 12960
rect 24768 12922 24820 12928
rect 24872 12850 24900 13466
rect 25148 13394 25176 13631
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25148 12986 25176 13330
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24504 11558 24532 12174
rect 24596 11898 24624 12242
rect 24688 12220 24716 12786
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25240 12442 25268 12718
rect 25332 12714 25360 13330
rect 25424 13326 25452 14010
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 26160 13025 26188 15438
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26252 13734 26280 14758
rect 26712 14618 26740 15642
rect 26804 14822 26832 15846
rect 27540 15688 27568 16594
rect 27710 15872 27766 15881
rect 27710 15807 27766 15816
rect 27620 15700 27672 15706
rect 27540 15660 27620 15688
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 27080 14822 27108 15574
rect 26792 14816 26844 14822
rect 27068 14816 27120 14822
rect 26792 14758 26844 14764
rect 27066 14784 27068 14793
rect 27120 14784 27122 14793
rect 27066 14719 27122 14728
rect 27540 14618 27568 15660
rect 27620 15642 27672 15648
rect 27724 15502 27752 15807
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27724 15162 27752 15438
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 27528 14612 27580 14618
rect 27528 14554 27580 14560
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26436 13938 26464 14486
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26252 13462 26280 13670
rect 27172 13530 27200 14418
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27540 14074 27568 14350
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 26146 13016 26202 13025
rect 26146 12951 26202 12960
rect 26160 12918 26188 12951
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 27264 12850 27292 13126
rect 27448 12986 27476 13806
rect 27632 13138 27660 14758
rect 27724 14414 27752 15098
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27724 14074 27752 14350
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 27816 13938 27844 18906
rect 27908 18698 27936 19450
rect 28092 18970 28120 19926
rect 28184 19378 28212 20266
rect 29012 20097 29040 20334
rect 28998 20088 29054 20097
rect 28998 20023 29000 20032
rect 29052 20023 29054 20032
rect 29000 19994 29052 20000
rect 28172 19372 28224 19378
rect 28172 19314 28224 19320
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27908 18426 27936 18634
rect 27896 18420 27948 18426
rect 27896 18362 27948 18368
rect 28644 18290 28672 19110
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 27894 17912 27950 17921
rect 27894 17847 27896 17856
rect 27948 17847 27950 17856
rect 27896 17818 27948 17824
rect 28722 17640 28778 17649
rect 28722 17575 28778 17584
rect 28736 17338 28764 17575
rect 28724 17332 28776 17338
rect 28724 17274 28776 17280
rect 28172 17128 28224 17134
rect 28172 17070 28224 17076
rect 28184 16726 28212 17070
rect 28736 17066 28764 17274
rect 28908 17128 28960 17134
rect 28908 17070 28960 17076
rect 28724 17060 28776 17066
rect 28724 17002 28776 17008
rect 28172 16720 28224 16726
rect 28172 16662 28224 16668
rect 28184 16250 28212 16662
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28630 15736 28686 15745
rect 28630 15671 28686 15680
rect 28724 15700 28776 15706
rect 28644 15638 28672 15671
rect 28724 15642 28776 15648
rect 28632 15632 28684 15638
rect 28632 15574 28684 15580
rect 28644 15434 28672 15574
rect 28632 15428 28684 15434
rect 28632 15370 28684 15376
rect 28446 15192 28502 15201
rect 28446 15127 28448 15136
rect 28500 15127 28502 15136
rect 28448 15098 28500 15104
rect 28460 14958 28488 15098
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28644 14618 28672 15370
rect 28736 15162 28764 15642
rect 28816 15360 28868 15366
rect 28816 15302 28868 15308
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 28828 14550 28856 15302
rect 28920 15042 28948 17070
rect 29000 16992 29052 16998
rect 28998 16960 29000 16969
rect 29052 16960 29054 16969
rect 28998 16895 29054 16904
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 29012 16046 29040 16594
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 29012 15162 29040 15438
rect 29104 15178 29132 25894
rect 29460 25900 29512 25906
rect 29460 25842 29512 25848
rect 29472 25498 29500 25842
rect 29460 25492 29512 25498
rect 29380 25452 29460 25480
rect 29380 25294 29408 25452
rect 29460 25434 29512 25440
rect 29368 25288 29420 25294
rect 29368 25230 29420 25236
rect 29380 24750 29408 25230
rect 29368 24744 29420 24750
rect 29368 24686 29420 24692
rect 29380 24410 29408 24686
rect 29368 24404 29420 24410
rect 29368 24346 29420 24352
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 29564 23866 29592 24210
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29184 23180 29236 23186
rect 29184 23122 29236 23128
rect 29196 22574 29224 23122
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 29196 22030 29224 22510
rect 30012 22500 30064 22506
rect 30012 22442 30064 22448
rect 29276 22432 29328 22438
rect 29276 22374 29328 22380
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29288 22234 29316 22374
rect 29276 22228 29328 22234
rect 29276 22170 29328 22176
rect 29748 22098 29776 22374
rect 29460 22092 29512 22098
rect 29460 22034 29512 22040
rect 29736 22092 29788 22098
rect 29736 22034 29788 22040
rect 29184 22024 29236 22030
rect 29184 21966 29236 21972
rect 29196 21690 29224 21966
rect 29184 21684 29236 21690
rect 29184 21626 29236 21632
rect 29196 21078 29224 21626
rect 29184 21072 29236 21078
rect 29184 21014 29236 21020
rect 29276 20596 29328 20602
rect 29276 20538 29328 20544
rect 29288 20398 29316 20538
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29288 19310 29316 20334
rect 29380 19718 29408 20334
rect 29472 20233 29500 22034
rect 29828 21412 29880 21418
rect 29828 21354 29880 21360
rect 29736 21140 29788 21146
rect 29736 21082 29788 21088
rect 29748 20466 29776 21082
rect 29840 20806 29868 21354
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29736 20256 29788 20262
rect 29458 20224 29514 20233
rect 29736 20198 29788 20204
rect 29458 20159 29514 20168
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29380 19553 29408 19654
rect 29366 19544 29422 19553
rect 29366 19479 29422 19488
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29184 19236 29236 19242
rect 29184 19178 29236 19184
rect 29196 18970 29224 19178
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 29196 18426 29224 18906
rect 29472 18902 29500 20159
rect 29748 19378 29776 20198
rect 29840 19922 29868 20742
rect 30024 20398 30052 22442
rect 30116 21894 30144 22578
rect 30104 21888 30156 21894
rect 30104 21830 30156 21836
rect 30116 21486 30144 21830
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 30116 21146 30144 21422
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30012 20392 30064 20398
rect 30012 20334 30064 20340
rect 30102 20224 30158 20233
rect 30102 20159 30158 20168
rect 30116 19990 30144 20159
rect 30104 19984 30156 19990
rect 30104 19926 30156 19932
rect 29828 19916 29880 19922
rect 29828 19858 29880 19864
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 29918 19000 29974 19009
rect 29918 18935 29920 18944
rect 29972 18935 29974 18944
rect 29920 18906 29972 18912
rect 29460 18896 29512 18902
rect 29460 18838 29512 18844
rect 29472 18426 29500 18838
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 29460 18420 29512 18426
rect 29460 18362 29512 18368
rect 29920 17604 29972 17610
rect 29920 17546 29972 17552
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29748 17202 29776 17478
rect 29736 17196 29788 17202
rect 29736 17138 29788 17144
rect 29748 16794 29776 17138
rect 29932 16998 29960 17546
rect 29920 16992 29972 16998
rect 29920 16934 29972 16940
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 29564 15434 29592 15982
rect 29748 15978 29776 16730
rect 29736 15972 29788 15978
rect 29736 15914 29788 15920
rect 29748 15706 29776 15914
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29000 15156 29052 15162
rect 29104 15150 29224 15178
rect 29000 15098 29052 15104
rect 29090 15056 29146 15065
rect 28920 15014 29040 15042
rect 29012 14958 29040 15014
rect 29090 14991 29146 15000
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 29012 14618 29040 14894
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 28816 14544 28868 14550
rect 28816 14486 28868 14492
rect 29104 14482 29132 14991
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 27896 14272 27948 14278
rect 27896 14214 27948 14220
rect 27908 14006 27936 14214
rect 29104 14074 29132 14418
rect 29196 14074 29224 15150
rect 29932 14618 29960 16934
rect 29920 14612 29972 14618
rect 29920 14554 29972 14560
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29184 14068 29236 14074
rect 29184 14010 29236 14016
rect 27896 14000 27948 14006
rect 27896 13942 27948 13948
rect 28540 14000 28592 14006
rect 28540 13942 28592 13948
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27908 13326 27936 13942
rect 28552 13705 28580 13942
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28538 13696 28594 13705
rect 28538 13631 28594 13640
rect 28644 13530 28672 13874
rect 29828 13728 29880 13734
rect 28998 13696 29054 13705
rect 28998 13631 29054 13640
rect 29748 13676 29828 13682
rect 29748 13670 29880 13676
rect 29748 13654 29868 13670
rect 29012 13530 29040 13631
rect 28632 13524 28684 13530
rect 28632 13466 28684 13472
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 27540 13110 27660 13138
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27540 12850 27568 13110
rect 27816 12986 27844 13262
rect 27804 12980 27856 12986
rect 27632 12940 27804 12968
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27528 12844 27580 12850
rect 27528 12786 27580 12792
rect 25320 12708 25372 12714
rect 25320 12650 25372 12656
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 24768 12232 24820 12238
rect 24688 12192 24768 12220
rect 24768 12174 24820 12180
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24596 11354 24624 11834
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24492 10532 24544 10538
rect 24492 10474 24544 10480
rect 24504 9382 24532 10474
rect 24582 9752 24638 9761
rect 24582 9687 24638 9696
rect 24596 9450 24624 9687
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24504 9110 24532 9318
rect 24596 9110 24624 9386
rect 24688 9178 24716 11494
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24780 10266 24808 11154
rect 25044 11008 25096 11014
rect 25044 10950 25096 10956
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25056 10470 25084 10950
rect 25424 10810 25452 10950
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 25884 10606 25912 12582
rect 26700 12232 26752 12238
rect 26700 12174 26752 12180
rect 26712 11694 26740 12174
rect 26988 12102 27016 12582
rect 27344 12368 27396 12374
rect 27344 12310 27396 12316
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26712 11218 26740 11630
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26700 11212 26752 11218
rect 26700 11154 26752 11160
rect 26896 11014 26924 11562
rect 26884 11008 26936 11014
rect 26884 10950 26936 10956
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 25056 10130 25084 10406
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 25884 9926 25912 10542
rect 26148 10532 26200 10538
rect 26148 10474 26200 10480
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25872 9920 25924 9926
rect 25872 9862 25924 9868
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24492 9104 24544 9110
rect 24492 9046 24544 9052
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24504 8634 24532 9046
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24400 8560 24452 8566
rect 24400 8502 24452 8508
rect 24596 8498 24624 9046
rect 25332 9042 25360 9862
rect 26160 9722 26188 10474
rect 26988 10266 27016 12038
rect 27356 10810 27384 12310
rect 27632 12306 27660 12940
rect 27804 12922 27856 12928
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27724 12442 27752 12786
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27632 11898 27660 12242
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27632 11801 27660 11834
rect 27618 11792 27674 11801
rect 27618 11727 27674 11736
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27436 11008 27488 11014
rect 27436 10950 27488 10956
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 27264 9761 27292 10406
rect 27356 10130 27384 10746
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27448 10062 27476 10950
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 27540 10282 27568 10474
rect 27632 10282 27660 11494
rect 27724 11286 27752 12378
rect 27908 12374 27936 13262
rect 28184 12986 28212 13330
rect 29748 13326 29776 13654
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29184 13320 29236 13326
rect 29184 13262 29236 13268
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 28172 12980 28224 12986
rect 28172 12922 28224 12928
rect 29196 12442 29224 13262
rect 29460 13184 29512 13190
rect 29460 13126 29512 13132
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 29184 12436 29236 12442
rect 29184 12378 29236 12384
rect 27896 12368 27948 12374
rect 27896 12310 27948 12316
rect 29276 11688 29328 11694
rect 29276 11630 29328 11636
rect 27712 11280 27764 11286
rect 27712 11222 27764 11228
rect 27724 10810 27752 11222
rect 29288 11150 29316 11630
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 29276 11144 29328 11150
rect 29276 11086 29328 11092
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 28736 10470 28764 11086
rect 29380 10674 29408 12922
rect 29472 12918 29500 13126
rect 29840 12986 29868 13330
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 29920 12980 29972 12986
rect 29920 12922 29972 12928
rect 29460 12912 29512 12918
rect 29460 12854 29512 12860
rect 29932 12782 29960 12922
rect 29920 12776 29972 12782
rect 29920 12718 29972 12724
rect 30024 12442 30052 13262
rect 29552 12436 29604 12442
rect 29552 12378 29604 12384
rect 30012 12436 30064 12442
rect 30012 12378 30064 12384
rect 29564 11898 29592 12378
rect 30010 12336 30066 12345
rect 30010 12271 30012 12280
rect 30064 12271 30066 12280
rect 30012 12242 30064 12248
rect 29552 11892 29604 11898
rect 29552 11834 29604 11840
rect 29564 11286 29592 11834
rect 30024 11558 30052 12242
rect 30012 11552 30064 11558
rect 30012 11494 30064 11500
rect 29552 11280 29604 11286
rect 29552 11222 29604 11228
rect 29564 10810 29592 11222
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 28724 10464 28776 10470
rect 28724 10406 28776 10412
rect 27540 10266 27660 10282
rect 27528 10260 27660 10266
rect 27580 10254 27660 10260
rect 27528 10202 27580 10208
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27250 9752 27306 9761
rect 26148 9716 26200 9722
rect 27448 9722 27476 9998
rect 27250 9687 27306 9696
rect 27436 9716 27488 9722
rect 26148 9658 26200 9664
rect 27436 9658 27488 9664
rect 27632 9654 27660 9998
rect 27620 9648 27672 9654
rect 27620 9590 27672 9596
rect 28264 9580 28316 9586
rect 28264 9522 28316 9528
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 26700 9444 26752 9450
rect 26700 9386 26752 9392
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 25332 8430 25360 8978
rect 26712 8634 26740 9386
rect 27344 9376 27396 9382
rect 27344 9318 27396 9324
rect 27436 9376 27488 9382
rect 27436 9318 27488 9324
rect 27160 9036 27212 9042
rect 27160 8978 27212 8984
rect 27172 8634 27200 8978
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 25332 7886 25360 8366
rect 26712 8022 26740 8570
rect 27356 8498 27384 9318
rect 27448 9178 27476 9318
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 26700 8016 26752 8022
rect 26700 7958 26752 7964
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26252 7546 26280 7822
rect 26712 7546 26740 7958
rect 27448 7750 27476 9114
rect 27632 8566 27660 9454
rect 28276 8974 28304 9522
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 28264 8968 28316 8974
rect 28316 8916 28396 8922
rect 28264 8910 28396 8916
rect 27712 8832 27764 8838
rect 27712 8774 27764 8780
rect 27620 8560 27672 8566
rect 27620 8502 27672 8508
rect 27724 8430 27752 8774
rect 28184 8634 28212 8910
rect 28276 8894 28396 8910
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27724 8090 27752 8366
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 27448 7342 27476 7686
rect 28184 7546 28212 8570
rect 28276 8498 28304 8774
rect 28368 8498 28396 8894
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28368 8090 28396 8434
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27252 7268 27304 7274
rect 27252 7210 27304 7216
rect 27264 6798 27292 7210
rect 27448 7002 27476 7278
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 28184 6934 28212 7482
rect 28172 6928 28224 6934
rect 28172 6870 28224 6876
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27264 6254 27292 6734
rect 27356 6458 27384 6802
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 27252 6248 27304 6254
rect 27252 6190 27304 6196
rect 28368 5710 28396 8026
rect 28736 7886 28764 10406
rect 28816 9036 28868 9042
rect 28816 8978 28868 8984
rect 29644 9036 29696 9042
rect 29644 8978 29696 8984
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 28736 7342 28764 7822
rect 28828 7410 28856 8978
rect 29000 8968 29052 8974
rect 28920 8916 29000 8922
rect 28920 8910 29052 8916
rect 28920 8894 29040 8910
rect 28816 7404 28868 7410
rect 28816 7346 28868 7352
rect 28724 7336 28776 7342
rect 28724 7278 28776 7284
rect 28828 6730 28856 7346
rect 28816 6724 28868 6730
rect 28816 6666 28868 6672
rect 28920 5914 28948 8894
rect 29656 8634 29684 8978
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29748 8634 29776 8910
rect 29932 8838 29960 8910
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29932 8401 29960 8774
rect 29918 8392 29974 8401
rect 29918 8327 29974 8336
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 29012 7546 29040 7890
rect 30208 7834 30236 33487
rect 33048 30592 33100 30598
rect 33048 30534 33100 30540
rect 33060 30258 33088 30534
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 32220 30048 32272 30054
rect 32220 29990 32272 29996
rect 32496 30048 32548 30054
rect 32496 29990 32548 29996
rect 32772 30048 32824 30054
rect 32772 29990 32824 29996
rect 31484 29096 31536 29102
rect 31484 29038 31536 29044
rect 31208 28960 31260 28966
rect 31208 28902 31260 28908
rect 31220 28762 31248 28902
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31220 28014 31248 28698
rect 31496 28422 31524 29038
rect 32232 28626 32260 29990
rect 32220 28620 32272 28626
rect 32220 28562 32272 28568
rect 31484 28416 31536 28422
rect 31484 28358 31536 28364
rect 31208 28008 31260 28014
rect 31208 27950 31260 27956
rect 31496 27946 31524 28358
rect 32232 28218 32260 28562
rect 32220 28212 32272 28218
rect 32220 28154 32272 28160
rect 31024 27940 31076 27946
rect 31024 27882 31076 27888
rect 31484 27940 31536 27946
rect 31484 27882 31536 27888
rect 31036 27674 31064 27882
rect 32312 27872 32364 27878
rect 32312 27814 32364 27820
rect 32324 27674 32352 27814
rect 31024 27668 31076 27674
rect 31024 27610 31076 27616
rect 32312 27668 32364 27674
rect 32312 27610 32364 27616
rect 30840 27532 30892 27538
rect 30840 27474 30892 27480
rect 30852 27130 30880 27474
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30852 26586 30880 26794
rect 31036 26586 31064 27610
rect 32128 27328 32180 27334
rect 31666 27296 31722 27305
rect 32128 27270 32180 27276
rect 31666 27231 31722 27240
rect 31680 27130 31708 27231
rect 31668 27124 31720 27130
rect 31668 27066 31720 27072
rect 32036 26784 32088 26790
rect 32036 26726 32088 26732
rect 32048 26586 32076 26726
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 31024 26580 31076 26586
rect 31024 26522 31076 26528
rect 32036 26580 32088 26586
rect 32036 26522 32088 26528
rect 31574 26480 31630 26489
rect 30288 26444 30340 26450
rect 31574 26415 31630 26424
rect 30288 26386 30340 26392
rect 30300 26058 30328 26386
rect 31300 26376 31352 26382
rect 31298 26344 31300 26353
rect 31352 26344 31354 26353
rect 31298 26279 31354 26288
rect 31208 26240 31260 26246
rect 31208 26182 31260 26188
rect 30300 26042 30420 26058
rect 31220 26042 31248 26182
rect 31588 26042 31616 26415
rect 31760 26240 31812 26246
rect 31760 26182 31812 26188
rect 30300 26036 30432 26042
rect 30300 26030 30380 26036
rect 30380 25978 30432 25984
rect 31208 26036 31260 26042
rect 31208 25978 31260 25984
rect 31576 26036 31628 26042
rect 31576 25978 31628 25984
rect 31588 25838 31616 25978
rect 31576 25832 31628 25838
rect 31576 25774 31628 25780
rect 30748 25764 30800 25770
rect 30748 25706 30800 25712
rect 30760 25498 30788 25706
rect 30748 25492 30800 25498
rect 30748 25434 30800 25440
rect 30564 24676 30616 24682
rect 30564 24618 30616 24624
rect 30576 24410 30604 24618
rect 30760 24410 30788 25434
rect 31772 24886 31800 26182
rect 32140 25362 32168 27270
rect 32324 27130 32352 27610
rect 32508 27606 32536 29990
rect 32784 29714 32812 29990
rect 32772 29708 32824 29714
rect 32772 29650 32824 29656
rect 32680 28960 32732 28966
rect 32680 28902 32732 28908
rect 32692 28626 32720 28902
rect 32680 28620 32732 28626
rect 32680 28562 32732 28568
rect 33060 28082 33088 30194
rect 34532 29866 34560 35566
rect 34808 34921 34836 37182
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35636 35834 35664 39335
rect 35806 36952 35862 36961
rect 35806 36887 35862 36896
rect 35624 35828 35676 35834
rect 35624 35770 35676 35776
rect 35622 35728 35678 35737
rect 35622 35663 35678 35672
rect 35530 35320 35586 35329
rect 35530 35255 35532 35264
rect 35584 35255 35586 35264
rect 35532 35226 35584 35232
rect 34794 34912 34850 34921
rect 34794 34847 34850 34856
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 35438 34640 35494 34649
rect 35438 34575 35494 34584
rect 35452 34202 35480 34575
rect 35532 34536 35584 34542
rect 35532 34478 35584 34484
rect 35440 34196 35492 34202
rect 35440 34138 35492 34144
rect 35256 34060 35308 34066
rect 35256 34002 35308 34008
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35268 33522 35296 34002
rect 35256 33516 35308 33522
rect 35256 33458 35308 33464
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34532 29838 34652 29866
rect 33600 29708 33652 29714
rect 33600 29650 33652 29656
rect 34520 29708 34572 29714
rect 34520 29650 34572 29656
rect 33508 29640 33560 29646
rect 33508 29582 33560 29588
rect 33520 29034 33548 29582
rect 33508 29028 33560 29034
rect 33508 28970 33560 28976
rect 33612 28966 33640 29650
rect 33600 28960 33652 28966
rect 33600 28902 33652 28908
rect 34244 28960 34296 28966
rect 34244 28902 34296 28908
rect 33612 28762 33640 28902
rect 33600 28756 33652 28762
rect 33600 28698 33652 28704
rect 34152 28688 34204 28694
rect 34152 28630 34204 28636
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 33048 28076 33100 28082
rect 33048 28018 33100 28024
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 32784 27606 32812 28018
rect 33796 27878 33824 28018
rect 33968 27940 34020 27946
rect 33968 27882 34020 27888
rect 33784 27872 33836 27878
rect 33782 27840 33784 27849
rect 33836 27840 33838 27849
rect 33782 27775 33838 27784
rect 32496 27600 32548 27606
rect 32496 27542 32548 27548
rect 32772 27600 32824 27606
rect 32772 27542 32824 27548
rect 32312 27124 32364 27130
rect 32312 27066 32364 27072
rect 32784 26994 32812 27542
rect 33508 27464 33560 27470
rect 33508 27406 33560 27412
rect 33232 27328 33284 27334
rect 33230 27296 33232 27305
rect 33284 27296 33286 27305
rect 33230 27231 33286 27240
rect 32772 26988 32824 26994
rect 32772 26930 32824 26936
rect 32680 26512 32732 26518
rect 32680 26454 32732 26460
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 32324 26042 32352 26318
rect 32692 26042 32720 26454
rect 32784 26382 32812 26930
rect 33244 26926 33272 27231
rect 33520 26994 33548 27406
rect 33508 26988 33560 26994
rect 33508 26930 33560 26936
rect 33232 26920 33284 26926
rect 33232 26862 33284 26868
rect 33048 26784 33100 26790
rect 33048 26726 33100 26732
rect 33232 26784 33284 26790
rect 33232 26726 33284 26732
rect 33060 26586 33088 26726
rect 33048 26580 33100 26586
rect 33048 26522 33100 26528
rect 33244 26489 33272 26726
rect 33230 26480 33286 26489
rect 33520 26450 33548 26930
rect 33784 26512 33836 26518
rect 33784 26454 33836 26460
rect 33230 26415 33286 26424
rect 33508 26444 33560 26450
rect 33508 26386 33560 26392
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 33140 26240 33192 26246
rect 33140 26182 33192 26188
rect 33692 26240 33744 26246
rect 33692 26182 33744 26188
rect 32312 26036 32364 26042
rect 32312 25978 32364 25984
rect 32680 26036 32732 26042
rect 32680 25978 32732 25984
rect 33152 25974 33180 26182
rect 33140 25968 33192 25974
rect 33140 25910 33192 25916
rect 33152 25838 33180 25910
rect 33140 25832 33192 25838
rect 33140 25774 33192 25780
rect 32772 25696 32824 25702
rect 32772 25638 32824 25644
rect 32864 25696 32916 25702
rect 32864 25638 32916 25644
rect 31944 25356 31996 25362
rect 31944 25298 31996 25304
rect 32128 25356 32180 25362
rect 32128 25298 32180 25304
rect 31300 24880 31352 24886
rect 31300 24822 31352 24828
rect 31760 24880 31812 24886
rect 31760 24822 31812 24828
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30748 24404 30800 24410
rect 30748 24346 30800 24352
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 30300 23322 30328 23666
rect 30576 23594 30604 24346
rect 31312 23866 31340 24822
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31864 24410 31892 24550
rect 31956 24410 31984 25298
rect 32034 24984 32090 24993
rect 32140 24954 32168 25298
rect 32784 25294 32812 25638
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32784 24954 32812 25230
rect 32876 25158 32904 25638
rect 33704 25362 33732 26182
rect 33796 25702 33824 26454
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 33888 25702 33916 26386
rect 33784 25696 33836 25702
rect 33784 25638 33836 25644
rect 33876 25696 33928 25702
rect 33876 25638 33928 25644
rect 33796 25498 33824 25638
rect 33784 25492 33836 25498
rect 33784 25434 33836 25440
rect 33692 25356 33744 25362
rect 33692 25298 33744 25304
rect 32864 25152 32916 25158
rect 32864 25094 32916 25100
rect 33416 25152 33468 25158
rect 33416 25094 33468 25100
rect 32034 24919 32090 24928
rect 32128 24948 32180 24954
rect 31852 24404 31904 24410
rect 31852 24346 31904 24352
rect 31944 24404 31996 24410
rect 31944 24346 31996 24352
rect 31956 24041 31984 24346
rect 32048 24274 32076 24919
rect 32128 24890 32180 24896
rect 32772 24948 32824 24954
rect 32772 24890 32824 24896
rect 32772 24812 32824 24818
rect 32772 24754 32824 24760
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 31942 24032 31998 24041
rect 31942 23967 31998 23976
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 30564 23588 30616 23594
rect 30564 23530 30616 23536
rect 30576 23322 30604 23530
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30564 23316 30616 23322
rect 30564 23258 30616 23264
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31220 22778 31248 23054
rect 31956 22778 31984 23967
rect 32048 23866 32076 24210
rect 32784 23866 32812 24754
rect 32876 24410 32904 25094
rect 33140 24948 33192 24954
rect 33140 24890 33192 24896
rect 32864 24404 32916 24410
rect 32864 24346 32916 24352
rect 33048 24404 33100 24410
rect 33048 24346 33100 24352
rect 32036 23860 32088 23866
rect 32036 23802 32088 23808
rect 32772 23860 32824 23866
rect 32772 23802 32824 23808
rect 33060 23186 33088 24346
rect 33152 23866 33180 24890
rect 33428 23866 33456 25094
rect 33704 24410 33732 25298
rect 33888 24954 33916 25638
rect 33876 24948 33928 24954
rect 33876 24890 33928 24896
rect 33876 24676 33928 24682
rect 33876 24618 33928 24624
rect 33692 24404 33744 24410
rect 33692 24346 33744 24352
rect 33888 23866 33916 24618
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 33416 23860 33468 23866
rect 33416 23802 33468 23808
rect 33876 23860 33928 23866
rect 33876 23802 33928 23808
rect 33152 23662 33180 23802
rect 33140 23656 33192 23662
rect 33140 23598 33192 23604
rect 33600 23248 33652 23254
rect 33600 23190 33652 23196
rect 33048 23180 33100 23186
rect 33048 23122 33100 23128
rect 33060 22778 33088 23122
rect 33232 22976 33284 22982
rect 33232 22918 33284 22924
rect 30748 22772 30800 22778
rect 30748 22714 30800 22720
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 31944 22772 31996 22778
rect 31944 22714 31996 22720
rect 33048 22772 33100 22778
rect 33048 22714 33100 22720
rect 30760 21418 30788 22714
rect 33140 22432 33192 22438
rect 33140 22374 33192 22380
rect 33152 22030 33180 22374
rect 32956 22024 33008 22030
rect 32956 21966 33008 21972
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 31208 21888 31260 21894
rect 31208 21830 31260 21836
rect 30748 21412 30800 21418
rect 30748 21354 30800 21360
rect 31220 21350 31248 21830
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31208 21344 31260 21350
rect 31208 21286 31260 21292
rect 31116 20256 31168 20262
rect 31022 20224 31078 20233
rect 31116 20198 31168 20204
rect 31022 20159 31078 20168
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30300 19174 30328 19314
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30484 18970 30512 19314
rect 30748 19304 30800 19310
rect 30748 19246 30800 19252
rect 30760 19174 30788 19246
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30932 19168 30984 19174
rect 30932 19110 30984 19116
rect 30944 18970 30972 19110
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 30484 18290 30512 18906
rect 30944 18426 30972 18906
rect 31036 18766 31064 20159
rect 31128 19378 31156 20198
rect 31116 19372 31168 19378
rect 31116 19314 31168 19320
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 31036 18426 31064 18702
rect 31220 18698 31248 21286
rect 31588 21146 31616 21490
rect 31852 21480 31904 21486
rect 31852 21422 31904 21428
rect 31668 21412 31720 21418
rect 31668 21354 31720 21360
rect 31576 21140 31628 21146
rect 31576 21082 31628 21088
rect 31588 20058 31616 21082
rect 31680 20466 31708 21354
rect 31864 21146 31892 21422
rect 32968 21146 32996 21966
rect 33140 21888 33192 21894
rect 33140 21830 33192 21836
rect 33152 21554 33180 21830
rect 33244 21690 33272 22918
rect 33612 22506 33640 23190
rect 33600 22500 33652 22506
rect 33600 22442 33652 22448
rect 33980 22234 34008 27882
rect 34058 25392 34114 25401
rect 34058 25327 34114 25336
rect 34072 25294 34100 25327
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 34072 24410 34100 25230
rect 34060 24404 34112 24410
rect 34060 24346 34112 24352
rect 34060 23112 34112 23118
rect 34060 23054 34112 23060
rect 34072 22234 34100 23054
rect 34164 22658 34192 28630
rect 34256 28422 34284 28902
rect 34244 28416 34296 28422
rect 34244 28358 34296 28364
rect 34256 27878 34284 28358
rect 34532 28234 34560 29650
rect 34348 28206 34560 28234
rect 34244 27872 34296 27878
rect 34244 27814 34296 27820
rect 34244 27328 34296 27334
rect 34244 27270 34296 27276
rect 34256 26382 34284 27270
rect 34348 27010 34376 28206
rect 34518 28112 34574 28121
rect 34518 28047 34574 28056
rect 34532 27554 34560 28047
rect 34624 27946 34652 29838
rect 34704 29504 34756 29510
rect 34704 29446 34756 29452
rect 34716 28966 34744 29446
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34980 29232 35032 29238
rect 34980 29174 35032 29180
rect 34704 28960 34756 28966
rect 34704 28902 34756 28908
rect 34716 28626 34744 28902
rect 34704 28620 34756 28626
rect 34704 28562 34756 28568
rect 34716 28218 34744 28562
rect 34704 28212 34756 28218
rect 34704 28154 34756 28160
rect 34612 27940 34664 27946
rect 34612 27882 34664 27888
rect 34704 27872 34756 27878
rect 34704 27814 34756 27820
rect 34440 27538 34560 27554
rect 34612 27600 34664 27606
rect 34612 27542 34664 27548
rect 34428 27532 34560 27538
rect 34480 27526 34560 27532
rect 34428 27474 34480 27480
rect 34440 27130 34468 27474
rect 34428 27124 34480 27130
rect 34428 27066 34480 27072
rect 34348 26982 34560 27010
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34244 26376 34296 26382
rect 34244 26318 34296 26324
rect 34256 25906 34284 26318
rect 34244 25900 34296 25906
rect 34244 25842 34296 25848
rect 34256 25498 34284 25842
rect 34244 25492 34296 25498
rect 34244 25434 34296 25440
rect 34440 24750 34468 26726
rect 34428 24744 34480 24750
rect 34428 24686 34480 24692
rect 34532 23769 34560 26982
rect 34518 23760 34574 23769
rect 34428 23724 34480 23730
rect 34518 23695 34574 23704
rect 34428 23666 34480 23672
rect 34244 23520 34296 23526
rect 34244 23462 34296 23468
rect 34256 23254 34284 23462
rect 34440 23254 34468 23666
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 34532 23322 34560 23598
rect 34520 23316 34572 23322
rect 34520 23258 34572 23264
rect 34244 23248 34296 23254
rect 34244 23190 34296 23196
rect 34428 23248 34480 23254
rect 34428 23190 34480 23196
rect 34440 22778 34468 23190
rect 34428 22772 34480 22778
rect 34428 22714 34480 22720
rect 34164 22630 34468 22658
rect 34244 22568 34296 22574
rect 34244 22510 34296 22516
rect 34152 22500 34204 22506
rect 34152 22442 34204 22448
rect 33968 22228 34020 22234
rect 33968 22170 34020 22176
rect 34060 22228 34112 22234
rect 34060 22170 34112 22176
rect 33600 22092 33652 22098
rect 33600 22034 33652 22040
rect 33232 21684 33284 21690
rect 33232 21626 33284 21632
rect 33140 21548 33192 21554
rect 33140 21490 33192 21496
rect 33244 21486 33272 21626
rect 33232 21480 33284 21486
rect 33232 21422 33284 21428
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 31852 21140 31904 21146
rect 31852 21082 31904 21088
rect 32956 21140 33008 21146
rect 32956 21082 33008 21088
rect 33140 20936 33192 20942
rect 33244 20913 33272 21286
rect 33612 21146 33640 22034
rect 33980 21570 34008 22170
rect 33980 21542 34100 21570
rect 34072 21486 34100 21542
rect 33968 21480 34020 21486
rect 33968 21422 34020 21428
rect 34060 21480 34112 21486
rect 34060 21422 34112 21428
rect 33876 21344 33928 21350
rect 33876 21286 33928 21292
rect 33600 21140 33652 21146
rect 33600 21082 33652 21088
rect 33692 20936 33744 20942
rect 33140 20878 33192 20884
rect 33230 20904 33286 20913
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31852 20460 31904 20466
rect 31852 20402 31904 20408
rect 31576 20052 31628 20058
rect 31576 19994 31628 20000
rect 31680 18970 31708 20402
rect 31760 20324 31812 20330
rect 31760 20266 31812 20272
rect 31772 20097 31800 20266
rect 31758 20088 31814 20097
rect 31864 20058 31892 20402
rect 32956 20256 33008 20262
rect 33152 20244 33180 20878
rect 33692 20878 33744 20884
rect 33230 20839 33286 20848
rect 33704 20602 33732 20878
rect 33692 20596 33744 20602
rect 33692 20538 33744 20544
rect 33008 20216 33180 20244
rect 33324 20256 33376 20262
rect 33322 20224 33324 20233
rect 33376 20224 33378 20233
rect 32956 20198 33008 20204
rect 31758 20023 31814 20032
rect 31852 20052 31904 20058
rect 31852 19994 31904 20000
rect 32968 19718 32996 20198
rect 33322 20159 33378 20168
rect 33704 20058 33732 20538
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 33692 20052 33744 20058
rect 33692 19994 33744 20000
rect 32956 19712 33008 19718
rect 33008 19660 33180 19666
rect 32956 19654 33180 19660
rect 32968 19638 33180 19654
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 31668 18964 31720 18970
rect 31668 18906 31720 18912
rect 31208 18692 31260 18698
rect 31208 18634 31260 18640
rect 32772 18624 32824 18630
rect 32772 18566 32824 18572
rect 30932 18420 30984 18426
rect 30932 18362 30984 18368
rect 31024 18420 31076 18426
rect 31024 18362 31076 18368
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30392 15706 30420 17614
rect 31668 17536 31720 17542
rect 31668 17478 31720 17484
rect 32128 17536 32180 17542
rect 32128 17478 32180 17484
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 30380 15700 30432 15706
rect 30380 15642 30432 15648
rect 30288 15360 30340 15366
rect 30286 15328 30288 15337
rect 30340 15328 30342 15337
rect 30286 15263 30342 15272
rect 30392 15162 30420 15642
rect 30484 15638 30512 17206
rect 31390 17096 31446 17105
rect 31680 17066 31708 17478
rect 31390 17031 31392 17040
rect 31444 17031 31446 17040
rect 31668 17060 31720 17066
rect 31392 17002 31444 17008
rect 31668 17002 31720 17008
rect 31852 17060 31904 17066
rect 31852 17002 31904 17008
rect 31116 16992 31168 16998
rect 31116 16934 31168 16940
rect 30564 16652 30616 16658
rect 30564 16594 30616 16600
rect 30576 15745 30604 16594
rect 30932 15904 30984 15910
rect 30932 15846 30984 15852
rect 30562 15736 30618 15745
rect 30562 15671 30618 15680
rect 30472 15632 30524 15638
rect 30472 15574 30524 15580
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30484 14618 30512 15574
rect 30944 15502 30972 15846
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 30932 15496 30984 15502
rect 30932 15438 30984 15444
rect 30944 15162 30972 15438
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 30472 14612 30524 14618
rect 30472 14554 30524 14560
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30392 13938 30420 14214
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 30300 13530 30328 13806
rect 31036 13530 31064 15642
rect 31128 15434 31156 16934
rect 31208 15904 31260 15910
rect 31208 15846 31260 15852
rect 31116 15428 31168 15434
rect 31116 15370 31168 15376
rect 31128 14958 31156 15370
rect 31116 14952 31168 14958
rect 31116 14894 31168 14900
rect 31116 13864 31168 13870
rect 31116 13806 31168 13812
rect 30288 13524 30340 13530
rect 30288 13466 30340 13472
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 30300 12782 30328 13466
rect 30656 13252 30708 13258
rect 30656 13194 30708 13200
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30378 11792 30434 11801
rect 30378 11727 30434 11736
rect 30392 11354 30420 11727
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30668 10606 30696 13194
rect 31036 12986 31064 13466
rect 31024 12980 31076 12986
rect 31024 12922 31076 12928
rect 31036 12238 31064 12922
rect 31128 12442 31156 13806
rect 31220 12594 31248 15846
rect 31864 15473 31892 17002
rect 32140 16794 32168 17478
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 32036 16652 32088 16658
rect 32036 16594 32088 16600
rect 32048 16114 32076 16594
rect 32140 16130 32168 16730
rect 32140 16114 32260 16130
rect 32036 16108 32088 16114
rect 32140 16108 32272 16114
rect 32140 16102 32220 16108
rect 32036 16050 32088 16056
rect 32220 16050 32272 16056
rect 32048 15706 32076 16050
rect 32036 15700 32088 15706
rect 32036 15642 32088 15648
rect 32416 15638 32444 18226
rect 32784 18222 32812 18566
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32680 18080 32732 18086
rect 32678 18048 32680 18057
rect 32732 18048 32734 18057
rect 32678 17983 32734 17992
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32508 16794 32536 17682
rect 32680 17672 32732 17678
rect 32680 17614 32732 17620
rect 32692 16998 32720 17614
rect 32680 16992 32732 16998
rect 32680 16934 32732 16940
rect 32496 16788 32548 16794
rect 32496 16730 32548 16736
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32508 15910 32536 16186
rect 32588 16040 32640 16046
rect 32588 15982 32640 15988
rect 32496 15904 32548 15910
rect 32496 15846 32548 15852
rect 32404 15632 32456 15638
rect 32404 15574 32456 15580
rect 31850 15464 31906 15473
rect 31850 15399 31906 15408
rect 32416 15162 32444 15574
rect 32600 15366 32628 15982
rect 32588 15360 32640 15366
rect 32784 15337 32812 18158
rect 32864 17740 32916 17746
rect 32864 17682 32916 17688
rect 32876 17066 32904 17682
rect 32864 17060 32916 17066
rect 32864 17002 32916 17008
rect 32588 15302 32640 15308
rect 32770 15328 32826 15337
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31300 14476 31352 14482
rect 31300 14418 31352 14424
rect 31312 14074 31340 14418
rect 31496 14278 31524 14758
rect 32600 14482 32628 15302
rect 32770 15263 32826 15272
rect 32784 14550 32812 15263
rect 32876 14618 32904 17002
rect 33060 16980 33088 19450
rect 33152 19394 33180 19638
rect 33244 19514 33272 19994
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33232 19508 33284 19514
rect 33232 19450 33284 19456
rect 33152 19366 33272 19394
rect 33428 19378 33456 19790
rect 33244 18970 33272 19366
rect 33416 19372 33468 19378
rect 33416 19314 33468 19320
rect 33704 19174 33732 19790
rect 33888 19360 33916 21286
rect 33980 20942 34008 21422
rect 33968 20936 34020 20942
rect 33968 20878 34020 20884
rect 33980 20602 34008 20878
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 33888 19332 34008 19360
rect 33782 19272 33838 19281
rect 33782 19207 33784 19216
rect 33836 19207 33838 19216
rect 33784 19178 33836 19184
rect 33692 19168 33744 19174
rect 33692 19110 33744 19116
rect 33232 18964 33284 18970
rect 33232 18906 33284 18912
rect 32968 16952 33180 16980
rect 32968 16250 32996 16952
rect 33152 16794 33180 16952
rect 33048 16788 33100 16794
rect 33048 16730 33100 16736
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 32954 15464 33010 15473
rect 32954 15399 33010 15408
rect 32864 14612 32916 14618
rect 32864 14554 32916 14560
rect 32772 14544 32824 14550
rect 32772 14486 32824 14492
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 31484 14272 31536 14278
rect 31484 14214 31536 14220
rect 31496 14074 31524 14214
rect 31300 14068 31352 14074
rect 31300 14010 31352 14016
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31760 14000 31812 14006
rect 31760 13942 31812 13948
rect 31668 13864 31720 13870
rect 31668 13806 31720 13812
rect 31680 13258 31708 13806
rect 31772 13530 31800 13942
rect 32600 13734 32628 14418
rect 32784 14074 32812 14486
rect 32968 14414 32996 15399
rect 33060 15026 33088 16730
rect 33244 16674 33272 18906
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 33796 18426 33824 18702
rect 33784 18420 33836 18426
rect 33784 18362 33836 18368
rect 33416 18148 33468 18154
rect 33416 18090 33468 18096
rect 33324 17740 33376 17746
rect 33324 17682 33376 17688
rect 33336 16998 33364 17682
rect 33324 16992 33376 16998
rect 33324 16934 33376 16940
rect 33152 16658 33272 16674
rect 33140 16652 33272 16658
rect 33192 16646 33272 16652
rect 33140 16594 33192 16600
rect 33152 15162 33180 16594
rect 33232 16584 33284 16590
rect 33336 16572 33364 16934
rect 33428 16658 33456 18090
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33284 16544 33364 16572
rect 33232 16526 33284 16532
rect 33244 16454 33272 16526
rect 33232 16448 33284 16454
rect 33232 16390 33284 16396
rect 33244 16114 33272 16390
rect 33428 16250 33456 16594
rect 33416 16244 33468 16250
rect 33416 16186 33468 16192
rect 33232 16108 33284 16114
rect 33232 16050 33284 16056
rect 33876 15496 33928 15502
rect 33876 15438 33928 15444
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 33888 14822 33916 15438
rect 33876 14816 33928 14822
rect 33876 14758 33928 14764
rect 32956 14408 33008 14414
rect 32956 14350 33008 14356
rect 32968 14074 32996 14350
rect 33888 14278 33916 14758
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33876 14272 33928 14278
rect 33876 14214 33928 14220
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32956 14068 33008 14074
rect 32956 14010 33008 14016
rect 32588 13728 32640 13734
rect 32588 13670 32640 13676
rect 31760 13524 31812 13530
rect 31760 13466 31812 13472
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 31300 12640 31352 12646
rect 31220 12588 31300 12594
rect 31220 12582 31352 12588
rect 31220 12566 31340 12582
rect 31116 12436 31168 12442
rect 31116 12378 31168 12384
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 31128 11694 31156 12378
rect 31116 11688 31168 11694
rect 31220 11665 31248 12566
rect 32404 12300 32456 12306
rect 32404 12242 32456 12248
rect 31944 12232 31996 12238
rect 31944 12174 31996 12180
rect 31116 11630 31168 11636
rect 31206 11656 31262 11665
rect 31206 11591 31262 11600
rect 31666 11656 31722 11665
rect 31666 11591 31668 11600
rect 31220 10690 31248 11591
rect 31720 11591 31722 11600
rect 31668 11562 31720 11568
rect 31760 11552 31812 11558
rect 31760 11494 31812 11500
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31220 10662 31340 10690
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 31208 10600 31260 10606
rect 31208 10542 31260 10548
rect 30668 10266 30696 10542
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 30852 10266 30880 10406
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30840 10260 30892 10266
rect 30840 10202 30892 10208
rect 31036 10198 31064 10406
rect 31024 10192 31076 10198
rect 31024 10134 31076 10140
rect 31116 9920 31168 9926
rect 31116 9862 31168 9868
rect 31128 9518 31156 9862
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 31128 9178 31156 9454
rect 31220 9382 31248 10542
rect 31208 9376 31260 9382
rect 31208 9318 31260 9324
rect 31220 9178 31248 9318
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 31208 9172 31260 9178
rect 31208 9114 31260 9120
rect 30840 8900 30892 8906
rect 30840 8842 30892 8848
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30300 8498 30328 8774
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 30024 7806 30236 7834
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 29012 5846 29040 7482
rect 29276 7336 29328 7342
rect 29276 7278 29328 7284
rect 29092 6928 29144 6934
rect 29092 6870 29144 6876
rect 29104 6458 29132 6870
rect 29288 6866 29316 7278
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29092 6452 29144 6458
rect 29092 6394 29144 6400
rect 29104 5914 29132 6394
rect 29564 6254 29592 6802
rect 29552 6248 29604 6254
rect 29552 6190 29604 6196
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29092 5908 29144 5914
rect 29092 5850 29144 5856
rect 29000 5840 29052 5846
rect 28920 5788 29000 5794
rect 28920 5782 29052 5788
rect 28920 5766 29040 5782
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 28368 5370 28396 5646
rect 28920 5370 28948 5766
rect 29104 5370 29132 5850
rect 29564 5846 29592 6190
rect 29840 5914 29868 6190
rect 29828 5908 29880 5914
rect 29828 5850 29880 5856
rect 29552 5840 29604 5846
rect 29552 5782 29604 5788
rect 28356 5364 28408 5370
rect 28356 5306 28408 5312
rect 28908 5364 28960 5370
rect 28908 5306 28960 5312
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 23294 4040 23350 4049
rect 23294 3975 23350 3984
rect 23938 4040 23994 4049
rect 23938 3975 23994 3984
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 16670 3360 16726 3369
rect 4220 3292 4516 3312
rect 16670 3295 16726 3304
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 3330 2408 3386 2417
rect 3330 2343 3386 2352
rect 3344 480 3372 2343
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 9968 480 9996 2246
rect 16684 480 16712 3295
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 23308 480 23336 3975
rect 30024 480 30052 7806
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 6934 30144 7686
rect 30104 6928 30156 6934
rect 30104 6870 30156 6876
rect 30300 6746 30328 8298
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 30392 7478 30420 8230
rect 30852 8090 30880 8842
rect 30840 8084 30892 8090
rect 30840 8026 30892 8032
rect 30380 7472 30432 7478
rect 30380 7414 30432 7420
rect 30932 7472 30984 7478
rect 30932 7414 30984 7420
rect 30300 6718 30420 6746
rect 30392 6662 30420 6718
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30392 6254 30420 6598
rect 30944 6458 30972 7414
rect 30932 6452 30984 6458
rect 30932 6394 30984 6400
rect 30380 6248 30432 6254
rect 30380 6190 30432 6196
rect 31312 3369 31340 10662
rect 31496 10266 31524 11086
rect 31772 10810 31800 11494
rect 31956 11354 31984 12174
rect 32036 12096 32088 12102
rect 32036 12038 32088 12044
rect 32048 11830 32076 12038
rect 32416 11898 32444 12242
rect 32600 12102 32628 13670
rect 32956 13524 33008 13530
rect 32956 13466 33008 13472
rect 32968 12714 32996 13466
rect 33520 13326 33548 14214
rect 33692 13388 33744 13394
rect 33692 13330 33744 13336
rect 33508 13320 33560 13326
rect 33508 13262 33560 13268
rect 33048 12912 33100 12918
rect 33048 12854 33100 12860
rect 32956 12708 33008 12714
rect 32956 12650 33008 12656
rect 32496 12096 32548 12102
rect 32496 12038 32548 12044
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32404 11892 32456 11898
rect 32404 11834 32456 11840
rect 32036 11824 32088 11830
rect 32036 11766 32088 11772
rect 32416 11626 32444 11834
rect 32508 11626 32536 12038
rect 32404 11620 32456 11626
rect 32404 11562 32456 11568
rect 32496 11620 32548 11626
rect 32496 11562 32548 11568
rect 32508 11354 32536 11562
rect 31944 11348 31996 11354
rect 31944 11290 31996 11296
rect 32496 11348 32548 11354
rect 32496 11290 32548 11296
rect 31760 10804 31812 10810
rect 31760 10746 31812 10752
rect 31772 10606 31800 10746
rect 32508 10674 32536 11290
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 31760 10600 31812 10606
rect 31760 10542 31812 10548
rect 32692 10538 32720 11154
rect 32968 10810 32996 12650
rect 33060 11370 33088 12854
rect 33520 12782 33548 13262
rect 33704 12850 33732 13330
rect 33692 12844 33744 12850
rect 33692 12786 33744 12792
rect 33416 12776 33468 12782
rect 33416 12718 33468 12724
rect 33508 12776 33560 12782
rect 33508 12718 33560 12724
rect 33428 12238 33456 12718
rect 33232 12232 33284 12238
rect 33232 12174 33284 12180
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33244 11694 33272 12174
rect 33520 11898 33548 12718
rect 33704 11898 33732 12786
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 33980 11762 34008 19332
rect 34060 19168 34112 19174
rect 34060 19110 34112 19116
rect 34072 18834 34100 19110
rect 34164 18970 34192 22442
rect 34256 21010 34284 22510
rect 34440 21332 34468 22630
rect 34624 21978 34652 27542
rect 34716 27470 34744 27814
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34716 27010 34744 27406
rect 34808 27130 34836 29174
rect 34992 28694 35020 29174
rect 34980 28688 35032 28694
rect 34980 28630 35032 28636
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35072 28008 35124 28014
rect 35072 27950 35124 27956
rect 35084 27674 35112 27950
rect 35072 27668 35124 27674
rect 35072 27610 35124 27616
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34796 27124 34848 27130
rect 34796 27066 34848 27072
rect 34716 26982 34836 27010
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 34716 26042 34744 26386
rect 34808 26382 34836 26982
rect 34980 26852 35032 26858
rect 34980 26794 35032 26800
rect 34992 26586 35020 26794
rect 34980 26580 35032 26586
rect 34980 26522 35032 26528
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 34808 25702 34836 26318
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34704 25424 34756 25430
rect 34704 25366 34756 25372
rect 34716 24954 34744 25366
rect 34808 25158 34836 25638
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34704 24948 34756 24954
rect 34808 24936 34836 25094
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34808 24908 34928 24936
rect 34704 24890 34756 24896
rect 34796 24608 34848 24614
rect 34796 24550 34848 24556
rect 34808 23662 34836 24550
rect 34900 24274 34928 24908
rect 34888 24268 34940 24274
rect 34888 24210 34940 24216
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 35268 23712 35296 33458
rect 35348 33312 35400 33318
rect 35348 33254 35400 33260
rect 35360 27606 35388 33254
rect 35440 31884 35492 31890
rect 35440 31826 35492 31832
rect 35452 31142 35480 31826
rect 35440 31136 35492 31142
rect 35440 31078 35492 31084
rect 35348 27600 35400 27606
rect 35348 27542 35400 27548
rect 35268 23684 35388 23712
rect 34796 23656 34848 23662
rect 34796 23598 34848 23604
rect 35254 23624 35310 23633
rect 35254 23559 35310 23568
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 34888 22568 34940 22574
rect 34888 22510 34940 22516
rect 34900 22234 34928 22510
rect 34888 22228 34940 22234
rect 34888 22170 34940 22176
rect 34704 22092 34756 22098
rect 34704 22034 34756 22040
rect 34532 21950 34652 21978
rect 34532 21622 34560 21950
rect 34716 21690 34744 22034
rect 34796 22024 34848 22030
rect 35268 22001 35296 23559
rect 34796 21966 34848 21972
rect 35254 21992 35310 22001
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 34520 21616 34572 21622
rect 34520 21558 34572 21564
rect 34532 21486 34560 21558
rect 34808 21486 34836 21966
rect 35254 21927 35310 21936
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35360 21672 35388 23684
rect 35176 21644 35388 21672
rect 34520 21480 34572 21486
rect 34520 21422 34572 21428
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 34796 21480 34848 21486
rect 34796 21422 34848 21428
rect 34612 21412 34664 21418
rect 34612 21354 34664 21360
rect 34440 21304 34560 21332
rect 34244 21004 34296 21010
rect 34244 20946 34296 20952
rect 34256 20602 34284 20946
rect 34244 20596 34296 20602
rect 34244 20538 34296 20544
rect 34256 20040 34284 20538
rect 34336 20052 34388 20058
rect 34256 20012 34336 20040
rect 34336 19994 34388 20000
rect 34428 19780 34480 19786
rect 34428 19722 34480 19728
rect 34242 19544 34298 19553
rect 34242 19479 34298 19488
rect 34152 18964 34204 18970
rect 34152 18906 34204 18912
rect 34060 18828 34112 18834
rect 34060 18770 34112 18776
rect 34072 18426 34100 18770
rect 34164 18426 34192 18906
rect 34060 18420 34112 18426
rect 34060 18362 34112 18368
rect 34152 18420 34204 18426
rect 34152 18362 34204 18368
rect 34152 18148 34204 18154
rect 34152 18090 34204 18096
rect 34164 12594 34192 18090
rect 34256 17882 34284 19479
rect 34440 18698 34468 19722
rect 34428 18692 34480 18698
rect 34428 18634 34480 18640
rect 34244 17876 34296 17882
rect 34244 17818 34296 17824
rect 34256 17338 34284 17818
rect 34336 17536 34388 17542
rect 34336 17478 34388 17484
rect 34244 17332 34296 17338
rect 34244 17274 34296 17280
rect 34256 16794 34284 17274
rect 34348 17202 34376 17478
rect 34336 17196 34388 17202
rect 34336 17138 34388 17144
rect 34428 17060 34480 17066
rect 34428 17002 34480 17008
rect 34244 16788 34296 16794
rect 34244 16730 34296 16736
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 34244 15564 34296 15570
rect 34244 15506 34296 15512
rect 34256 15366 34284 15506
rect 34348 15502 34376 15982
rect 34336 15496 34388 15502
rect 34336 15438 34388 15444
rect 34244 15360 34296 15366
rect 34244 15302 34296 15308
rect 34256 15162 34284 15302
rect 34440 15162 34468 17002
rect 34244 15156 34296 15162
rect 34244 15098 34296 15104
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34256 15026 34284 15098
rect 34244 15020 34296 15026
rect 34244 14962 34296 14968
rect 34256 14618 34284 14962
rect 34244 14612 34296 14618
rect 34244 14554 34296 14560
rect 34428 13728 34480 13734
rect 34428 13670 34480 13676
rect 34164 12566 34284 12594
rect 34256 12442 34284 12566
rect 34244 12436 34296 12442
rect 34244 12378 34296 12384
rect 34244 12300 34296 12306
rect 34244 12242 34296 12248
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 34164 11898 34192 12174
rect 34152 11892 34204 11898
rect 34152 11834 34204 11840
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 34152 11756 34204 11762
rect 34152 11698 34204 11704
rect 33232 11688 33284 11694
rect 33232 11630 33284 11636
rect 33060 11342 33180 11370
rect 33152 11286 33180 11342
rect 33140 11280 33192 11286
rect 33140 11222 33192 11228
rect 32956 10804 33008 10810
rect 32956 10746 33008 10752
rect 33046 10704 33102 10713
rect 32968 10662 33046 10690
rect 32680 10532 32732 10538
rect 32680 10474 32732 10480
rect 32404 10464 32456 10470
rect 32404 10406 32456 10412
rect 32416 10266 32444 10406
rect 31484 10260 31536 10266
rect 31484 10202 31536 10208
rect 32404 10260 32456 10266
rect 32404 10202 32456 10208
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 32496 10192 32548 10198
rect 32496 10134 32548 10140
rect 32508 9722 32536 10134
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32600 9654 32628 10202
rect 32588 9648 32640 9654
rect 32588 9590 32640 9596
rect 31576 9444 31628 9450
rect 31576 9386 31628 9392
rect 31588 9217 31616 9386
rect 31574 9208 31630 9217
rect 31574 9143 31630 9152
rect 32692 9110 32720 10474
rect 32968 9586 32996 10662
rect 33046 10639 33048 10648
rect 33100 10639 33102 10648
rect 33048 10610 33100 10616
rect 33140 10600 33192 10606
rect 33060 10548 33140 10554
rect 33060 10542 33192 10548
rect 33060 10526 33180 10542
rect 33416 10532 33468 10538
rect 33060 9654 33088 10526
rect 33416 10474 33468 10480
rect 33428 10062 33456 10474
rect 33692 10464 33744 10470
rect 33692 10406 33744 10412
rect 33704 10266 33732 10406
rect 33692 10260 33744 10266
rect 33692 10202 33744 10208
rect 33968 10124 34020 10130
rect 33968 10066 34020 10072
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33980 9722 34008 10066
rect 34164 9722 34192 11698
rect 34256 10266 34284 12242
rect 34440 11354 34468 13670
rect 34428 11348 34480 11354
rect 34428 11290 34480 11296
rect 34440 10810 34468 11290
rect 34532 11082 34560 21304
rect 34624 17338 34652 21354
rect 34716 18154 34744 21422
rect 35176 21350 35204 21644
rect 35452 21593 35480 31078
rect 35544 29714 35572 34478
rect 35636 33658 35664 35663
rect 35716 35148 35768 35154
rect 35716 35090 35768 35096
rect 35728 34542 35756 35090
rect 35820 34746 35848 36887
rect 36096 35601 36124 39520
rect 36726 38176 36782 38185
rect 36726 38111 36782 38120
rect 36082 35592 36138 35601
rect 36082 35527 36138 35536
rect 36740 34746 36768 38111
rect 37200 35193 37228 39520
rect 38304 35329 38332 39520
rect 38290 35320 38346 35329
rect 38290 35255 38346 35264
rect 37186 35184 37242 35193
rect 37186 35119 37242 35128
rect 35808 34740 35860 34746
rect 35808 34682 35860 34688
rect 36728 34740 36780 34746
rect 36728 34682 36780 34688
rect 39408 34649 39436 39520
rect 39394 34640 39450 34649
rect 39394 34575 39450 34584
rect 35716 34536 35768 34542
rect 37096 34536 37148 34542
rect 35716 34478 35768 34484
rect 35806 34504 35862 34513
rect 35624 33652 35676 33658
rect 35624 33594 35676 33600
rect 35728 33561 35756 34478
rect 37096 34478 37148 34484
rect 35806 34439 35862 34448
rect 35714 33552 35770 33561
rect 35714 33487 35770 33496
rect 35622 33280 35678 33289
rect 35622 33215 35678 33224
rect 35636 30938 35664 33215
rect 35714 32056 35770 32065
rect 35820 32026 35848 34439
rect 35714 31991 35770 32000
rect 35808 32020 35860 32026
rect 35624 30932 35676 30938
rect 35624 30874 35676 30880
rect 35624 30796 35676 30802
rect 35624 30738 35676 30744
rect 35636 30054 35664 30738
rect 35728 30326 35756 31991
rect 35808 31962 35860 31968
rect 35898 30832 35954 30841
rect 35898 30767 35954 30776
rect 35716 30320 35768 30326
rect 35716 30262 35768 30268
rect 35716 30184 35768 30190
rect 35716 30126 35768 30132
rect 35624 30048 35676 30054
rect 35624 29990 35676 29996
rect 35532 29708 35584 29714
rect 35532 29650 35584 29656
rect 35530 29608 35586 29617
rect 35530 29543 35586 29552
rect 35544 26042 35572 29543
rect 35636 27826 35664 29990
rect 35728 29238 35756 30126
rect 35912 29850 35940 30767
rect 35900 29844 35952 29850
rect 35900 29786 35952 29792
rect 35808 29708 35860 29714
rect 35808 29650 35860 29656
rect 35716 29232 35768 29238
rect 35716 29174 35768 29180
rect 35716 29096 35768 29102
rect 35716 29038 35768 29044
rect 35728 28762 35756 29038
rect 35820 29034 35848 29650
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 35912 29170 35940 29446
rect 35900 29164 35952 29170
rect 35900 29106 35952 29112
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35716 28756 35768 28762
rect 35716 28698 35768 28704
rect 35728 28014 35756 28698
rect 35716 28008 35768 28014
rect 35716 27950 35768 27956
rect 35636 27798 35756 27826
rect 35624 26240 35676 26246
rect 35624 26182 35676 26188
rect 35532 26036 35584 26042
rect 35532 25978 35584 25984
rect 35544 25770 35572 25978
rect 35636 25838 35664 26182
rect 35624 25832 35676 25838
rect 35624 25774 35676 25780
rect 35532 25764 35584 25770
rect 35532 25706 35584 25712
rect 35636 25430 35664 25774
rect 35624 25424 35676 25430
rect 35624 25366 35676 25372
rect 35532 24268 35584 24274
rect 35532 24210 35584 24216
rect 35544 23322 35572 24210
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35636 23730 35664 24006
rect 35624 23724 35676 23730
rect 35624 23666 35676 23672
rect 35532 23316 35584 23322
rect 35532 23258 35584 23264
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35544 22574 35572 22918
rect 35532 22568 35584 22574
rect 35532 22510 35584 22516
rect 35728 21978 35756 27798
rect 35544 21950 35756 21978
rect 35254 21584 35310 21593
rect 35254 21519 35310 21528
rect 35438 21584 35494 21593
rect 35438 21519 35494 21528
rect 35164 21344 35216 21350
rect 35164 21286 35216 21292
rect 35176 21146 35204 21286
rect 35164 21140 35216 21146
rect 35164 21082 35216 21088
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34796 20596 34848 20602
rect 34796 20538 34848 20544
rect 34808 19145 34836 20538
rect 35164 20392 35216 20398
rect 35164 20334 35216 20340
rect 35176 20058 35204 20334
rect 35164 20052 35216 20058
rect 35164 19994 35216 20000
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 34794 19136 34850 19145
rect 34794 19071 34850 19080
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34704 18148 34756 18154
rect 34704 18090 34756 18096
rect 34702 18048 34758 18057
rect 34702 17983 34758 17992
rect 34612 17332 34664 17338
rect 34612 17274 34664 17280
rect 34610 17232 34666 17241
rect 34610 17167 34666 17176
rect 34624 15201 34652 17167
rect 34610 15192 34666 15201
rect 34610 15127 34666 15136
rect 34716 14890 34744 17983
rect 34888 17672 34940 17678
rect 34888 17614 34940 17620
rect 34900 17524 34928 17614
rect 34808 17496 34928 17524
rect 34808 16794 34836 17496
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35164 17264 35216 17270
rect 35164 17206 35216 17212
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 35176 16538 35204 17206
rect 35268 16658 35296 21519
rect 35440 21412 35492 21418
rect 35440 21354 35492 21360
rect 35452 20330 35480 21354
rect 35440 20324 35492 20330
rect 35440 20266 35492 20272
rect 35346 19816 35402 19825
rect 35346 19751 35402 19760
rect 35360 17649 35388 19751
rect 35452 19378 35480 20266
rect 35440 19372 35492 19378
rect 35440 19314 35492 19320
rect 35346 17640 35402 17649
rect 35346 17575 35402 17584
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 35256 16652 35308 16658
rect 35256 16594 35308 16600
rect 35176 16510 35296 16538
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35268 16232 35296 16510
rect 35360 16250 35388 17478
rect 35440 16992 35492 16998
rect 35438 16960 35440 16969
rect 35544 16980 35572 21950
rect 35716 21888 35768 21894
rect 35636 21848 35716 21876
rect 35636 21486 35664 21848
rect 35716 21830 35768 21836
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 35636 21146 35664 21422
rect 35714 21176 35770 21185
rect 35624 21140 35676 21146
rect 35714 21111 35770 21120
rect 35624 21082 35676 21088
rect 35728 19961 35756 21111
rect 35714 19952 35770 19961
rect 35714 19887 35770 19896
rect 35716 18964 35768 18970
rect 35716 18906 35768 18912
rect 35624 18624 35676 18630
rect 35624 18566 35676 18572
rect 35492 16960 35572 16980
rect 35494 16952 35572 16960
rect 35438 16895 35494 16904
rect 35440 16448 35492 16454
rect 35440 16390 35492 16396
rect 35176 16204 35296 16232
rect 35348 16244 35400 16250
rect 35176 15892 35204 16204
rect 35348 16186 35400 16192
rect 35452 16046 35480 16390
rect 35530 16280 35586 16289
rect 35530 16215 35586 16224
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35176 15864 35480 15892
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34704 14884 34756 14890
rect 34704 14826 34756 14832
rect 35164 14884 35216 14890
rect 35164 14826 35216 14832
rect 35176 14618 35204 14826
rect 35164 14612 35216 14618
rect 35164 14554 35216 14560
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 35348 13184 35400 13190
rect 35348 13126 35400 13132
rect 34716 12986 34744 13126
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34704 12980 34756 12986
rect 34704 12922 34756 12928
rect 34716 12753 34744 12922
rect 34702 12744 34758 12753
rect 35360 12714 35388 13126
rect 34702 12679 34758 12688
rect 35348 12708 35400 12714
rect 35348 12650 35400 12656
rect 34610 12472 34666 12481
rect 34610 12407 34666 12416
rect 34704 12436 34756 12442
rect 34624 11218 34652 12407
rect 34704 12378 34756 12384
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 34520 11076 34572 11082
rect 34520 11018 34572 11024
rect 34428 10804 34480 10810
rect 34428 10746 34480 10752
rect 34244 10260 34296 10266
rect 34244 10202 34296 10208
rect 34532 10033 34560 11018
rect 34624 10266 34652 11154
rect 34612 10260 34664 10266
rect 34612 10202 34664 10208
rect 34612 10124 34664 10130
rect 34612 10066 34664 10072
rect 34518 10024 34574 10033
rect 34518 9959 34574 9968
rect 34624 9722 34652 10066
rect 33968 9716 34020 9722
rect 33968 9658 34020 9664
rect 34152 9716 34204 9722
rect 34152 9658 34204 9664
rect 34612 9716 34664 9722
rect 34612 9658 34664 9664
rect 33048 9648 33100 9654
rect 33048 9590 33100 9596
rect 33876 9648 33928 9654
rect 33876 9590 33928 9596
rect 32956 9580 33008 9586
rect 32956 9522 33008 9528
rect 33232 9512 33284 9518
rect 33232 9454 33284 9460
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 32968 9110 32996 9318
rect 33244 9178 33272 9454
rect 33232 9172 33284 9178
rect 33232 9114 33284 9120
rect 32680 9104 32732 9110
rect 32680 9046 32732 9052
rect 32956 9104 33008 9110
rect 32956 9046 33008 9052
rect 32036 9036 32088 9042
rect 32036 8978 32088 8984
rect 33324 9036 33376 9042
rect 33324 8978 33376 8984
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 31864 8090 31892 8434
rect 31942 8392 31998 8401
rect 32048 8362 32076 8978
rect 32312 8832 32364 8838
rect 32312 8774 32364 8780
rect 32324 8634 32352 8774
rect 32312 8628 32364 8634
rect 32312 8570 32364 8576
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 31942 8327 31998 8336
rect 32036 8356 32088 8362
rect 31852 8084 31904 8090
rect 31852 8026 31904 8032
rect 31956 7886 31984 8327
rect 32036 8298 32088 8304
rect 31944 7880 31996 7886
rect 31944 7822 31996 7828
rect 31484 7336 31536 7342
rect 31484 7278 31536 7284
rect 31496 6798 31524 7278
rect 31956 7002 31984 7822
rect 32048 7818 32076 8298
rect 32128 8288 32180 8294
rect 32128 8230 32180 8236
rect 32140 8090 32168 8230
rect 32128 8084 32180 8090
rect 32128 8026 32180 8032
rect 32036 7812 32088 7818
rect 32036 7754 32088 7760
rect 32140 7002 32168 8026
rect 32496 7948 32548 7954
rect 32496 7890 32548 7896
rect 32508 7546 32536 7890
rect 32496 7540 32548 7546
rect 32496 7482 32548 7488
rect 32600 7478 32628 8434
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32588 7472 32640 7478
rect 32588 7414 32640 7420
rect 31944 6996 31996 7002
rect 31944 6938 31996 6944
rect 32128 6996 32180 7002
rect 32128 6938 32180 6944
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 31760 6248 31812 6254
rect 31760 6190 31812 6196
rect 31772 5846 31800 6190
rect 32508 5846 32536 6734
rect 32600 6254 32628 7414
rect 32784 6866 32812 8366
rect 33336 8294 33364 8978
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 33704 8634 33732 8910
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 33784 8560 33836 8566
rect 33784 8502 33836 8508
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33324 8288 33376 8294
rect 33324 8230 33376 8236
rect 33336 8090 33364 8230
rect 33704 8090 33732 8366
rect 33324 8084 33376 8090
rect 33324 8026 33376 8032
rect 33692 8084 33744 8090
rect 33692 8026 33744 8032
rect 33232 7540 33284 7546
rect 33232 7482 33284 7488
rect 32772 6860 32824 6866
rect 32772 6802 32824 6808
rect 32784 6458 32812 6802
rect 32772 6452 32824 6458
rect 32772 6394 32824 6400
rect 32588 6248 32640 6254
rect 32588 6190 32640 6196
rect 32784 5914 32812 6394
rect 33244 5914 33272 7482
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33704 6118 33732 6598
rect 33692 6112 33744 6118
rect 33692 6054 33744 6060
rect 32772 5908 32824 5914
rect 32772 5850 32824 5856
rect 33232 5908 33284 5914
rect 33232 5850 33284 5856
rect 31760 5840 31812 5846
rect 31760 5782 31812 5788
rect 32496 5840 32548 5846
rect 32496 5782 32548 5788
rect 33600 5772 33652 5778
rect 33600 5714 33652 5720
rect 33612 5302 33640 5714
rect 33704 5710 33732 6054
rect 33796 5710 33824 8502
rect 33692 5704 33744 5710
rect 33692 5646 33744 5652
rect 33784 5704 33836 5710
rect 33784 5646 33836 5652
rect 33704 5370 33732 5646
rect 33796 5370 33824 5646
rect 33692 5364 33744 5370
rect 33692 5306 33744 5312
rect 33784 5364 33836 5370
rect 33784 5306 33836 5312
rect 33600 5296 33652 5302
rect 33600 5238 33652 5244
rect 31298 3360 31354 3369
rect 31298 3295 31354 3304
rect 33888 2650 33916 9590
rect 33980 9518 34008 9658
rect 34520 9648 34572 9654
rect 34520 9590 34572 9596
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 34334 9208 34390 9217
rect 34334 9143 34336 9152
rect 34388 9143 34390 9152
rect 34336 9114 34388 9120
rect 34348 8974 34376 9114
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 34532 8106 34560 9590
rect 34612 9580 34664 9586
rect 34612 9522 34664 9528
rect 34624 9382 34652 9522
rect 34612 9376 34664 9382
rect 34612 9318 34664 9324
rect 34624 8566 34652 9318
rect 34612 8560 34664 8566
rect 34612 8502 34664 8508
rect 34440 8090 34560 8106
rect 34428 8084 34560 8090
rect 34480 8078 34560 8084
rect 34428 8026 34480 8032
rect 34334 7984 34390 7993
rect 34334 7919 34390 7928
rect 34348 7886 34376 7919
rect 34152 7880 34204 7886
rect 34152 7822 34204 7828
rect 34336 7880 34388 7886
rect 34336 7822 34388 7828
rect 34164 7206 34192 7822
rect 34152 7200 34204 7206
rect 34152 7142 34204 7148
rect 34348 7002 34376 7822
rect 34440 7546 34468 8026
rect 34428 7540 34480 7546
rect 34428 7482 34480 7488
rect 34428 7200 34480 7206
rect 34612 7200 34664 7206
rect 34480 7148 34560 7154
rect 34428 7142 34560 7148
rect 34612 7142 34664 7148
rect 34440 7126 34560 7142
rect 34336 6996 34388 7002
rect 34336 6938 34388 6944
rect 34532 5914 34560 7126
rect 34624 7002 34652 7142
rect 34612 6996 34664 7002
rect 34612 6938 34664 6944
rect 34520 5908 34572 5914
rect 34520 5850 34572 5856
rect 34624 5778 34652 6938
rect 34612 5772 34664 5778
rect 34612 5714 34664 5720
rect 34716 5273 34744 12378
rect 35256 12232 35308 12238
rect 35256 12174 35308 12180
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34808 11830 34836 12038
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34796 11824 34848 11830
rect 34796 11766 34848 11772
rect 35268 11694 35296 12174
rect 35256 11688 35308 11694
rect 35256 11630 35308 11636
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34794 10568 34850 10577
rect 34794 10503 34850 10512
rect 34808 6769 34836 10503
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 35346 9752 35402 9761
rect 35256 9716 35308 9722
rect 35346 9687 35402 9696
rect 35256 9658 35308 9664
rect 35268 9625 35296 9658
rect 35254 9616 35310 9625
rect 35254 9551 35310 9560
rect 35256 9444 35308 9450
rect 35256 9386 35308 9392
rect 35268 8838 35296 9386
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 35268 8362 35296 8774
rect 35256 8356 35308 8362
rect 35256 8298 35308 8304
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34888 7336 34940 7342
rect 34888 7278 34940 7284
rect 34900 6916 34928 7278
rect 35072 6928 35124 6934
rect 34900 6888 35072 6916
rect 34794 6760 34850 6769
rect 34794 6695 34850 6704
rect 34900 6644 34928 6888
rect 35072 6870 35124 6876
rect 34808 6616 34928 6644
rect 34808 6254 34836 6616
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34796 6248 34848 6254
rect 34796 6190 34848 6196
rect 34808 5846 34836 6190
rect 34796 5840 34848 5846
rect 34796 5782 34848 5788
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34702 5264 34758 5273
rect 34702 5199 34758 5208
rect 35360 5114 35388 9687
rect 35452 9081 35480 15864
rect 35544 15065 35572 16215
rect 35530 15056 35586 15065
rect 35530 14991 35586 15000
rect 35532 14816 35584 14822
rect 35532 14758 35584 14764
rect 35544 10266 35572 14758
rect 35532 10260 35584 10266
rect 35532 10202 35584 10208
rect 35636 10198 35664 18566
rect 35728 18426 35756 18906
rect 35716 18420 35768 18426
rect 35716 18362 35768 18368
rect 35716 16720 35768 16726
rect 35716 16662 35768 16668
rect 35728 15706 35756 16662
rect 35716 15700 35768 15706
rect 35716 15642 35768 15648
rect 35820 13530 35848 28970
rect 35912 27849 35940 29106
rect 36360 27872 36412 27878
rect 35898 27840 35954 27849
rect 36360 27814 36412 27820
rect 35898 27775 35954 27784
rect 35912 27606 35940 27775
rect 35900 27600 35952 27606
rect 35900 27542 35952 27548
rect 36372 27538 36400 27814
rect 37004 27600 37056 27606
rect 37004 27542 37056 27548
rect 36360 27532 36412 27538
rect 36360 27474 36412 27480
rect 36372 27130 36400 27474
rect 36820 27328 36872 27334
rect 36820 27270 36872 27276
rect 36360 27124 36412 27130
rect 36360 27066 36412 27072
rect 36372 26926 36400 27066
rect 36636 26988 36688 26994
rect 36636 26930 36688 26936
rect 36360 26920 36412 26926
rect 36360 26862 36412 26868
rect 36450 26072 36506 26081
rect 36450 26007 36506 26016
rect 36360 25152 36412 25158
rect 36360 25094 36412 25100
rect 36372 24954 36400 25094
rect 36360 24948 36412 24954
rect 36360 24890 36412 24896
rect 35900 24812 35952 24818
rect 35900 24754 35952 24760
rect 35912 24342 35940 24754
rect 35900 24336 35952 24342
rect 35900 24278 35952 24284
rect 35912 23866 35940 24278
rect 36464 24274 36492 26007
rect 36648 24954 36676 26930
rect 36832 26790 36860 27270
rect 37016 26994 37044 27542
rect 37004 26988 37056 26994
rect 37004 26930 37056 26936
rect 37016 26874 37044 26930
rect 36924 26846 37044 26874
rect 36820 26784 36872 26790
rect 36820 26726 36872 26732
rect 36832 26450 36860 26726
rect 36820 26444 36872 26450
rect 36820 26386 36872 26392
rect 36924 26314 36952 26846
rect 36912 26308 36964 26314
rect 36912 26250 36964 26256
rect 36820 25696 36872 25702
rect 36820 25638 36872 25644
rect 36832 25401 36860 25638
rect 36818 25392 36874 25401
rect 36818 25327 36874 25336
rect 36636 24948 36688 24954
rect 36636 24890 36688 24896
rect 36924 24410 36952 26250
rect 36912 24404 36964 24410
rect 36912 24346 36964 24352
rect 36452 24268 36504 24274
rect 36452 24210 36504 24216
rect 36464 23866 36492 24210
rect 35900 23860 35952 23866
rect 35900 23802 35952 23808
rect 36452 23860 36504 23866
rect 36452 23802 36504 23808
rect 35992 23588 36044 23594
rect 35992 23530 36044 23536
rect 36004 23322 36032 23530
rect 35992 23316 36044 23322
rect 35992 23258 36044 23264
rect 36636 22500 36688 22506
rect 36636 22442 36688 22448
rect 36268 22432 36320 22438
rect 36082 22400 36138 22409
rect 36268 22374 36320 22380
rect 36082 22335 36138 22344
rect 35900 21344 35952 21350
rect 35900 21286 35952 21292
rect 35912 20398 35940 21286
rect 36096 20602 36124 22335
rect 36280 22166 36308 22374
rect 36268 22160 36320 22166
rect 36268 22102 36320 22108
rect 36648 21690 36676 22442
rect 36636 21684 36688 21690
rect 36636 21626 36688 21632
rect 36174 20904 36230 20913
rect 36174 20839 36230 20848
rect 36084 20596 36136 20602
rect 36084 20538 36136 20544
rect 35900 20392 35952 20398
rect 35900 20334 35952 20340
rect 35912 18834 35940 20334
rect 36084 20256 36136 20262
rect 36084 20198 36136 20204
rect 35992 19916 36044 19922
rect 35992 19858 36044 19864
rect 36004 19310 36032 19858
rect 35992 19304 36044 19310
rect 35990 19272 35992 19281
rect 36044 19272 36046 19281
rect 36096 19242 36124 20198
rect 35990 19207 36046 19216
rect 36084 19236 36136 19242
rect 36004 19181 36032 19207
rect 36084 19178 36136 19184
rect 35900 18828 35952 18834
rect 35900 18770 35952 18776
rect 35912 18426 35940 18770
rect 36096 18766 36124 19178
rect 36188 18902 36216 20839
rect 36912 19848 36964 19854
rect 36912 19790 36964 19796
rect 36924 19174 36952 19790
rect 36912 19168 36964 19174
rect 36912 19110 36964 19116
rect 36176 18896 36228 18902
rect 36176 18838 36228 18844
rect 36084 18760 36136 18766
rect 36084 18702 36136 18708
rect 36188 18426 36216 18838
rect 36542 18728 36598 18737
rect 36542 18663 36598 18672
rect 35900 18420 35952 18426
rect 35900 18362 35952 18368
rect 36176 18420 36228 18426
rect 36176 18362 36228 18368
rect 36556 17746 36584 18663
rect 36544 17740 36596 17746
rect 36544 17682 36596 17688
rect 35992 17536 36044 17542
rect 35992 17478 36044 17484
rect 36084 17536 36136 17542
rect 36084 17478 36136 17484
rect 36004 17202 36032 17478
rect 35992 17196 36044 17202
rect 35992 17138 36044 17144
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35912 15706 35940 16934
rect 36004 16794 36032 17138
rect 35992 16788 36044 16794
rect 35992 16730 36044 16736
rect 35992 16652 36044 16658
rect 35992 16594 36044 16600
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 36004 14822 36032 16594
rect 36096 15881 36124 17478
rect 36556 17338 36584 17682
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 36820 15904 36872 15910
rect 36082 15872 36138 15881
rect 36820 15846 36872 15852
rect 36082 15807 36138 15816
rect 36832 15473 36860 15846
rect 36818 15464 36874 15473
rect 36818 15399 36874 15408
rect 36082 15056 36138 15065
rect 36082 14991 36138 15000
rect 35992 14816 36044 14822
rect 35992 14758 36044 14764
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35716 13320 35768 13326
rect 35716 13262 35768 13268
rect 35728 11626 35756 13262
rect 35716 11620 35768 11626
rect 35716 11562 35768 11568
rect 35716 10260 35768 10266
rect 35716 10202 35768 10208
rect 35624 10192 35676 10198
rect 35624 10134 35676 10140
rect 35532 9988 35584 9994
rect 35532 9930 35584 9936
rect 35544 9382 35572 9930
rect 35622 9752 35678 9761
rect 35622 9687 35678 9696
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35438 9072 35494 9081
rect 35544 9042 35572 9318
rect 35438 9007 35494 9016
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 35544 8650 35572 8978
rect 35452 8634 35572 8650
rect 35440 8628 35572 8634
rect 35492 8622 35572 8628
rect 35440 8570 35492 8576
rect 35440 8424 35492 8430
rect 35440 8366 35492 8372
rect 35452 8022 35480 8366
rect 35440 8016 35492 8022
rect 35440 7958 35492 7964
rect 35452 7342 35480 7958
rect 35440 7336 35492 7342
rect 35440 7278 35492 7284
rect 35440 6248 35492 6254
rect 35440 6190 35492 6196
rect 35452 5846 35480 6190
rect 35532 5908 35584 5914
rect 35532 5850 35584 5856
rect 35440 5840 35492 5846
rect 35440 5782 35492 5788
rect 35452 5302 35480 5782
rect 35544 5370 35572 5850
rect 35532 5364 35584 5370
rect 35532 5306 35584 5312
rect 35440 5296 35492 5302
rect 35440 5238 35492 5244
rect 35360 5086 35480 5114
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 33876 2644 33928 2650
rect 33876 2586 33928 2592
rect 33506 2408 33562 2417
rect 33506 2343 33508 2352
rect 33560 2343 33562 2352
rect 33508 2314 33560 2320
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35452 1737 35480 5086
rect 35636 2961 35664 9687
rect 35728 4185 35756 10202
rect 35714 4176 35770 4185
rect 35714 4111 35770 4120
rect 35622 2952 35678 2961
rect 35622 2887 35678 2896
rect 35438 1728 35494 1737
rect 35438 1663 35494 1672
rect 35820 649 35848 13466
rect 35992 12640 36044 12646
rect 35992 12582 36044 12588
rect 36004 12374 36032 12582
rect 35992 12368 36044 12374
rect 35992 12310 36044 12316
rect 36004 11898 36032 12310
rect 35992 11892 36044 11898
rect 35992 11834 36044 11840
rect 36096 11286 36124 14991
rect 36544 13388 36596 13394
rect 36544 13330 36596 13336
rect 36452 13320 36504 13326
rect 36452 13262 36504 13268
rect 36268 13184 36320 13190
rect 36268 13126 36320 13132
rect 36280 12306 36308 13126
rect 36464 12986 36492 13262
rect 36452 12980 36504 12986
rect 36452 12922 36504 12928
rect 36556 12918 36584 13330
rect 36820 12980 36872 12986
rect 36820 12922 36872 12928
rect 36544 12912 36596 12918
rect 36544 12854 36596 12860
rect 36542 12744 36598 12753
rect 36542 12679 36598 12688
rect 36268 12300 36320 12306
rect 36268 12242 36320 12248
rect 36280 11898 36308 12242
rect 36268 11892 36320 11898
rect 36268 11834 36320 11840
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36266 11520 36322 11529
rect 36266 11455 36322 11464
rect 36084 11280 36136 11286
rect 36084 11222 36136 11228
rect 35992 11008 36044 11014
rect 35992 10950 36044 10956
rect 36004 10606 36032 10950
rect 35992 10600 36044 10606
rect 35992 10542 36044 10548
rect 35900 9920 35952 9926
rect 35900 9862 35952 9868
rect 35912 9722 35940 9862
rect 35900 9716 35952 9722
rect 35900 9658 35952 9664
rect 35898 9616 35954 9625
rect 35898 9551 35954 9560
rect 35912 7857 35940 9551
rect 36004 9110 36032 10542
rect 36096 10266 36124 11222
rect 36176 11212 36228 11218
rect 36176 11154 36228 11160
rect 36188 10538 36216 11154
rect 36176 10532 36228 10538
rect 36176 10474 36228 10480
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 36280 10130 36308 11455
rect 36464 11354 36492 11630
rect 36452 11348 36504 11354
rect 36452 11290 36504 11296
rect 36556 10130 36584 12679
rect 36832 12442 36860 12922
rect 36820 12436 36872 12442
rect 36820 12378 36872 12384
rect 36832 12345 36860 12378
rect 36818 12336 36874 12345
rect 36818 12271 36874 12280
rect 36636 11552 36688 11558
rect 36636 11494 36688 11500
rect 36648 10713 36676 11494
rect 36634 10704 36690 10713
rect 36634 10639 36690 10648
rect 36924 10305 36952 19110
rect 37108 18630 37136 34478
rect 37464 27940 37516 27946
rect 37464 27882 37516 27888
rect 37186 27296 37242 27305
rect 37186 27231 37242 27240
rect 37200 24818 37228 27231
rect 37476 27130 37504 27882
rect 37464 27124 37516 27130
rect 37464 27066 37516 27072
rect 37188 24812 37240 24818
rect 37188 24754 37240 24760
rect 37280 20256 37332 20262
rect 37280 20198 37332 20204
rect 37188 18964 37240 18970
rect 37292 18952 37320 20198
rect 37240 18924 37320 18952
rect 37188 18906 37240 18912
rect 37096 18624 37148 18630
rect 37096 18566 37148 18572
rect 37186 13968 37242 13977
rect 37186 13903 37242 13912
rect 37096 10464 37148 10470
rect 37096 10406 37148 10412
rect 36910 10296 36966 10305
rect 36910 10231 36966 10240
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 36544 10124 36596 10130
rect 36544 10066 36596 10072
rect 36280 9654 36308 10066
rect 36556 9722 36584 10066
rect 36728 9920 36780 9926
rect 36728 9862 36780 9868
rect 36544 9716 36596 9722
rect 36544 9658 36596 9664
rect 36268 9648 36320 9654
rect 36268 9590 36320 9596
rect 35992 9104 36044 9110
rect 35992 9046 36044 9052
rect 36004 8430 36032 9046
rect 35992 8424 36044 8430
rect 35992 8366 36044 8372
rect 36636 8288 36688 8294
rect 36636 8230 36688 8236
rect 36648 8090 36676 8230
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36740 7993 36768 9862
rect 36912 9376 36964 9382
rect 36912 9318 36964 9324
rect 36924 9217 36952 9318
rect 36910 9208 36966 9217
rect 37108 9178 37136 10406
rect 37200 9654 37228 13903
rect 37556 13252 37608 13258
rect 37556 13194 37608 13200
rect 37568 12986 37596 13194
rect 37556 12980 37608 12986
rect 37556 12922 37608 12928
rect 37188 9648 37240 9654
rect 37188 9590 37240 9596
rect 36910 9143 36966 9152
rect 37096 9172 37148 9178
rect 37096 9114 37148 9120
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 36832 8634 36860 8978
rect 36820 8628 36872 8634
rect 36820 8570 36872 8576
rect 37096 8288 37148 8294
rect 37096 8230 37148 8236
rect 36726 7984 36782 7993
rect 36544 7948 36596 7954
rect 36726 7919 36782 7928
rect 36544 7890 36596 7896
rect 35898 7848 35954 7857
rect 35898 7783 35954 7792
rect 36556 7206 36584 7890
rect 37108 7546 37136 8230
rect 37096 7540 37148 7546
rect 37096 7482 37148 7488
rect 35900 7200 35952 7206
rect 35900 7142 35952 7148
rect 36544 7200 36596 7206
rect 36544 7142 36596 7148
rect 35912 6254 35940 7142
rect 36556 6458 36584 7142
rect 37108 6458 37136 7482
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 37096 6452 37148 6458
rect 37096 6394 37148 6400
rect 35900 6248 35952 6254
rect 35900 6190 35952 6196
rect 36556 5914 36584 6394
rect 36544 5908 36596 5914
rect 36544 5850 36596 5856
rect 36636 2508 36688 2514
rect 36636 2450 36688 2456
rect 35806 640 35862 649
rect 35806 575 35862 584
rect 36648 480 36676 2450
rect 3330 0 3386 480
rect 9954 0 10010 480
rect 16670 0 16726 480
rect 23294 0 23350 480
rect 30010 0 30066 480
rect 36634 0 36690 480
<< via2 >>
rect 2042 35128 2098 35184
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4710 35400 4766 35456
rect 7470 36524 7472 36544
rect 7472 36524 7524 36544
rect 7524 36524 7526 36544
rect 7470 36488 7526 36524
rect 7102 35672 7158 35728
rect 6090 35264 6146 35320
rect 4618 34992 4674 35048
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 3146 34604 3202 34640
rect 3146 34584 3148 34604
rect 3148 34584 3200 34604
rect 3200 34584 3202 34604
rect 2870 34076 2872 34096
rect 2872 34076 2924 34096
rect 2924 34076 2926 34096
rect 2870 34040 2926 34076
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4066 31864 4122 31920
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 1674 30660 1730 30696
rect 1674 30640 1676 30660
rect 1676 30640 1728 30660
rect 1728 30640 1730 30660
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 5630 31884 5686 31920
rect 5630 31864 5632 31884
rect 5632 31864 5684 31884
rect 5684 31864 5686 31884
rect 7746 35828 7802 35864
rect 7746 35808 7748 35828
rect 7748 35808 7800 35828
rect 7800 35808 7802 35828
rect 9402 35808 9458 35864
rect 9586 35808 9642 35864
rect 8850 35556 8906 35592
rect 8850 35536 8852 35556
rect 8852 35536 8904 35556
rect 8904 35536 8906 35556
rect 10506 35672 10562 35728
rect 10690 35672 10746 35728
rect 9586 35400 9642 35456
rect 9126 34740 9182 34776
rect 9126 34720 9128 34740
rect 9128 34720 9180 34740
rect 9180 34720 9182 34740
rect 9586 34348 9588 34368
rect 9588 34348 9640 34368
rect 9640 34348 9642 34368
rect 9586 34312 9642 34348
rect 10782 33532 10784 33552
rect 10784 33532 10836 33552
rect 10836 33532 10838 33552
rect 10782 33496 10838 33532
rect 11242 34312 11298 34368
rect 12714 35672 12770 35728
rect 11610 34720 11666 34776
rect 11610 34040 11666 34096
rect 9862 32544 9918 32600
rect 5906 30640 5962 30696
rect 7010 30660 7066 30696
rect 7010 30640 7012 30660
rect 7012 30640 7064 30660
rect 7064 30640 7066 30660
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 13634 34856 13690 34912
rect 12622 33904 12678 33960
rect 12806 33496 12862 33552
rect 12898 33224 12954 33280
rect 13266 32564 13322 32600
rect 13266 32544 13268 32564
rect 13268 32544 13320 32564
rect 13320 32544 13322 32564
rect 11886 31476 11942 31512
rect 11886 31456 11888 31476
rect 11888 31456 11940 31476
rect 11940 31456 11942 31476
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 8206 27784 8262 27840
rect 11150 30912 11206 30968
rect 10782 30368 10838 30424
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 7654 24520 7710 24576
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 10230 27820 10232 27840
rect 10232 27820 10284 27840
rect 10284 27820 10286 27840
rect 10230 27784 10286 27820
rect 10138 27512 10194 27568
rect 12714 31048 12770 31104
rect 12714 30368 12770 30424
rect 13726 30388 13782 30424
rect 13726 30368 13728 30388
rect 13728 30368 13780 30388
rect 13780 30368 13782 30388
rect 14186 34740 14242 34776
rect 14186 34720 14188 34740
rect 14188 34720 14240 34740
rect 14240 34720 14242 34740
rect 14094 32852 14096 32872
rect 14096 32852 14148 32872
rect 14148 32852 14150 32872
rect 14094 32816 14150 32852
rect 14922 32428 14978 32464
rect 15658 35708 15660 35728
rect 15660 35708 15712 35728
rect 15712 35708 15714 35728
rect 15658 35672 15714 35708
rect 15290 35128 15346 35184
rect 15750 34856 15806 34912
rect 16854 35012 16910 35048
rect 16854 34992 16856 35012
rect 16856 34992 16908 35012
rect 16908 34992 16910 35012
rect 16118 34720 16174 34776
rect 15658 33496 15714 33552
rect 15934 33516 15990 33552
rect 15934 33496 15936 33516
rect 15936 33496 15988 33516
rect 15988 33496 15990 33516
rect 16026 33224 16082 33280
rect 14922 32408 14924 32428
rect 14924 32408 14976 32428
rect 14976 32408 14978 32428
rect 14830 31456 14886 31512
rect 14370 30932 14426 30968
rect 14370 30912 14372 30932
rect 14372 30912 14424 30932
rect 14424 30912 14426 30932
rect 12714 27512 12770 27568
rect 10414 26288 10470 26344
rect 12530 26308 12586 26344
rect 12530 26288 12532 26308
rect 12532 26288 12584 26308
rect 12584 26288 12586 26308
rect 15474 31048 15530 31104
rect 16762 32816 16818 32872
rect 16670 32408 16726 32464
rect 16486 31592 16542 31648
rect 17958 35264 18014 35320
rect 17958 34856 18014 34912
rect 17038 33260 17040 33280
rect 17040 33260 17092 33280
rect 17092 33260 17094 33280
rect 17038 33224 17094 33260
rect 17590 32544 17646 32600
rect 17038 31476 17094 31512
rect 17038 31456 17040 31476
rect 17040 31456 17092 31476
rect 17092 31456 17094 31476
rect 18142 34620 18144 34640
rect 18144 34620 18196 34640
rect 18196 34620 18198 34640
rect 18142 34584 18198 34620
rect 16946 30368 17002 30424
rect 15842 29588 15844 29608
rect 15844 29588 15896 29608
rect 15896 29588 15898 29608
rect 15842 29552 15898 29588
rect 17038 27512 17094 27568
rect 8482 24792 8538 24848
rect 9218 24792 9274 24848
rect 11886 24812 11942 24848
rect 11886 24792 11888 24812
rect 11888 24792 11940 24812
rect 11940 24792 11942 24812
rect 12898 24828 12900 24848
rect 12900 24828 12952 24848
rect 12952 24828 12954 24848
rect 12898 24792 12954 24828
rect 11518 24556 11520 24576
rect 11520 24556 11572 24576
rect 11572 24556 11574 24576
rect 11518 24520 11574 24556
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 12714 23432 12770 23488
rect 12990 22888 13046 22944
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 12806 21936 12862 21992
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 14738 26424 14794 26480
rect 16394 24520 16450 24576
rect 15290 23568 15346 23624
rect 16486 23432 16542 23488
rect 16394 22924 16396 22944
rect 16396 22924 16448 22944
rect 16448 22924 16450 22944
rect 16394 22888 16450 22924
rect 14002 21936 14058 21992
rect 18970 34856 19026 34912
rect 18878 31456 18934 31512
rect 18878 29552 18934 29608
rect 19154 34740 19210 34776
rect 19154 34720 19156 34740
rect 19156 34720 19208 34740
rect 19208 34720 19210 34740
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 20258 35944 20314 36000
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 21178 35808 21234 35864
rect 20994 35264 21050 35320
rect 20534 34720 20590 34776
rect 20074 34196 20130 34232
rect 20074 34176 20076 34196
rect 20076 34176 20128 34196
rect 20128 34176 20130 34196
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19430 31592 19486 31648
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 20166 32564 20222 32600
rect 20166 32544 20168 32564
rect 20168 32544 20220 32564
rect 20220 32544 20222 32564
rect 21178 34720 21234 34776
rect 20626 30776 20682 30832
rect 22282 35980 22284 36000
rect 22284 35980 22336 36000
rect 22336 35980 22338 36000
rect 22282 35944 22338 35980
rect 22650 35264 22706 35320
rect 19890 27512 19946 27568
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 18602 24928 18658 24984
rect 18694 24792 18750 24848
rect 2778 20032 2834 20088
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 18694 24556 18696 24576
rect 18696 24556 18748 24576
rect 18748 24556 18750 24576
rect 18694 24520 18750 24556
rect 18050 23604 18052 23624
rect 18052 23604 18104 23624
rect 18104 23604 18106 23624
rect 18050 23568 18106 23604
rect 20166 26424 20222 26480
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19982 24248 20038 24304
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 570 6704 626 6760
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 23754 35536 23810 35592
rect 23570 34196 23626 34232
rect 23570 34176 23572 34196
rect 23572 34176 23624 34196
rect 23624 34176 23626 34196
rect 22558 30796 22614 30832
rect 22558 30776 22560 30796
rect 22560 30776 22612 30796
rect 22612 30776 22614 30796
rect 20626 25472 20682 25528
rect 20718 24928 20774 24984
rect 20902 24828 20904 24848
rect 20904 24828 20956 24848
rect 20956 24828 20958 24848
rect 20902 24792 20958 24828
rect 21822 28872 21878 28928
rect 23662 28872 23718 28928
rect 24950 34720 25006 34776
rect 24858 32952 24914 33008
rect 24766 31204 24822 31240
rect 24766 31184 24768 31204
rect 24768 31184 24820 31204
rect 24820 31184 24822 31204
rect 24398 30232 24454 30288
rect 24766 29280 24822 29336
rect 23846 26288 23902 26344
rect 22006 25472 22062 25528
rect 23662 25492 23718 25528
rect 23662 25472 23664 25492
rect 23664 25472 23716 25492
rect 23716 25472 23718 25492
rect 21362 24248 21418 24304
rect 25226 31884 25282 31920
rect 25226 31864 25228 31884
rect 25228 31864 25280 31884
rect 25280 31864 25282 31884
rect 27250 35672 27306 35728
rect 29458 35128 29514 35184
rect 27526 33904 27582 33960
rect 27526 33632 27582 33688
rect 35622 39344 35678 39400
rect 32770 34992 32826 35048
rect 33874 34992 33930 35048
rect 31666 34584 31722 34640
rect 30562 33904 30618 33960
rect 30194 33496 30250 33552
rect 29366 32972 29422 33008
rect 29366 32952 29368 32972
rect 29368 32952 29420 32972
rect 29420 32952 29422 32972
rect 29550 31864 29606 31920
rect 28170 31184 28226 31240
rect 26974 30232 27030 30288
rect 26422 29300 26478 29336
rect 26422 29280 26424 29300
rect 26424 29280 26476 29300
rect 26476 29280 26478 29300
rect 25870 28056 25926 28112
rect 27894 28056 27950 28112
rect 24214 26152 24270 26208
rect 25594 26288 25650 26344
rect 26238 26324 26240 26344
rect 26240 26324 26292 26344
rect 26292 26324 26294 26344
rect 26238 26288 26294 26324
rect 26238 25492 26294 25528
rect 26974 26152 27030 26208
rect 26238 25472 26240 25492
rect 26240 25472 26292 25492
rect 26292 25472 26294 25492
rect 26606 25064 26662 25120
rect 25042 24792 25098 24848
rect 28446 26288 28502 26344
rect 27802 24928 27858 24984
rect 28722 25064 28778 25120
rect 21546 22752 21602 22808
rect 20166 20712 20222 20768
rect 19522 20304 19578 20360
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 21362 20032 21418 20088
rect 22190 20304 22246 20360
rect 19246 18264 19302 18320
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19246 17176 19302 17232
rect 19246 17040 19302 17096
rect 20074 18148 20130 18184
rect 20074 18128 20076 18148
rect 20076 18128 20128 18148
rect 20128 18128 20130 18148
rect 20350 17992 20406 18048
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 21086 18128 21142 18184
rect 21546 17312 21602 17368
rect 21730 17060 21786 17096
rect 21730 17040 21732 17060
rect 21732 17040 21784 17060
rect 21784 17040 21786 17060
rect 20258 16632 20314 16688
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 22374 18264 22430 18320
rect 22282 17992 22338 18048
rect 23662 20052 23718 20088
rect 23662 20032 23664 20052
rect 23664 20032 23716 20052
rect 23716 20032 23718 20052
rect 23754 19216 23810 19272
rect 23846 18164 23848 18184
rect 23848 18164 23900 18184
rect 23900 18164 23902 18184
rect 23846 18128 23902 18164
rect 22282 17176 22338 17232
rect 22282 16632 22338 16688
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 21178 12824 21234 12880
rect 23294 14728 23350 14784
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 570 5616 626 5672
rect 17498 5616 17554 5672
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 24490 22480 24546 22536
rect 24674 21548 24730 21584
rect 24674 21528 24676 21548
rect 24676 21528 24728 21548
rect 24728 21528 24730 21548
rect 25686 22772 25742 22808
rect 25686 22752 25688 22772
rect 25688 22752 25740 22772
rect 25740 22752 25742 22772
rect 24306 20460 24362 20496
rect 24306 20440 24308 20460
rect 24308 20440 24360 20460
rect 24360 20440 24362 20460
rect 24214 19352 24270 19408
rect 24030 18944 24086 19000
rect 24490 19352 24546 19408
rect 26882 22516 26884 22536
rect 26884 22516 26936 22536
rect 26936 22516 26938 22536
rect 26882 22480 26938 22516
rect 26698 21528 26754 21584
rect 26054 20204 26056 20224
rect 26056 20204 26108 20224
rect 26108 20204 26110 20224
rect 26054 20168 26110 20204
rect 26514 19916 26570 19952
rect 26514 19896 26516 19916
rect 26516 19896 26568 19916
rect 26568 19896 26570 19916
rect 25778 19116 25780 19136
rect 25780 19116 25832 19136
rect 25832 19116 25834 19136
rect 25778 19080 25834 19116
rect 27710 20712 27766 20768
rect 27618 20596 27674 20632
rect 27618 20576 27620 20596
rect 27620 20576 27672 20596
rect 27672 20576 27674 20596
rect 26882 19252 26884 19272
rect 26884 19252 26936 19272
rect 26936 19252 26938 19272
rect 26882 19216 26938 19252
rect 26698 18964 26754 19000
rect 26698 18944 26700 18964
rect 26700 18944 26752 18964
rect 26752 18944 26754 18964
rect 27066 18944 27122 19000
rect 25226 17856 25282 17912
rect 28446 21936 28502 21992
rect 28906 23976 28962 24032
rect 27986 20440 28042 20496
rect 25226 17332 25282 17368
rect 25226 17312 25228 17332
rect 25228 17312 25280 17332
rect 25280 17312 25282 17332
rect 25502 17060 25558 17096
rect 25502 17040 25504 17060
rect 25504 17040 25556 17060
rect 25556 17040 25558 17060
rect 27434 16904 27490 16960
rect 24030 12824 24086 12880
rect 25134 13640 25190 13696
rect 24766 12980 24822 13016
rect 24766 12960 24768 12980
rect 24768 12960 24820 12980
rect 24820 12960 24822 12980
rect 27710 15816 27766 15872
rect 27066 14764 27068 14784
rect 27068 14764 27120 14784
rect 27120 14764 27122 14784
rect 27066 14728 27122 14764
rect 26146 12960 26202 13016
rect 28998 20052 29054 20088
rect 28998 20032 29000 20052
rect 29000 20032 29052 20052
rect 29052 20032 29054 20052
rect 27894 17876 27950 17912
rect 27894 17856 27896 17876
rect 27896 17856 27948 17876
rect 27948 17856 27950 17876
rect 28722 17584 28778 17640
rect 28630 15680 28686 15736
rect 28446 15156 28502 15192
rect 28446 15136 28448 15156
rect 28448 15136 28500 15156
rect 28500 15136 28502 15156
rect 28998 16940 29000 16960
rect 29000 16940 29052 16960
rect 29052 16940 29054 16960
rect 28998 16904 29054 16940
rect 29458 20168 29514 20224
rect 29366 19488 29422 19544
rect 30102 20168 30158 20224
rect 29918 18964 29974 19000
rect 29918 18944 29920 18964
rect 29920 18944 29972 18964
rect 29972 18944 29974 18964
rect 29090 15000 29146 15056
rect 28538 13640 28594 13696
rect 28998 13640 29054 13696
rect 24582 9696 24638 9752
rect 27618 11736 27674 11792
rect 30010 12300 30066 12336
rect 30010 12280 30012 12300
rect 30012 12280 30064 12300
rect 30064 12280 30066 12300
rect 27250 9696 27306 9752
rect 29918 8336 29974 8392
rect 31666 27240 31722 27296
rect 31574 26424 31630 26480
rect 31298 26324 31300 26344
rect 31300 26324 31352 26344
rect 31352 26324 31354 26344
rect 31298 26288 31354 26324
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 35806 36896 35862 36952
rect 35622 35672 35678 35728
rect 35530 35284 35586 35320
rect 35530 35264 35532 35284
rect 35532 35264 35584 35284
rect 35584 35264 35586 35284
rect 34794 34856 34850 34912
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 35438 34584 35494 34640
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 33782 27820 33784 27840
rect 33784 27820 33836 27840
rect 33836 27820 33838 27840
rect 33782 27784 33838 27820
rect 33230 27276 33232 27296
rect 33232 27276 33284 27296
rect 33284 27276 33286 27296
rect 33230 27240 33286 27276
rect 33230 26424 33286 26480
rect 32034 24928 32090 24984
rect 31942 23976 31998 24032
rect 31022 20168 31078 20224
rect 34058 25336 34114 25392
rect 34518 28056 34574 28112
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34518 23704 34574 23760
rect 31758 20032 31814 20088
rect 33230 20848 33286 20904
rect 33322 20204 33324 20224
rect 33324 20204 33376 20224
rect 33376 20204 33378 20224
rect 33322 20168 33378 20204
rect 30286 15308 30288 15328
rect 30288 15308 30340 15328
rect 30340 15308 30342 15328
rect 30286 15272 30342 15308
rect 31390 17060 31446 17096
rect 31390 17040 31392 17060
rect 31392 17040 31444 17060
rect 31444 17040 31446 17060
rect 30562 15680 30618 15736
rect 30378 11736 30434 11792
rect 32678 18028 32680 18048
rect 32680 18028 32732 18048
rect 32732 18028 32734 18048
rect 32678 17992 32734 18028
rect 31850 15408 31906 15464
rect 32770 15272 32826 15328
rect 33782 19236 33838 19272
rect 33782 19216 33784 19236
rect 33784 19216 33836 19236
rect 33836 19216 33838 19236
rect 32954 15408 33010 15464
rect 31206 11600 31262 11656
rect 31666 11620 31722 11656
rect 31666 11600 31668 11620
rect 31668 11600 31720 11620
rect 31720 11600 31722 11620
rect 23294 3984 23350 4040
rect 23938 3984 23994 4040
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 16670 3304 16726 3360
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 3330 2352 3386 2408
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 35254 23568 35310 23624
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 35254 21936 35310 21992
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34242 19488 34298 19544
rect 33046 10668 33102 10704
rect 31574 9152 31630 9208
rect 33046 10648 33048 10668
rect 33048 10648 33100 10668
rect 33100 10648 33102 10668
rect 36726 38120 36782 38176
rect 36082 35536 36138 35592
rect 38290 35264 38346 35320
rect 37186 35128 37242 35184
rect 39394 34584 39450 34640
rect 35806 34448 35862 34504
rect 35714 33496 35770 33552
rect 35622 33224 35678 33280
rect 35714 32000 35770 32056
rect 35898 30776 35954 30832
rect 35530 29552 35586 29608
rect 35254 21528 35310 21584
rect 35438 21528 35494 21584
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34794 19080 34850 19136
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34702 17992 34758 18048
rect 34610 17176 34666 17232
rect 34610 15136 34666 15192
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35346 19760 35402 19816
rect 35346 17584 35402 17640
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 35714 21120 35770 21176
rect 35714 19896 35770 19952
rect 35438 16940 35440 16960
rect 35440 16940 35492 16960
rect 35492 16940 35494 16960
rect 35438 16904 35494 16940
rect 35530 16224 35586 16280
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34702 12688 34758 12744
rect 34610 12416 34666 12472
rect 34518 9968 34574 10024
rect 31942 8336 31998 8392
rect 31298 3304 31354 3360
rect 34334 9172 34390 9208
rect 34334 9152 34336 9172
rect 34336 9152 34388 9172
rect 34388 9152 34390 9172
rect 34334 7928 34390 7984
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34794 10512 34850 10568
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 35346 9696 35402 9752
rect 35254 9560 35310 9616
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34794 6704 34850 6760
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34702 5208 34758 5264
rect 35530 15000 35586 15056
rect 35898 27784 35954 27840
rect 36450 26016 36506 26072
rect 36818 25336 36874 25392
rect 36082 22344 36138 22400
rect 36174 20848 36230 20904
rect 35990 19252 35992 19272
rect 35992 19252 36044 19272
rect 36044 19252 36046 19272
rect 35990 19216 36046 19252
rect 36542 18672 36598 18728
rect 36082 15816 36138 15872
rect 36818 15408 36874 15464
rect 36082 15000 36138 15056
rect 35622 9696 35678 9752
rect 35438 9016 35494 9072
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 33506 2372 33562 2408
rect 33506 2352 33508 2372
rect 33508 2352 33560 2372
rect 33560 2352 33562 2372
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 35714 4120 35770 4176
rect 35622 2896 35678 2952
rect 35438 1672 35494 1728
rect 36542 12688 36598 12744
rect 36266 11464 36322 11520
rect 35898 9560 35954 9616
rect 36818 12280 36874 12336
rect 36634 10648 36690 10704
rect 37186 27240 37242 27296
rect 37186 13912 37242 13968
rect 36910 10240 36966 10296
rect 36910 9152 36966 9208
rect 36726 7928 36782 7984
rect 35898 7792 35954 7848
rect 35806 584 35862 640
<< metal3 >>
rect 35617 39402 35683 39405
rect 39520 39402 40000 39432
rect 35617 39400 40000 39402
rect 35617 39344 35622 39400
rect 35678 39344 40000 39400
rect 35617 39342 40000 39344
rect 35617 39339 35683 39342
rect 39520 39312 40000 39342
rect 36721 38178 36787 38181
rect 39520 38178 40000 38208
rect 36721 38176 40000 38178
rect 36721 38120 36726 38176
rect 36782 38120 40000 38176
rect 36721 38118 40000 38120
rect 36721 38115 36787 38118
rect 39520 38088 40000 38118
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 35801 36954 35867 36957
rect 39520 36954 40000 36984
rect 35801 36952 40000 36954
rect 35801 36896 35806 36952
rect 35862 36896 40000 36952
rect 35801 36894 40000 36896
rect 35801 36891 35867 36894
rect 39520 36864 40000 36894
rect 7465 36546 7531 36549
rect 8150 36546 8156 36548
rect 7465 36544 8156 36546
rect 7465 36488 7470 36544
rect 7526 36488 8156 36544
rect 7465 36486 8156 36488
rect 7465 36483 7531 36486
rect 8150 36484 8156 36486
rect 8220 36484 8226 36548
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 20253 36002 20319 36005
rect 22277 36002 22343 36005
rect 20253 36000 22343 36002
rect 20253 35944 20258 36000
rect 20314 35944 22282 36000
rect 22338 35944 22343 36000
rect 20253 35942 22343 35944
rect 20253 35939 20319 35942
rect 22277 35939 22343 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 7741 35866 7807 35869
rect 9397 35866 9463 35869
rect 7741 35864 9463 35866
rect 7741 35808 7746 35864
rect 7802 35808 9402 35864
rect 9458 35808 9463 35864
rect 7741 35806 9463 35808
rect 7741 35803 7807 35806
rect 9397 35803 9463 35806
rect 9581 35866 9647 35869
rect 21173 35866 21239 35869
rect 9581 35864 21239 35866
rect 9581 35808 9586 35864
rect 9642 35808 21178 35864
rect 21234 35808 21239 35864
rect 9581 35806 21239 35808
rect 9581 35803 9647 35806
rect 21173 35803 21239 35806
rect 7097 35730 7163 35733
rect 10501 35730 10567 35733
rect 7097 35728 10567 35730
rect 7097 35672 7102 35728
rect 7158 35672 10506 35728
rect 10562 35672 10567 35728
rect 7097 35670 10567 35672
rect 7097 35667 7163 35670
rect 10501 35667 10567 35670
rect 10685 35730 10751 35733
rect 12709 35730 12775 35733
rect 10685 35728 12775 35730
rect 10685 35672 10690 35728
rect 10746 35672 12714 35728
rect 12770 35672 12775 35728
rect 10685 35670 12775 35672
rect 10685 35667 10751 35670
rect 12709 35667 12775 35670
rect 15653 35730 15719 35733
rect 27245 35730 27311 35733
rect 15653 35728 27311 35730
rect 15653 35672 15658 35728
rect 15714 35672 27250 35728
rect 27306 35672 27311 35728
rect 15653 35670 27311 35672
rect 15653 35667 15719 35670
rect 27245 35667 27311 35670
rect 35617 35730 35683 35733
rect 39520 35730 40000 35760
rect 35617 35728 40000 35730
rect 35617 35672 35622 35728
rect 35678 35672 40000 35728
rect 35617 35670 40000 35672
rect 35617 35667 35683 35670
rect 39520 35640 40000 35670
rect 8845 35594 8911 35597
rect 23749 35594 23815 35597
rect 8845 35592 24778 35594
rect 8845 35536 8850 35592
rect 8906 35536 23754 35592
rect 23810 35536 24778 35592
rect 8845 35534 24778 35536
rect 8845 35531 8911 35534
rect 23749 35531 23815 35534
rect 4705 35458 4771 35461
rect 9581 35458 9647 35461
rect 4705 35456 9647 35458
rect 4705 35400 4710 35456
rect 4766 35400 9586 35456
rect 9642 35400 9647 35456
rect 4705 35398 9647 35400
rect 4705 35395 4771 35398
rect 9581 35395 9647 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 6085 35322 6151 35325
rect 17953 35322 18019 35325
rect 6085 35320 18019 35322
rect 6085 35264 6090 35320
rect 6146 35264 17958 35320
rect 18014 35264 18019 35320
rect 6085 35262 18019 35264
rect 6085 35259 6151 35262
rect 17953 35259 18019 35262
rect 20989 35322 21055 35325
rect 22645 35322 22711 35325
rect 20989 35320 22711 35322
rect 20989 35264 20994 35320
rect 21050 35264 22650 35320
rect 22706 35264 22711 35320
rect 20989 35262 22711 35264
rect 24718 35322 24778 35534
rect 24894 35532 24900 35596
rect 24964 35594 24970 35596
rect 36077 35594 36143 35597
rect 24964 35592 36143 35594
rect 24964 35536 36082 35592
rect 36138 35536 36143 35592
rect 24964 35534 36143 35536
rect 24964 35532 24970 35534
rect 36077 35531 36143 35534
rect 35525 35322 35591 35325
rect 38285 35322 38351 35325
rect 24718 35262 29746 35322
rect 20989 35259 21055 35262
rect 22645 35259 22711 35262
rect 2037 35186 2103 35189
rect 15285 35186 15351 35189
rect 29453 35186 29519 35189
rect 2037 35184 29519 35186
rect 2037 35128 2042 35184
rect 2098 35128 15290 35184
rect 15346 35128 29458 35184
rect 29514 35128 29519 35184
rect 2037 35126 29519 35128
rect 29686 35186 29746 35262
rect 35525 35320 38351 35322
rect 35525 35264 35530 35320
rect 35586 35264 38290 35320
rect 38346 35264 38351 35320
rect 35525 35262 38351 35264
rect 35525 35259 35591 35262
rect 38285 35259 38351 35262
rect 37181 35186 37247 35189
rect 29686 35184 37247 35186
rect 29686 35128 37186 35184
rect 37242 35128 37247 35184
rect 29686 35126 37247 35128
rect 2037 35123 2103 35126
rect 15285 35123 15351 35126
rect 29453 35123 29519 35126
rect 37181 35123 37247 35126
rect 4613 35050 4679 35053
rect 16849 35050 16915 35053
rect 32765 35050 32831 35053
rect 4613 35048 32831 35050
rect 4613 34992 4618 35048
rect 4674 34992 16854 35048
rect 16910 34992 32770 35048
rect 32826 34992 32831 35048
rect 4613 34990 32831 34992
rect 4613 34987 4679 34990
rect 16849 34987 16915 34990
rect 32765 34987 32831 34990
rect 33174 34988 33180 35052
rect 33244 35050 33250 35052
rect 33869 35050 33935 35053
rect 33244 35048 33935 35050
rect 33244 34992 33874 35048
rect 33930 34992 33935 35048
rect 33244 34990 33935 34992
rect 33244 34988 33250 34990
rect 33869 34987 33935 34990
rect 13629 34914 13695 34917
rect 15745 34914 15811 34917
rect 13629 34912 15811 34914
rect 13629 34856 13634 34912
rect 13690 34856 15750 34912
rect 15806 34856 15811 34912
rect 13629 34854 15811 34856
rect 13629 34851 13695 34854
rect 15745 34851 15811 34854
rect 17953 34914 18019 34917
rect 18965 34914 19031 34917
rect 34789 34914 34855 34917
rect 17953 34912 34855 34914
rect 17953 34856 17958 34912
rect 18014 34856 18970 34912
rect 19026 34856 34794 34912
rect 34850 34856 34855 34912
rect 17953 34854 34855 34856
rect 17953 34851 18019 34854
rect 18965 34851 19031 34854
rect 34789 34851 34855 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 9121 34778 9187 34781
rect 11605 34778 11671 34781
rect 9121 34776 11671 34778
rect 9121 34720 9126 34776
rect 9182 34720 11610 34776
rect 11666 34720 11671 34776
rect 9121 34718 11671 34720
rect 9121 34715 9187 34718
rect 11605 34715 11671 34718
rect 14181 34778 14247 34781
rect 16113 34778 16179 34781
rect 14181 34776 16179 34778
rect 14181 34720 14186 34776
rect 14242 34720 16118 34776
rect 16174 34720 16179 34776
rect 14181 34718 16179 34720
rect 14181 34715 14247 34718
rect 16113 34715 16179 34718
rect 19149 34778 19215 34781
rect 20529 34778 20595 34781
rect 19149 34776 20595 34778
rect 19149 34720 19154 34776
rect 19210 34720 20534 34776
rect 20590 34720 20595 34776
rect 19149 34718 20595 34720
rect 19149 34715 19215 34718
rect 20529 34715 20595 34718
rect 21173 34778 21239 34781
rect 24945 34780 25011 34781
rect 21582 34778 21588 34780
rect 21173 34776 21588 34778
rect 21173 34720 21178 34776
rect 21234 34720 21588 34776
rect 21173 34718 21588 34720
rect 21173 34715 21239 34718
rect 21582 34716 21588 34718
rect 21652 34716 21658 34780
rect 24894 34716 24900 34780
rect 24964 34778 25011 34780
rect 24964 34776 25056 34778
rect 25006 34720 25056 34776
rect 24964 34718 25056 34720
rect 24964 34716 25011 34718
rect 24945 34715 25011 34716
rect 3141 34642 3207 34645
rect 18137 34642 18203 34645
rect 31661 34642 31727 34645
rect 3141 34640 31727 34642
rect 3141 34584 3146 34640
rect 3202 34584 18142 34640
rect 18198 34584 31666 34640
rect 31722 34584 31727 34640
rect 3141 34582 31727 34584
rect 3141 34579 3207 34582
rect 18137 34579 18203 34582
rect 31661 34579 31727 34582
rect 35433 34642 35499 34645
rect 39389 34642 39455 34645
rect 35433 34640 39455 34642
rect 35433 34584 35438 34640
rect 35494 34584 39394 34640
rect 39450 34584 39455 34640
rect 35433 34582 39455 34584
rect 35433 34579 35499 34582
rect 39389 34579 39455 34582
rect 35801 34506 35867 34509
rect 39520 34506 40000 34536
rect 35801 34504 40000 34506
rect 35801 34448 35806 34504
rect 35862 34448 40000 34504
rect 35801 34446 40000 34448
rect 35801 34443 35867 34446
rect 39520 34416 40000 34446
rect 9581 34370 9647 34373
rect 11237 34370 11303 34373
rect 9581 34368 11303 34370
rect 9581 34312 9586 34368
rect 9642 34312 11242 34368
rect 11298 34312 11303 34368
rect 9581 34310 11303 34312
rect 9581 34307 9647 34310
rect 11237 34307 11303 34310
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 20069 34234 20135 34237
rect 23565 34234 23631 34237
rect 20069 34232 23631 34234
rect 20069 34176 20074 34232
rect 20130 34176 23570 34232
rect 23626 34176 23631 34232
rect 20069 34174 23631 34176
rect 20069 34171 20135 34174
rect 23565 34171 23631 34174
rect 2865 34098 2931 34101
rect 11605 34098 11671 34101
rect 2865 34096 11671 34098
rect 2865 34040 2870 34096
rect 2926 34040 11610 34096
rect 11666 34040 11671 34096
rect 2865 34038 11671 34040
rect 2865 34035 2931 34038
rect 11605 34035 11671 34038
rect 12617 33962 12683 33965
rect 17902 33962 17908 33964
rect 12617 33960 17908 33962
rect 12617 33904 12622 33960
rect 12678 33904 17908 33960
rect 12617 33902 17908 33904
rect 12617 33899 12683 33902
rect 17902 33900 17908 33902
rect 17972 33900 17978 33964
rect 27521 33962 27587 33965
rect 30557 33962 30623 33965
rect 27521 33960 30623 33962
rect 27521 33904 27526 33960
rect 27582 33904 30562 33960
rect 30618 33904 30623 33960
rect 27521 33902 30623 33904
rect 27521 33899 27587 33902
rect 30557 33899 30623 33902
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 17902 33628 17908 33692
rect 17972 33690 17978 33692
rect 27521 33690 27587 33693
rect 17972 33688 27587 33690
rect 17972 33632 27526 33688
rect 27582 33632 27587 33688
rect 17972 33630 27587 33632
rect 17972 33628 17978 33630
rect 27521 33627 27587 33630
rect 10777 33554 10843 33557
rect 12801 33554 12867 33557
rect 15653 33554 15719 33557
rect 10777 33552 15719 33554
rect 10777 33496 10782 33552
rect 10838 33496 12806 33552
rect 12862 33496 15658 33552
rect 15714 33496 15719 33552
rect 10777 33494 15719 33496
rect 10777 33491 10843 33494
rect 12801 33491 12867 33494
rect 15653 33491 15719 33494
rect 15929 33554 15995 33557
rect 30189 33554 30255 33557
rect 35709 33554 35775 33557
rect 15929 33552 35775 33554
rect 15929 33496 15934 33552
rect 15990 33496 30194 33552
rect 30250 33496 35714 33552
rect 35770 33496 35775 33552
rect 15929 33494 35775 33496
rect 15929 33491 15995 33494
rect 30189 33491 30255 33494
rect 35709 33491 35775 33494
rect 0 33328 480 33448
rect 12893 33282 12959 33285
rect 16021 33282 16087 33285
rect 17033 33282 17099 33285
rect 12893 33280 17099 33282
rect 12893 33224 12898 33280
rect 12954 33224 16026 33280
rect 16082 33224 17038 33280
rect 17094 33224 17099 33280
rect 12893 33222 17099 33224
rect 12893 33219 12959 33222
rect 16021 33219 16087 33222
rect 17033 33219 17099 33222
rect 35617 33282 35683 33285
rect 39520 33282 40000 33312
rect 35617 33280 40000 33282
rect 35617 33224 35622 33280
rect 35678 33224 40000 33280
rect 35617 33222 40000 33224
rect 35617 33219 35683 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 39520 33192 40000 33222
rect 19568 33151 19888 33152
rect 24853 33010 24919 33013
rect 29361 33010 29427 33013
rect 24853 33008 29427 33010
rect 24853 32952 24858 33008
rect 24914 32952 29366 33008
rect 29422 32952 29427 33008
rect 24853 32950 29427 32952
rect 24853 32947 24919 32950
rect 29361 32947 29427 32950
rect 14089 32874 14155 32877
rect 16757 32874 16823 32877
rect 14089 32872 16823 32874
rect 14089 32816 14094 32872
rect 14150 32816 16762 32872
rect 16818 32816 16823 32872
rect 14089 32814 16823 32816
rect 14089 32811 14155 32814
rect 16757 32811 16823 32814
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 9857 32602 9923 32605
rect 13261 32602 13327 32605
rect 9857 32600 13327 32602
rect 9857 32544 9862 32600
rect 9918 32544 13266 32600
rect 13322 32544 13327 32600
rect 9857 32542 13327 32544
rect 9857 32539 9923 32542
rect 13261 32539 13327 32542
rect 17585 32602 17651 32605
rect 20161 32602 20227 32605
rect 17585 32600 20227 32602
rect 17585 32544 17590 32600
rect 17646 32544 20166 32600
rect 20222 32544 20227 32600
rect 17585 32542 20227 32544
rect 17585 32539 17651 32542
rect 20161 32539 20227 32542
rect 14917 32466 14983 32469
rect 16665 32466 16731 32469
rect 14917 32464 16731 32466
rect 14917 32408 14922 32464
rect 14978 32408 16670 32464
rect 16726 32408 16731 32464
rect 14917 32406 16731 32408
rect 14917 32403 14983 32406
rect 16665 32403 16731 32406
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 35709 32058 35775 32061
rect 39520 32058 40000 32088
rect 35709 32056 40000 32058
rect 35709 32000 35714 32056
rect 35770 32000 40000 32056
rect 35709 31998 40000 32000
rect 35709 31995 35775 31998
rect 39520 31968 40000 31998
rect 4061 31922 4127 31925
rect 5625 31922 5691 31925
rect 4061 31920 5691 31922
rect 4061 31864 4066 31920
rect 4122 31864 5630 31920
rect 5686 31864 5691 31920
rect 4061 31862 5691 31864
rect 4061 31859 4127 31862
rect 5625 31859 5691 31862
rect 25221 31922 25287 31925
rect 29545 31922 29611 31925
rect 25221 31920 29611 31922
rect 25221 31864 25226 31920
rect 25282 31864 29550 31920
rect 29606 31864 29611 31920
rect 25221 31862 29611 31864
rect 25221 31859 25287 31862
rect 29545 31859 29611 31862
rect 16481 31650 16547 31653
rect 19425 31650 19491 31653
rect 16481 31648 19491 31650
rect 16481 31592 16486 31648
rect 16542 31592 19430 31648
rect 19486 31592 19491 31648
rect 16481 31590 19491 31592
rect 16481 31587 16547 31590
rect 19425 31587 19491 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 11881 31514 11947 31517
rect 14825 31514 14891 31517
rect 11881 31512 14891 31514
rect 11881 31456 11886 31512
rect 11942 31456 14830 31512
rect 14886 31456 14891 31512
rect 11881 31454 14891 31456
rect 11881 31451 11947 31454
rect 14825 31451 14891 31454
rect 17033 31514 17099 31517
rect 18873 31514 18939 31517
rect 17033 31512 18939 31514
rect 17033 31456 17038 31512
rect 17094 31456 18878 31512
rect 18934 31456 18939 31512
rect 17033 31454 18939 31456
rect 17033 31451 17099 31454
rect 18873 31451 18939 31454
rect 24761 31242 24827 31245
rect 28165 31242 28231 31245
rect 24761 31240 28231 31242
rect 24761 31184 24766 31240
rect 24822 31184 28170 31240
rect 28226 31184 28231 31240
rect 24761 31182 28231 31184
rect 24761 31179 24827 31182
rect 28165 31179 28231 31182
rect 12709 31106 12775 31109
rect 15469 31106 15535 31109
rect 12709 31104 15535 31106
rect 12709 31048 12714 31104
rect 12770 31048 15474 31104
rect 15530 31048 15535 31104
rect 12709 31046 15535 31048
rect 12709 31043 12775 31046
rect 15469 31043 15535 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 11145 30970 11211 30973
rect 14365 30970 14431 30973
rect 11145 30968 14431 30970
rect 11145 30912 11150 30968
rect 11206 30912 14370 30968
rect 14426 30912 14431 30968
rect 11145 30910 14431 30912
rect 11145 30907 11211 30910
rect 14365 30907 14431 30910
rect 20621 30834 20687 30837
rect 22553 30834 22619 30837
rect 20621 30832 22619 30834
rect 20621 30776 20626 30832
rect 20682 30776 22558 30832
rect 22614 30776 22619 30832
rect 20621 30774 22619 30776
rect 20621 30771 20687 30774
rect 22553 30771 22619 30774
rect 35893 30834 35959 30837
rect 39520 30834 40000 30864
rect 35893 30832 40000 30834
rect 35893 30776 35898 30832
rect 35954 30776 40000 30832
rect 35893 30774 40000 30776
rect 35893 30771 35959 30774
rect 39520 30744 40000 30774
rect 1669 30698 1735 30701
rect 5901 30698 5967 30701
rect 7005 30698 7071 30701
rect 1669 30696 7071 30698
rect 1669 30640 1674 30696
rect 1730 30640 5906 30696
rect 5962 30640 7010 30696
rect 7066 30640 7071 30696
rect 1669 30638 7071 30640
rect 1669 30635 1735 30638
rect 5901 30635 5967 30638
rect 7005 30635 7071 30638
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 10777 30426 10843 30429
rect 12709 30426 12775 30429
rect 10777 30424 12775 30426
rect 10777 30368 10782 30424
rect 10838 30368 12714 30424
rect 12770 30368 12775 30424
rect 10777 30366 12775 30368
rect 10777 30363 10843 30366
rect 12709 30363 12775 30366
rect 13721 30426 13787 30429
rect 16941 30426 17007 30429
rect 13721 30424 17007 30426
rect 13721 30368 13726 30424
rect 13782 30368 16946 30424
rect 17002 30368 17007 30424
rect 13721 30366 17007 30368
rect 13721 30363 13787 30366
rect 16941 30363 17007 30366
rect 24393 30290 24459 30293
rect 26969 30290 27035 30293
rect 24393 30288 27035 30290
rect 24393 30232 24398 30288
rect 24454 30232 26974 30288
rect 27030 30232 27035 30288
rect 24393 30230 27035 30232
rect 24393 30227 24459 30230
rect 26969 30227 27035 30230
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 15837 29610 15903 29613
rect 18873 29610 18939 29613
rect 15837 29608 18939 29610
rect 15837 29552 15842 29608
rect 15898 29552 18878 29608
rect 18934 29552 18939 29608
rect 15837 29550 18939 29552
rect 15837 29547 15903 29550
rect 18873 29547 18939 29550
rect 35525 29610 35591 29613
rect 39520 29610 40000 29640
rect 35525 29608 40000 29610
rect 35525 29552 35530 29608
rect 35586 29552 40000 29608
rect 35525 29550 40000 29552
rect 35525 29547 35591 29550
rect 39520 29520 40000 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 24761 29338 24827 29341
rect 26417 29338 26483 29341
rect 24761 29336 26483 29338
rect 24761 29280 24766 29336
rect 24822 29280 26422 29336
rect 26478 29280 26483 29336
rect 24761 29278 26483 29280
rect 24761 29275 24827 29278
rect 26417 29275 26483 29278
rect 21817 28930 21883 28933
rect 23657 28930 23723 28933
rect 21817 28928 23723 28930
rect 21817 28872 21822 28928
rect 21878 28872 23662 28928
rect 23718 28872 23723 28928
rect 21817 28870 23723 28872
rect 21817 28867 21883 28870
rect 23657 28867 23723 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 39520 28386 40000 28416
rect 35574 28326 40000 28386
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 25865 28114 25931 28117
rect 27889 28114 27955 28117
rect 25865 28112 27955 28114
rect 25865 28056 25870 28112
rect 25926 28056 27894 28112
rect 27950 28056 27955 28112
rect 25865 28054 27955 28056
rect 25865 28051 25931 28054
rect 27889 28051 27955 28054
rect 34513 28114 34579 28117
rect 35574 28114 35634 28326
rect 39520 28296 40000 28326
rect 34513 28112 35634 28114
rect 34513 28056 34518 28112
rect 34574 28056 35634 28112
rect 34513 28054 35634 28056
rect 34513 28051 34579 28054
rect 8201 27842 8267 27845
rect 10225 27842 10291 27845
rect 8201 27840 10291 27842
rect 8201 27784 8206 27840
rect 8262 27784 10230 27840
rect 10286 27784 10291 27840
rect 8201 27782 10291 27784
rect 8201 27779 8267 27782
rect 10225 27779 10291 27782
rect 33777 27842 33843 27845
rect 35893 27842 35959 27845
rect 33777 27840 35959 27842
rect 33777 27784 33782 27840
rect 33838 27784 35898 27840
rect 35954 27784 35959 27840
rect 33777 27782 35959 27784
rect 33777 27779 33843 27782
rect 35893 27779 35959 27782
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 10133 27570 10199 27573
rect 12709 27570 12775 27573
rect 10133 27568 12775 27570
rect 10133 27512 10138 27568
rect 10194 27512 12714 27568
rect 12770 27512 12775 27568
rect 10133 27510 12775 27512
rect 10133 27507 10199 27510
rect 12709 27507 12775 27510
rect 17033 27570 17099 27573
rect 19885 27570 19951 27573
rect 17033 27568 19951 27570
rect 17033 27512 17038 27568
rect 17094 27512 19890 27568
rect 19946 27512 19951 27568
rect 17033 27510 19951 27512
rect 17033 27507 17099 27510
rect 19885 27507 19951 27510
rect 31661 27298 31727 27301
rect 33225 27298 33291 27301
rect 31661 27296 33291 27298
rect 31661 27240 31666 27296
rect 31722 27240 33230 27296
rect 33286 27240 33291 27296
rect 31661 27238 33291 27240
rect 31661 27235 31727 27238
rect 33225 27235 33291 27238
rect 37181 27298 37247 27301
rect 39520 27298 40000 27328
rect 37181 27296 40000 27298
rect 37181 27240 37186 27296
rect 37242 27240 40000 27296
rect 37181 27238 40000 27240
rect 37181 27235 37247 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 39520 27208 40000 27238
rect 34928 27167 35248 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 14733 26482 14799 26485
rect 20161 26482 20227 26485
rect 14733 26480 20227 26482
rect 14733 26424 14738 26480
rect 14794 26424 20166 26480
rect 20222 26424 20227 26480
rect 14733 26422 20227 26424
rect 14733 26419 14799 26422
rect 20161 26419 20227 26422
rect 31569 26482 31635 26485
rect 33225 26482 33291 26485
rect 31569 26480 33291 26482
rect 31569 26424 31574 26480
rect 31630 26424 33230 26480
rect 33286 26424 33291 26480
rect 31569 26422 33291 26424
rect 31569 26419 31635 26422
rect 33225 26419 33291 26422
rect 10409 26346 10475 26349
rect 12525 26346 12591 26349
rect 10409 26344 12591 26346
rect 10409 26288 10414 26344
rect 10470 26288 12530 26344
rect 12586 26288 12591 26344
rect 10409 26286 12591 26288
rect 10409 26283 10475 26286
rect 12525 26283 12591 26286
rect 23841 26346 23907 26349
rect 25589 26346 25655 26349
rect 26233 26346 26299 26349
rect 23841 26344 26299 26346
rect 23841 26288 23846 26344
rect 23902 26288 25594 26344
rect 25650 26288 26238 26344
rect 26294 26288 26299 26344
rect 23841 26286 26299 26288
rect 23841 26283 23907 26286
rect 25589 26283 25655 26286
rect 26233 26283 26299 26286
rect 28441 26346 28507 26349
rect 31293 26346 31359 26349
rect 28441 26344 31359 26346
rect 28441 26288 28446 26344
rect 28502 26288 31298 26344
rect 31354 26288 31359 26344
rect 28441 26286 31359 26288
rect 28441 26283 28507 26286
rect 31293 26283 31359 26286
rect 24209 26210 24275 26213
rect 26969 26210 27035 26213
rect 24209 26208 27035 26210
rect 24209 26152 24214 26208
rect 24270 26152 26974 26208
rect 27030 26152 27035 26208
rect 24209 26150 27035 26152
rect 24209 26147 24275 26150
rect 26969 26147 27035 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 36445 26074 36511 26077
rect 39520 26074 40000 26104
rect 36445 26072 40000 26074
rect 36445 26016 36450 26072
rect 36506 26016 40000 26072
rect 36445 26014 40000 26016
rect 36445 26011 36511 26014
rect 39520 25984 40000 26014
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 20621 25530 20687 25533
rect 22001 25530 22067 25533
rect 23657 25530 23723 25533
rect 26233 25530 26299 25533
rect 20621 25528 26299 25530
rect 20621 25472 20626 25528
rect 20682 25472 22006 25528
rect 22062 25472 23662 25528
rect 23718 25472 26238 25528
rect 26294 25472 26299 25528
rect 20621 25470 26299 25472
rect 20621 25467 20687 25470
rect 22001 25467 22067 25470
rect 23657 25467 23723 25470
rect 26233 25467 26299 25470
rect 34053 25394 34119 25397
rect 36813 25394 36879 25397
rect 34053 25392 36879 25394
rect 34053 25336 34058 25392
rect 34114 25336 36818 25392
rect 36874 25336 36879 25392
rect 34053 25334 36879 25336
rect 34053 25331 34119 25334
rect 36813 25331 36879 25334
rect 26601 25122 26667 25125
rect 28717 25122 28783 25125
rect 26601 25120 28783 25122
rect 26601 25064 26606 25120
rect 26662 25064 28722 25120
rect 28778 25064 28783 25120
rect 26601 25062 28783 25064
rect 26601 25059 26667 25062
rect 28717 25059 28783 25062
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 18597 24986 18663 24989
rect 20713 24986 20779 24989
rect 18597 24984 20779 24986
rect 18597 24928 18602 24984
rect 18658 24928 20718 24984
rect 20774 24928 20779 24984
rect 18597 24926 20779 24928
rect 18597 24923 18663 24926
rect 20713 24923 20779 24926
rect 27797 24986 27863 24989
rect 32029 24986 32095 24989
rect 27797 24984 32095 24986
rect 27797 24928 27802 24984
rect 27858 24928 32034 24984
rect 32090 24928 32095 24984
rect 27797 24926 32095 24928
rect 27797 24923 27863 24926
rect 32029 24923 32095 24926
rect 8477 24850 8543 24853
rect 9213 24850 9279 24853
rect 11881 24850 11947 24853
rect 12893 24850 12959 24853
rect 8477 24848 12959 24850
rect 8477 24792 8482 24848
rect 8538 24792 9218 24848
rect 9274 24792 11886 24848
rect 11942 24792 12898 24848
rect 12954 24792 12959 24848
rect 8477 24790 12959 24792
rect 8477 24787 8543 24790
rect 9213 24787 9279 24790
rect 11881 24787 11947 24790
rect 12893 24787 12959 24790
rect 18689 24850 18755 24853
rect 20897 24850 20963 24853
rect 18689 24848 20963 24850
rect 18689 24792 18694 24848
rect 18750 24792 20902 24848
rect 20958 24792 20963 24848
rect 18689 24790 20963 24792
rect 18689 24787 18755 24790
rect 20897 24787 20963 24790
rect 25037 24850 25103 24853
rect 39520 24850 40000 24880
rect 25037 24848 40000 24850
rect 25037 24792 25042 24848
rect 25098 24792 40000 24848
rect 25037 24790 40000 24792
rect 25037 24787 25103 24790
rect 39520 24760 40000 24790
rect 7649 24578 7715 24581
rect 11513 24578 11579 24581
rect 7649 24576 11579 24578
rect 7649 24520 7654 24576
rect 7710 24520 11518 24576
rect 11574 24520 11579 24576
rect 7649 24518 11579 24520
rect 7649 24515 7715 24518
rect 11513 24515 11579 24518
rect 16389 24578 16455 24581
rect 18689 24578 18755 24581
rect 16389 24576 18755 24578
rect 16389 24520 16394 24576
rect 16450 24520 18694 24576
rect 18750 24520 18755 24576
rect 16389 24518 18755 24520
rect 16389 24515 16455 24518
rect 18689 24515 18755 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 19977 24306 20043 24309
rect 21357 24306 21423 24309
rect 19977 24304 21423 24306
rect 19977 24248 19982 24304
rect 20038 24248 21362 24304
rect 21418 24248 21423 24304
rect 19977 24246 21423 24248
rect 19977 24243 20043 24246
rect 21357 24243 21423 24246
rect 28901 24034 28967 24037
rect 31937 24034 32003 24037
rect 28901 24032 32003 24034
rect 28901 23976 28906 24032
rect 28962 23976 31942 24032
rect 31998 23976 32003 24032
rect 28901 23974 32003 23976
rect 28901 23971 28967 23974
rect 31937 23971 32003 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 34513 23762 34579 23765
rect 34646 23762 34652 23764
rect 34513 23760 34652 23762
rect 34513 23704 34518 23760
rect 34574 23704 34652 23760
rect 34513 23702 34652 23704
rect 34513 23699 34579 23702
rect 34646 23700 34652 23702
rect 34716 23700 34722 23764
rect 15285 23626 15351 23629
rect 18045 23626 18111 23629
rect 15285 23624 18111 23626
rect 15285 23568 15290 23624
rect 15346 23568 18050 23624
rect 18106 23568 18111 23624
rect 15285 23566 18111 23568
rect 15285 23563 15351 23566
rect 18045 23563 18111 23566
rect 35249 23626 35315 23629
rect 39520 23626 40000 23656
rect 35249 23624 40000 23626
rect 35249 23568 35254 23624
rect 35310 23568 40000 23624
rect 35249 23566 40000 23568
rect 35249 23563 35315 23566
rect 39520 23536 40000 23566
rect 12709 23490 12775 23493
rect 16481 23490 16547 23493
rect 12709 23488 16547 23490
rect 12709 23432 12714 23488
rect 12770 23432 16486 23488
rect 16542 23432 16547 23488
rect 12709 23430 16547 23432
rect 12709 23427 12775 23430
rect 16481 23427 16547 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 12985 22946 13051 22949
rect 16389 22946 16455 22949
rect 12985 22944 16455 22946
rect 12985 22888 12990 22944
rect 13046 22888 16394 22944
rect 16450 22888 16455 22944
rect 12985 22886 16455 22888
rect 12985 22883 13051 22886
rect 16389 22883 16455 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 21541 22810 21607 22813
rect 25681 22810 25747 22813
rect 21541 22808 25747 22810
rect 21541 22752 21546 22808
rect 21602 22752 25686 22808
rect 25742 22752 25747 22808
rect 21541 22750 25747 22752
rect 21541 22747 21607 22750
rect 25681 22747 25747 22750
rect 24485 22538 24551 22541
rect 26877 22538 26943 22541
rect 24485 22536 26943 22538
rect 24485 22480 24490 22536
rect 24546 22480 26882 22536
rect 26938 22480 26943 22536
rect 24485 22478 26943 22480
rect 24485 22475 24551 22478
rect 26877 22475 26943 22478
rect 36077 22402 36143 22405
rect 39520 22402 40000 22432
rect 36077 22400 40000 22402
rect 36077 22344 36082 22400
rect 36138 22344 40000 22400
rect 36077 22342 40000 22344
rect 36077 22339 36143 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 39520 22312 40000 22342
rect 19568 22271 19888 22272
rect 12801 21994 12867 21997
rect 13997 21994 14063 21997
rect 12801 21992 14063 21994
rect 12801 21936 12806 21992
rect 12862 21936 14002 21992
rect 14058 21936 14063 21992
rect 12801 21934 14063 21936
rect 12801 21931 12867 21934
rect 13997 21931 14063 21934
rect 28441 21994 28507 21997
rect 35249 21994 35315 21997
rect 28441 21992 35315 21994
rect 28441 21936 28446 21992
rect 28502 21936 35254 21992
rect 35310 21936 35315 21992
rect 28441 21934 35315 21936
rect 28441 21931 28507 21934
rect 35249 21931 35315 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 24669 21586 24735 21589
rect 26693 21586 26759 21589
rect 24669 21584 26759 21586
rect 24669 21528 24674 21584
rect 24730 21528 26698 21584
rect 26754 21528 26759 21584
rect 24669 21526 26759 21528
rect 24669 21523 24735 21526
rect 26693 21523 26759 21526
rect 35249 21586 35315 21589
rect 35433 21586 35499 21589
rect 35249 21584 35499 21586
rect 35249 21528 35254 21584
rect 35310 21528 35438 21584
rect 35494 21528 35499 21584
rect 35249 21526 35499 21528
rect 35249 21523 35315 21526
rect 35433 21523 35499 21526
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 35709 21178 35775 21181
rect 39520 21178 40000 21208
rect 35709 21176 40000 21178
rect 35709 21120 35714 21176
rect 35770 21120 40000 21176
rect 35709 21118 40000 21120
rect 35709 21115 35775 21118
rect 39520 21088 40000 21118
rect 33225 20906 33291 20909
rect 36169 20906 36235 20909
rect 33225 20904 36235 20906
rect 33225 20848 33230 20904
rect 33286 20848 36174 20904
rect 36230 20848 36235 20904
rect 33225 20846 36235 20848
rect 33225 20843 33291 20846
rect 36169 20843 36235 20846
rect 20161 20770 20227 20773
rect 27705 20770 27771 20773
rect 20161 20768 27771 20770
rect 20161 20712 20166 20768
rect 20222 20712 27710 20768
rect 27766 20712 27771 20768
rect 20161 20710 27771 20712
rect 20161 20707 20227 20710
rect 27705 20707 27771 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 27613 20634 27679 20637
rect 34646 20634 34652 20636
rect 27613 20632 34652 20634
rect 27613 20576 27618 20632
rect 27674 20576 34652 20632
rect 27613 20574 34652 20576
rect 27613 20571 27679 20574
rect 34646 20572 34652 20574
rect 34716 20572 34722 20636
rect 24301 20498 24367 20501
rect 27981 20498 28047 20501
rect 24301 20496 28047 20498
rect 24301 20440 24306 20496
rect 24362 20440 27986 20496
rect 28042 20440 28047 20496
rect 24301 20438 28047 20440
rect 24301 20435 24367 20438
rect 27981 20435 28047 20438
rect 19517 20362 19583 20365
rect 22185 20362 22251 20365
rect 19517 20360 22251 20362
rect 19517 20304 19522 20360
rect 19578 20304 22190 20360
rect 22246 20304 22251 20360
rect 19517 20302 22251 20304
rect 19517 20299 19583 20302
rect 22185 20299 22251 20302
rect 26049 20226 26115 20229
rect 29453 20226 29519 20229
rect 26049 20224 29519 20226
rect 26049 20168 26054 20224
rect 26110 20168 29458 20224
rect 29514 20168 29519 20224
rect 26049 20166 29519 20168
rect 26049 20163 26115 20166
rect 29453 20163 29519 20166
rect 30097 20226 30163 20229
rect 31017 20226 31083 20229
rect 33317 20226 33383 20229
rect 30097 20224 33383 20226
rect 30097 20168 30102 20224
rect 30158 20168 31022 20224
rect 31078 20168 33322 20224
rect 33378 20168 33383 20224
rect 30097 20166 33383 20168
rect 30097 20163 30163 20166
rect 31017 20163 31083 20166
rect 33317 20163 33383 20166
rect 19568 20160 19888 20161
rect 0 20090 480 20120
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 2773 20090 2839 20093
rect 0 20088 2839 20090
rect 0 20032 2778 20088
rect 2834 20032 2839 20088
rect 0 20030 2839 20032
rect 0 20000 480 20030
rect 2773 20027 2839 20030
rect 21357 20090 21423 20093
rect 23657 20090 23723 20093
rect 21357 20088 23723 20090
rect 21357 20032 21362 20088
rect 21418 20032 23662 20088
rect 23718 20032 23723 20088
rect 21357 20030 23723 20032
rect 21357 20027 21423 20030
rect 23657 20027 23723 20030
rect 28993 20090 29059 20093
rect 31753 20090 31819 20093
rect 28993 20088 31819 20090
rect 28993 20032 28998 20088
rect 29054 20032 31758 20088
rect 31814 20032 31819 20088
rect 28993 20030 31819 20032
rect 28993 20027 29059 20030
rect 31753 20027 31819 20030
rect 26509 19954 26575 19957
rect 35709 19954 35775 19957
rect 39520 19954 40000 19984
rect 26509 19952 35775 19954
rect 26509 19896 26514 19952
rect 26570 19896 35714 19952
rect 35770 19896 35775 19952
rect 26509 19894 35775 19896
rect 26509 19891 26575 19894
rect 35709 19891 35775 19894
rect 35942 19894 40000 19954
rect 35341 19818 35407 19821
rect 35942 19818 36002 19894
rect 39520 19864 40000 19894
rect 35341 19816 36002 19818
rect 35341 19760 35346 19816
rect 35402 19760 36002 19816
rect 35341 19758 36002 19760
rect 35341 19755 35407 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 29361 19546 29427 19549
rect 34237 19546 34303 19549
rect 29361 19544 34303 19546
rect 29361 19488 29366 19544
rect 29422 19488 34242 19544
rect 34298 19488 34303 19544
rect 29361 19486 34303 19488
rect 29361 19483 29427 19486
rect 34237 19483 34303 19486
rect 24209 19410 24275 19413
rect 24485 19410 24551 19413
rect 24209 19408 24551 19410
rect 24209 19352 24214 19408
rect 24270 19352 24490 19408
rect 24546 19352 24551 19408
rect 24209 19350 24551 19352
rect 24209 19347 24275 19350
rect 24485 19347 24551 19350
rect 23749 19274 23815 19277
rect 26877 19274 26943 19277
rect 23749 19272 26943 19274
rect 23749 19216 23754 19272
rect 23810 19216 26882 19272
rect 26938 19216 26943 19272
rect 23749 19214 26943 19216
rect 23749 19211 23815 19214
rect 26877 19211 26943 19214
rect 33777 19274 33843 19277
rect 35985 19274 36051 19277
rect 33777 19272 36051 19274
rect 33777 19216 33782 19272
rect 33838 19216 35990 19272
rect 36046 19216 36051 19272
rect 33777 19214 36051 19216
rect 33777 19211 33843 19214
rect 35985 19211 36051 19214
rect 25773 19138 25839 19141
rect 34789 19138 34855 19141
rect 25773 19136 34855 19138
rect 25773 19080 25778 19136
rect 25834 19080 34794 19136
rect 34850 19080 34855 19136
rect 25773 19078 34855 19080
rect 25773 19075 25839 19078
rect 34789 19075 34855 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 24025 19002 24091 19005
rect 26693 19002 26759 19005
rect 24025 19000 26759 19002
rect 24025 18944 24030 19000
rect 24086 18944 26698 19000
rect 26754 18944 26759 19000
rect 24025 18942 26759 18944
rect 24025 18939 24091 18942
rect 26693 18939 26759 18942
rect 27061 19002 27127 19005
rect 29913 19002 29979 19005
rect 27061 19000 29979 19002
rect 27061 18944 27066 19000
rect 27122 18944 29918 19000
rect 29974 18944 29979 19000
rect 27061 18942 29979 18944
rect 27061 18939 27127 18942
rect 29913 18939 29979 18942
rect 36537 18730 36603 18733
rect 39520 18730 40000 18760
rect 36537 18728 40000 18730
rect 36537 18672 36542 18728
rect 36598 18672 40000 18728
rect 36537 18670 40000 18672
rect 36537 18667 36603 18670
rect 39520 18640 40000 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 19241 18322 19307 18325
rect 22369 18322 22435 18325
rect 19241 18320 22435 18322
rect 19241 18264 19246 18320
rect 19302 18264 22374 18320
rect 22430 18264 22435 18320
rect 19241 18262 22435 18264
rect 19241 18259 19307 18262
rect 22369 18259 22435 18262
rect 20069 18186 20135 18189
rect 21081 18186 21147 18189
rect 23841 18186 23907 18189
rect 20069 18184 23907 18186
rect 20069 18128 20074 18184
rect 20130 18128 21086 18184
rect 21142 18128 23846 18184
rect 23902 18128 23907 18184
rect 20069 18126 23907 18128
rect 20069 18123 20135 18126
rect 21081 18123 21147 18126
rect 23841 18123 23907 18126
rect 20345 18050 20411 18053
rect 22277 18050 22343 18053
rect 20345 18048 22343 18050
rect 20345 17992 20350 18048
rect 20406 17992 22282 18048
rect 22338 17992 22343 18048
rect 20345 17990 22343 17992
rect 20345 17987 20411 17990
rect 22277 17987 22343 17990
rect 32673 18050 32739 18053
rect 34697 18050 34763 18053
rect 32673 18048 34763 18050
rect 32673 17992 32678 18048
rect 32734 17992 34702 18048
rect 34758 17992 34763 18048
rect 32673 17990 34763 17992
rect 32673 17987 32739 17990
rect 34697 17987 34763 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 25221 17914 25287 17917
rect 27889 17914 27955 17917
rect 25221 17912 27955 17914
rect 25221 17856 25226 17912
rect 25282 17856 27894 17912
rect 27950 17856 27955 17912
rect 25221 17854 27955 17856
rect 25221 17851 25287 17854
rect 27889 17851 27955 17854
rect 28717 17642 28783 17645
rect 35341 17642 35407 17645
rect 28717 17640 35407 17642
rect 28717 17584 28722 17640
rect 28778 17584 35346 17640
rect 35402 17584 35407 17640
rect 28717 17582 35407 17584
rect 28717 17579 28783 17582
rect 35341 17579 35407 17582
rect 39520 17506 40000 17536
rect 35390 17446 40000 17506
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 21541 17370 21607 17373
rect 25221 17370 25287 17373
rect 21541 17368 25287 17370
rect 21541 17312 21546 17368
rect 21602 17312 25226 17368
rect 25282 17312 25287 17368
rect 21541 17310 25287 17312
rect 21541 17307 21607 17310
rect 25221 17307 25287 17310
rect 19241 17234 19307 17237
rect 22277 17234 22343 17237
rect 19241 17232 22343 17234
rect 19241 17176 19246 17232
rect 19302 17176 22282 17232
rect 22338 17176 22343 17232
rect 19241 17174 22343 17176
rect 19241 17171 19307 17174
rect 22277 17171 22343 17174
rect 34605 17234 34671 17237
rect 35390 17234 35450 17446
rect 39520 17416 40000 17446
rect 34605 17232 35450 17234
rect 34605 17176 34610 17232
rect 34666 17176 35450 17232
rect 34605 17174 35450 17176
rect 34605 17171 34671 17174
rect 19241 17098 19307 17101
rect 21725 17098 21791 17101
rect 19241 17096 21791 17098
rect 19241 17040 19246 17096
rect 19302 17040 21730 17096
rect 21786 17040 21791 17096
rect 19241 17038 21791 17040
rect 19241 17035 19307 17038
rect 21725 17035 21791 17038
rect 25497 17098 25563 17101
rect 31385 17098 31451 17101
rect 25497 17096 31451 17098
rect 25497 17040 25502 17096
rect 25558 17040 31390 17096
rect 31446 17040 31451 17096
rect 25497 17038 31451 17040
rect 25497 17035 25563 17038
rect 31385 17035 31451 17038
rect 27429 16962 27495 16965
rect 28993 16962 29059 16965
rect 27429 16960 29059 16962
rect 27429 16904 27434 16960
rect 27490 16904 28998 16960
rect 29054 16904 29059 16960
rect 27429 16902 29059 16904
rect 27429 16899 27495 16902
rect 28993 16899 29059 16902
rect 35433 16962 35499 16965
rect 35566 16962 35572 16964
rect 35433 16960 35572 16962
rect 35433 16904 35438 16960
rect 35494 16904 35572 16960
rect 35433 16902 35572 16904
rect 35433 16899 35499 16902
rect 35566 16900 35572 16902
rect 35636 16900 35642 16964
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 20253 16690 20319 16693
rect 22277 16690 22343 16693
rect 20253 16688 22343 16690
rect 20253 16632 20258 16688
rect 20314 16632 22282 16688
rect 22338 16632 22343 16688
rect 20253 16630 22343 16632
rect 20253 16627 20319 16630
rect 22277 16627 22343 16630
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 35525 16282 35591 16285
rect 39520 16282 40000 16312
rect 35525 16280 40000 16282
rect 35525 16224 35530 16280
rect 35586 16224 40000 16280
rect 35525 16222 40000 16224
rect 35525 16219 35591 16222
rect 39520 16192 40000 16222
rect 27705 15874 27771 15877
rect 36077 15874 36143 15877
rect 27705 15872 36143 15874
rect 27705 15816 27710 15872
rect 27766 15816 36082 15872
rect 36138 15816 36143 15872
rect 27705 15814 36143 15816
rect 27705 15811 27771 15814
rect 36077 15811 36143 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 28625 15738 28691 15741
rect 30557 15738 30623 15741
rect 28625 15736 30623 15738
rect 28625 15680 28630 15736
rect 28686 15680 30562 15736
rect 30618 15680 30623 15736
rect 28625 15678 30623 15680
rect 28625 15675 28691 15678
rect 30557 15675 30623 15678
rect 31845 15466 31911 15469
rect 32949 15466 33015 15469
rect 36813 15466 36879 15469
rect 31845 15464 36879 15466
rect 31845 15408 31850 15464
rect 31906 15408 32954 15464
rect 33010 15408 36818 15464
rect 36874 15408 36879 15464
rect 31845 15406 36879 15408
rect 31845 15403 31911 15406
rect 32949 15403 33015 15406
rect 36813 15403 36879 15406
rect 30281 15330 30347 15333
rect 32765 15330 32831 15333
rect 30281 15328 32831 15330
rect 30281 15272 30286 15328
rect 30342 15272 32770 15328
rect 32826 15272 32831 15328
rect 30281 15270 32831 15272
rect 30281 15267 30347 15270
rect 32765 15267 32831 15270
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 28441 15194 28507 15197
rect 34605 15194 34671 15197
rect 28441 15192 34671 15194
rect 28441 15136 28446 15192
rect 28502 15136 34610 15192
rect 34666 15136 34671 15192
rect 28441 15134 34671 15136
rect 28441 15131 28507 15134
rect 34605 15131 34671 15134
rect 29085 15058 29151 15061
rect 35525 15058 35591 15061
rect 29085 15056 35591 15058
rect 29085 15000 29090 15056
rect 29146 15000 35530 15056
rect 35586 15000 35591 15056
rect 29085 14998 35591 15000
rect 29085 14995 29151 14998
rect 35525 14995 35591 14998
rect 36077 15058 36143 15061
rect 39520 15058 40000 15088
rect 36077 15056 40000 15058
rect 36077 15000 36082 15056
rect 36138 15000 40000 15056
rect 36077 14998 40000 15000
rect 36077 14995 36143 14998
rect 39520 14968 40000 14998
rect 23289 14786 23355 14789
rect 27061 14786 27127 14789
rect 23289 14784 27127 14786
rect 23289 14728 23294 14784
rect 23350 14728 27066 14784
rect 27122 14728 27127 14784
rect 23289 14726 27127 14728
rect 23289 14723 23355 14726
rect 27061 14723 27127 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 37181 13970 37247 13973
rect 39520 13970 40000 14000
rect 37181 13968 40000 13970
rect 37181 13912 37186 13968
rect 37242 13912 40000 13968
rect 37181 13910 40000 13912
rect 37181 13907 37247 13910
rect 39520 13880 40000 13910
rect 25129 13698 25195 13701
rect 28533 13698 28599 13701
rect 28993 13698 29059 13701
rect 25129 13696 29059 13698
rect 25129 13640 25134 13696
rect 25190 13640 28538 13696
rect 28594 13640 28998 13696
rect 29054 13640 29059 13696
rect 25129 13638 29059 13640
rect 25129 13635 25195 13638
rect 28533 13635 28599 13638
rect 28993 13635 29059 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 24761 13018 24827 13021
rect 26141 13018 26207 13021
rect 24761 13016 26207 13018
rect 24761 12960 24766 13016
rect 24822 12960 26146 13016
rect 26202 12960 26207 13016
rect 24761 12958 26207 12960
rect 24761 12955 24827 12958
rect 26141 12955 26207 12958
rect 21173 12882 21239 12885
rect 24025 12882 24091 12885
rect 21173 12880 24091 12882
rect 21173 12824 21178 12880
rect 21234 12824 24030 12880
rect 24086 12824 24091 12880
rect 21173 12822 24091 12824
rect 21173 12819 21239 12822
rect 24025 12819 24091 12822
rect 34697 12746 34763 12749
rect 34654 12744 34763 12746
rect 34654 12688 34702 12744
rect 34758 12688 34763 12744
rect 34654 12683 34763 12688
rect 36537 12746 36603 12749
rect 39520 12746 40000 12776
rect 36537 12744 40000 12746
rect 36537 12688 36542 12744
rect 36598 12688 40000 12744
rect 36537 12686 40000 12688
rect 36537 12683 36603 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 34654 12477 34714 12683
rect 39520 12656 40000 12686
rect 34605 12472 34714 12477
rect 34605 12416 34610 12472
rect 34666 12416 34714 12472
rect 34605 12414 34714 12416
rect 34605 12411 34671 12414
rect 30005 12338 30071 12341
rect 36813 12338 36879 12341
rect 30005 12336 36879 12338
rect 30005 12280 30010 12336
rect 30066 12280 36818 12336
rect 36874 12280 36879 12336
rect 30005 12278 36879 12280
rect 30005 12275 30071 12278
rect 36813 12275 36879 12278
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 27613 11794 27679 11797
rect 30373 11794 30439 11797
rect 27613 11792 30439 11794
rect 27613 11736 27618 11792
rect 27674 11736 30378 11792
rect 30434 11736 30439 11792
rect 27613 11734 30439 11736
rect 27613 11731 27679 11734
rect 30373 11731 30439 11734
rect 31201 11658 31267 11661
rect 31661 11658 31727 11661
rect 31201 11656 31727 11658
rect 31201 11600 31206 11656
rect 31262 11600 31666 11656
rect 31722 11600 31727 11656
rect 31201 11598 31727 11600
rect 31201 11595 31267 11598
rect 31661 11595 31727 11598
rect 36261 11522 36327 11525
rect 39520 11522 40000 11552
rect 36261 11520 40000 11522
rect 36261 11464 36266 11520
rect 36322 11464 40000 11520
rect 36261 11462 40000 11464
rect 36261 11459 36327 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 39520 11432 40000 11462
rect 19568 11391 19888 11392
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 33041 10706 33107 10709
rect 36629 10706 36695 10709
rect 33041 10704 36695 10706
rect 33041 10648 33046 10704
rect 33102 10648 36634 10704
rect 36690 10648 36695 10704
rect 33041 10646 36695 10648
rect 33041 10643 33107 10646
rect 36629 10643 36695 10646
rect 34646 10508 34652 10572
rect 34716 10570 34722 10572
rect 34789 10570 34855 10573
rect 34716 10568 34855 10570
rect 34716 10512 34794 10568
rect 34850 10512 34855 10568
rect 34716 10510 34855 10512
rect 34716 10508 34722 10510
rect 34789 10507 34855 10510
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 36905 10298 36971 10301
rect 39520 10298 40000 10328
rect 36905 10296 40000 10298
rect 36905 10240 36910 10296
rect 36966 10240 40000 10296
rect 36905 10238 40000 10240
rect 36905 10235 36971 10238
rect 39520 10208 40000 10238
rect 34513 10026 34579 10029
rect 34513 10024 35404 10026
rect 34513 9968 34518 10024
rect 34574 9968 35404 10024
rect 34513 9966 35404 9968
rect 34513 9963 34579 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 35344 9757 35404 9966
rect 24577 9754 24643 9757
rect 27245 9754 27311 9757
rect 24577 9752 27311 9754
rect 24577 9696 24582 9752
rect 24638 9696 27250 9752
rect 27306 9696 27311 9752
rect 24577 9694 27311 9696
rect 24577 9691 24643 9694
rect 27245 9691 27311 9694
rect 35341 9752 35407 9757
rect 35617 9756 35683 9757
rect 35566 9754 35572 9756
rect 35341 9696 35346 9752
rect 35402 9696 35407 9752
rect 35341 9691 35407 9696
rect 35526 9694 35572 9754
rect 35636 9752 35683 9756
rect 35678 9696 35683 9752
rect 35566 9692 35572 9694
rect 35636 9692 35683 9696
rect 35617 9691 35683 9692
rect 35249 9618 35315 9621
rect 35893 9618 35959 9621
rect 35249 9616 35959 9618
rect 35249 9560 35254 9616
rect 35310 9560 35898 9616
rect 35954 9560 35959 9616
rect 35249 9558 35959 9560
rect 35249 9555 35315 9558
rect 35893 9555 35959 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 31569 9210 31635 9213
rect 34329 9210 34395 9213
rect 36905 9210 36971 9213
rect 31569 9208 36971 9210
rect 31569 9152 31574 9208
rect 31630 9152 34334 9208
rect 34390 9152 36910 9208
rect 36966 9152 36971 9208
rect 31569 9150 36971 9152
rect 31569 9147 31635 9150
rect 34329 9147 34395 9150
rect 36905 9147 36971 9150
rect 35433 9074 35499 9077
rect 39520 9074 40000 9104
rect 35433 9072 40000 9074
rect 35433 9016 35438 9072
rect 35494 9016 40000 9072
rect 35433 9014 40000 9016
rect 35433 9011 35499 9014
rect 39520 8984 40000 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 29913 8394 29979 8397
rect 31937 8394 32003 8397
rect 29913 8392 32003 8394
rect 29913 8336 29918 8392
rect 29974 8336 31942 8392
rect 31998 8336 32003 8392
rect 29913 8334 32003 8336
rect 29913 8331 29979 8334
rect 31937 8331 32003 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 34329 7986 34395 7989
rect 36721 7986 36787 7989
rect 34329 7984 36787 7986
rect 34329 7928 34334 7984
rect 34390 7928 36726 7984
rect 36782 7928 36787 7984
rect 34329 7926 36787 7928
rect 34329 7923 34395 7926
rect 36721 7923 36787 7926
rect 35893 7850 35959 7853
rect 39520 7850 40000 7880
rect 35893 7848 40000 7850
rect 35893 7792 35898 7848
rect 35954 7792 40000 7848
rect 35893 7790 40000 7792
rect 35893 7787 35959 7790
rect 39520 7760 40000 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 0 6762 480 6792
rect 565 6762 631 6765
rect 0 6760 631 6762
rect 0 6704 570 6760
rect 626 6704 631 6760
rect 0 6702 631 6704
rect 0 6672 480 6702
rect 565 6699 631 6702
rect 34789 6762 34855 6765
rect 34789 6760 35450 6762
rect 34789 6704 34794 6760
rect 34850 6704 35450 6760
rect 34789 6702 35450 6704
rect 34789 6699 34855 6702
rect 35390 6626 35450 6702
rect 39520 6626 40000 6656
rect 35390 6566 40000 6626
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 39520 6536 40000 6566
rect 34928 6495 35248 6496
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 565 5674 631 5677
rect 17493 5674 17559 5677
rect 565 5672 17559 5674
rect 565 5616 570 5672
rect 626 5616 17498 5672
rect 17554 5616 17559 5672
rect 565 5614 17559 5616
rect 565 5611 631 5614
rect 17493 5611 17559 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 39520 5402 40000 5432
rect 35390 5342 40000 5402
rect 34697 5266 34763 5269
rect 35390 5266 35450 5342
rect 39520 5312 40000 5342
rect 34697 5264 35450 5266
rect 34697 5208 34702 5264
rect 34758 5208 35450 5264
rect 34697 5206 35450 5208
rect 34697 5203 34763 5206
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 35709 4178 35775 4181
rect 39520 4178 40000 4208
rect 35709 4176 40000 4178
rect 35709 4120 35714 4176
rect 35770 4120 40000 4176
rect 35709 4118 40000 4120
rect 35709 4115 35775 4118
rect 39520 4088 40000 4118
rect 23289 4042 23355 4045
rect 23933 4042 23999 4045
rect 23289 4040 23999 4042
rect 23289 3984 23294 4040
rect 23350 3984 23938 4040
rect 23994 3984 23999 4040
rect 23289 3982 23999 3984
rect 23289 3979 23355 3982
rect 23933 3979 23999 3982
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 16665 3362 16731 3365
rect 31293 3362 31359 3365
rect 16665 3360 31359 3362
rect 16665 3304 16670 3360
rect 16726 3304 31298 3360
rect 31354 3304 31359 3360
rect 16665 3302 31359 3304
rect 16665 3299 16731 3302
rect 31293 3299 31359 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 35617 2954 35683 2957
rect 39520 2954 40000 2984
rect 35617 2952 40000 2954
rect 35617 2896 35622 2952
rect 35678 2896 40000 2952
rect 35617 2894 40000 2896
rect 35617 2891 35683 2894
rect 39520 2864 40000 2894
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 3325 2410 3391 2413
rect 33501 2410 33567 2413
rect 3325 2408 33567 2410
rect 3325 2352 3330 2408
rect 3386 2352 33506 2408
rect 33562 2352 33567 2408
rect 3325 2350 33567 2352
rect 3325 2347 3391 2350
rect 33501 2347 33567 2350
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 35433 1730 35499 1733
rect 39520 1730 40000 1760
rect 35433 1728 40000 1730
rect 35433 1672 35438 1728
rect 35494 1672 40000 1728
rect 35433 1670 40000 1672
rect 35433 1667 35499 1670
rect 39520 1640 40000 1670
rect 35801 642 35867 645
rect 39520 642 40000 672
rect 35801 640 40000 642
rect 35801 584 35806 640
rect 35862 584 40000 640
rect 35801 582 40000 584
rect 35801 579 35867 582
rect 39520 552 40000 582
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 8156 36484 8220 36548
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 24900 35532 24964 35596
rect 33180 34988 33244 35052
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 21588 34716 21652 34780
rect 24900 34776 24964 34780
rect 24900 34720 24950 34776
rect 24950 34720 24964 34776
rect 24900 34716 24964 34720
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 17908 33900 17972 33964
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 17908 33628 17972 33692
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 34652 23700 34716 23764
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 34652 20572 34716 20636
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 35572 16900 35636 16964
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 34652 10508 34716 10572
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 35572 9752 35636 9756
rect 35572 9696 35622 9752
rect 35622 9696 35636 9752
rect 35572 9692 35636 9696
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 37024 4528 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 19568 37568 19888 37584
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 8155 36548 8221 36549
rect 8155 36484 8156 36548
rect 8220 36484 8221 36548
rect 8155 36483 8221 36484
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 8158 35818 8218 36483
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 19568 35392 19888 36416
rect 34928 37024 35248 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 24899 35532 24900 35582
rect 24964 35532 24965 35582
rect 24899 35531 24965 35532
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 21590 34781 21650 34902
rect 24902 34781 24962 35531
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 21587 34780 21653 34781
rect 21587 34716 21588 34780
rect 21652 34716 21653 34780
rect 21587 34715 21653 34716
rect 24899 34780 24965 34781
rect 24899 34716 24900 34780
rect 24964 34716 24965 34780
rect 24899 34715 24965 34716
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 17907 33964 17973 33965
rect 17907 33900 17908 33964
rect 17972 33900 17973 33964
rect 17907 33899 17973 33900
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 17910 33693 17970 33899
rect 17907 33692 17973 33693
rect 17907 33628 17908 33692
rect 17972 33628 17973 33692
rect 17907 33627 17973 33628
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34651 23764 34717 23765
rect 34651 23700 34652 23764
rect 34716 23700 34717 23764
rect 34651 23699 34717 23700
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 34654 20637 34714 23699
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34651 20636 34717 20637
rect 34651 20572 34652 20636
rect 34716 20572 34717 20636
rect 34651 20571 34717 20572
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 34654 10573 34714 20571
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 35571 16964 35637 16965
rect 35571 16900 35572 16964
rect 35636 16900 35637 16964
rect 35571 16899 35637 16900
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34651 10572 34717 10573
rect 34651 10508 34652 10572
rect 34716 10508 34717 10572
rect 34651 10507 34717 10508
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 35574 9757 35634 16899
rect 35571 9756 35637 9757
rect 35571 9692 35572 9756
rect 35636 9692 35637 9756
rect 35571 9691 35637 9692
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
<< via4 >>
rect 8070 35582 8306 35818
rect 24814 35596 25050 35818
rect 24814 35582 24900 35596
rect 24900 35582 24964 35596
rect 24964 35582 25050 35596
rect 21502 34902 21738 35138
rect 33094 35052 33330 35138
rect 33094 34988 33180 35052
rect 33180 34988 33244 35052
rect 33244 34988 33330 35052
rect 33094 34902 33330 34988
<< metal5 >>
rect 8028 35818 25092 35860
rect 8028 35582 8070 35818
rect 8306 35582 24814 35818
rect 25050 35582 25092 35818
rect 8028 35540 25092 35582
rect 21460 35138 33372 35180
rect 21460 34902 21502 35138
rect 21738 34902 33094 35138
rect 33330 34902 33372 35138
rect 21460 34860 33372 34902
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8188 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_81
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_292
timestamp 1604681595
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_304
timestamp 1604681595
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1604681595
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_311
timestamp 1604681595
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1604681595
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_306
timestamp 1604681595
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1604681595
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1604681595
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_342
timestamp 1604681595
transform 1 0 32568 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_330
timestamp 1604681595
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_342
timestamp 1604681595
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 33304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 33856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_354
timestamp 1604681595
transform 1 0 33672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_358
timestamp 1604681595
transform 1 0 34040 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_370
timestamp 1604681595
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_354
timestamp 1604681595
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1604681595
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_373
timestamp 1604681595
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_385
timestamp 1604681595
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1604681595
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_391
timestamp 1604681595
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1604681595
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1604681595
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1604681595
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1604681595
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_300
timestamp 1604681595
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_312
timestamp 1604681595
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_324
timestamp 1604681595
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_337
timestamp 1604681595
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_349
timestamp 1604681595
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_361
timestamp 1604681595
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_373
timestamp 1604681595
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_385
timestamp 1604681595
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1604681595
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1604681595
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1604681595
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1604681595
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_330
timestamp 1604681595
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_342
timestamp 1604681595
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_354
timestamp 1604681595
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1604681595
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1604681595
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1604681595
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1604681595
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1604681595
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_300
timestamp 1604681595
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_312
timestamp 1604681595
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1604681595
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_337
timestamp 1604681595
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_349
timestamp 1604681595
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_361
timestamp 1604681595
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_373
timestamp 1604681595
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_385
timestamp 1604681595
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_398
timestamp 1604681595
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1604681595
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1604681595
transform 1 0 28060 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_299
timestamp 1604681595
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_303
timestamp 1604681595
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 29440 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_306
timestamp 1604681595
transform 1 0 29256 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_310
timestamp 1604681595
transform 1 0 29624 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_322
timestamp 1604681595
transform 1 0 30728 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 33212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_334
timestamp 1604681595
transform 1 0 31832 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_346
timestamp 1604681595
transform 1 0 32936 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_351
timestamp 1604681595
transform 1 0 33396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 33580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_359
timestamp 1604681595
transform 1 0 34132 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_355
timestamp 1604681595
transform 1 0 33764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 33948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_363
timestamp 1604681595
transform 1 0 34500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_367
timestamp 1604681595
transform 1 0 34868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_371
timestamp 1604681595
transform 1 0 35236 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 35052 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 35420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_375
timestamp 1604681595
transform 1 0 35604 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_387
timestamp 1604681595
transform 1 0 36708 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_399
timestamp 1604681595
transform 1 0 37812 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1604681595
transform 1 0 26588 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_282
timestamp 1604681595
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_290
timestamp 1604681595
transform 1 0 27784 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_286
timestamp 1604681595
transform 1 0 27416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 27600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 27232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_301
timestamp 1604681595
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1604681595
transform 1 0 28520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_300
timestamp 1604681595
transform 1 0 28704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 28796 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_288
timestamp 1604681595
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 29532 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 29808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 30176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_310
timestamp 1604681595
transform 1 0 29624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_314
timestamp 1604681595
transform 1 0 29992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_318
timestamp 1604681595
transform 1 0 30360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_306
timestamp 1604681595
transform 1 0 29256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_325
timestamp 1604681595
transform 1 0 31004 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_337
timestamp 1604681595
transform 1 0 32108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_335
timestamp 1604681595
transform 1 0 31924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_330
timestamp 1604681595
transform 1 0 31464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 31740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 31556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_349
timestamp 1604681595
transform 1 0 33212 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_347
timestamp 1604681595
transform 1 0 33028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_343
timestamp 1604681595
transform 1 0 32660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 32844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 32476 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 33212 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 31740 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_7_357
timestamp 1604681595
transform 1 0 33948 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_358
timestamp 1604681595
transform 1 0 34040 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_362
timestamp 1604681595
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_364
timestamp 1604681595
transform 1 0 34592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 34684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 34868 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 34868 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 36524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_376
timestamp 1604681595
transform 1 0 35696 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_388
timestamp 1604681595
transform 1 0 36800 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_383
timestamp 1604681595
transform 1 0 36340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_387
timestamp 1604681595
transform 1 0 36708 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_396
timestamp 1604681595
transform 1 0 37536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_398
timestamp 1604681595
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1604681595
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_399
timestamp 1604681595
transform 1 0 37812 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_282
timestamp 1604681595
transform 1 0 27048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 27232 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 28888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_300
timestamp 1604681595
transform 1 0 28704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_304
timestamp 1604681595
transform 1 0 29072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 29440 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 29256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_324
timestamp 1604681595
transform 1 0 30912 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 32476 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 32292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 31832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 31464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_332
timestamp 1604681595
transform 1 0 31648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_337
timestamp 1604681595
transform 1 0 32108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 34684 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 34132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_357
timestamp 1604681595
transform 1 0 33948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_361
timestamp 1604681595
transform 1 0 34316 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_381
timestamp 1604681595
transform 1 0 36156 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_393
timestamp 1604681595
transform 1 0 37260 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1604681595
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1604681595
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 26864 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 26496 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_274
timestamp 1604681595
transform 1 0 26312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1604681595
transform 1 0 26680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_296
timestamp 1604681595
transform 1 0 28336 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_301
timestamp 1604681595
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 29256 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_322
timestamp 1604681595
transform 1 0 30728 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 31464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 31280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 33120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_346
timestamp 1604681595
transform 1 0 32936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 34868 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 33672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_350
timestamp 1604681595
transform 1 0 33304 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_356
timestamp 1604681595
transform 1 0 33856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_360
timestamp 1604681595
transform 1 0 34224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 36524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 36892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_383
timestamp 1604681595
transform 1 0 36340 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_387
timestamp 1604681595
transform 1 0 36708 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_391
timestamp 1604681595
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1604681595
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_252
timestamp 1604681595
transform 1 0 24288 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_260
timestamp 1604681595
transform 1 0 25024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_265
timestamp 1604681595
transform 1 0 25484 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_273
timestamp 1604681595
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 28704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 28152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_296
timestamp 1604681595
transform 1 0 28336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 30820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_316
timestamp 1604681595
transform 1 0 30176 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_322
timestamp 1604681595
transform 1 0 30728 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_325
timestamp 1604681595
transform 1 0 31004 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 32108 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 33212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 31832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_333
timestamp 1604681595
transform 1 0 31740 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_346
timestamp 1604681595
transform 1 0 32936 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 33672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 35236 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_351
timestamp 1604681595
transform 1 0 33396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_363
timestamp 1604681595
transform 1 0 34500 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_369
timestamp 1604681595
transform 1 0 35052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_387
timestamp 1604681595
transform 1 0 36708 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_395
timestamp 1604681595
transform 1 0 37444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_398
timestamp 1604681595
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1604681595
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 24104 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_249
timestamp 1604681595
transform 1 0 24012 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_252
timestamp 1604681595
transform 1 0 24288 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1604681595
transform 1 0 24656 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_260
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 25300 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 27048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_279
timestamp 1604681595
transform 1 0 26772 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 27600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_284
timestamp 1604681595
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_297
timestamp 1604681595
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_301
timestamp 1604681595
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 29624 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 29440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 30636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_306
timestamp 1604681595
transform 1 0 29256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_319
timestamp 1604681595
transform 1 0 30452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_323
timestamp 1604681595
transform 1 0 30820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 32108 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 31924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 31556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 33212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_329
timestamp 1604681595
transform 1 0 31372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_333
timestamp 1604681595
transform 1 0 31740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_346
timestamp 1604681595
transform 1 0 32936 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 33672 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 35236 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_351
timestamp 1604681595
transform 1 0 33396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_358
timestamp 1604681595
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp 1604681595
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_367
timestamp 1604681595
transform 1 0 34868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 35420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 37076 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_389
timestamp 1604681595
transform 1 0 36892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1604681595
transform 1 0 37260 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1604681595
transform 1 0 38364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 24104 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 23736 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_245
timestamp 1604681595
transform 1 0 23644 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_248
timestamp 1604681595
transform 1 0 23920 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_259
timestamp 1604681595
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 26956 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_283
timestamp 1604681595
transform 1 0 27140 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 27692 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 27324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 29072 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 28704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_287
timestamp 1604681595
transform 1 0 27508 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_298
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_302
timestamp 1604681595
transform 1 0 28888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 29256 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 30820 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 30268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_315
timestamp 1604681595
transform 1 0 30084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_319
timestamp 1604681595
transform 1 0 30452 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_327
timestamp 1604681595
transform 1 0 31188 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 33212 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 32108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 32844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_333
timestamp 1604681595
transform 1 0 31740 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_341
timestamp 1604681595
transform 1 0 32476 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_347
timestamp 1604681595
transform 1 0 33028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 35144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 34224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 34776 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_358
timestamp 1604681595
transform 1 0 34040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_362
timestamp 1604681595
transform 1 0 34408 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_368
timestamp 1604681595
transform 1 0 34960 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 35420 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_372
timestamp 1604681595
transform 1 0 35328 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_389
timestamp 1604681595
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1604681595
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1604681595
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604681595
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 22724 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_228
timestamp 1604681595
transform 1 0 22080 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1604681595
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1604681595
transform 1 0 22908 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_241
timestamp 1604681595
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_255
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_262
timestamp 1604681595
transform 1 0 25208 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 24748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 23736 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_267
timestamp 1604681595
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_270
timestamp 1604681595
transform 1 0 25944 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_280
timestamp 1604681595
transform 1 0 26864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1604681595
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_277
timestamp 1604681595
transform 1 0 26588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_273
timestamp 1604681595
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 26956 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 27324 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 28336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_294
timestamp 1604681595
transform 1 0 28152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_298
timestamp 1604681595
transform 1 0 28520 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_304
timestamp 1604681595
transform 1 0 29072 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_290
timestamp 1604681595
transform 1 0 27784 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_302
timestamp 1604681595
transform 1 0 28888 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1604681595
transform 1 0 29992 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_312
timestamp 1604681595
transform 1 0 29808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_306
timestamp 1604681595
transform 1 0 29256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 29992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 29440 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_321
timestamp 1604681595
transform 1 0 30636 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_318
timestamp 1604681595
transform 1 0 30360 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_321
timestamp 1604681595
transform 1 0 30636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_316
timestamp 1604681595
transform 1 0 30176 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1604681595
transform 1 0 30452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 30452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 31004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 30820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 31004 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_327
timestamp 1604681595
transform 1 0 31188 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_337
timestamp 1604681595
transform 1 0 32108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_332
timestamp 1604681595
transform 1 0 31648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1604681595
transform 1 0 31832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 31464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 31832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_342
timestamp 1604681595
transform 1 0 32568 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_338
timestamp 1604681595
transform 1 0 32200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32384 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 32844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_349
timestamp 1604681595
transform 1 0 33212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_353
timestamp 1604681595
transform 1 0 33580 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_359
timestamp 1604681595
transform 1 0 34132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_354
timestamp 1604681595
transform 1 0 33672 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 33396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 33948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 33948 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_369
timestamp 1604681595
transform 1 0 35052 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_365
timestamp 1604681595
transform 1 0 34684 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_361
timestamp 1604681595
transform 1 0 34316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_367
timestamp 1604681595
transform 1 0 34868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_363
timestamp 1604681595
transform 1 0 34500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 34500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 35144 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 35144 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_377
timestamp 1604681595
transform 1 0 35788 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_372
timestamp 1604681595
transform 1 0 35328 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_379
timestamp 1604681595
transform 1 0 35972 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 36064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 35420 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_382
timestamp 1604681595
transform 1 0 36248 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_383
timestamp 1604681595
transform 1 0 36340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 36524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 36156 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 36708 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 36524 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1604681595
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_391
timestamp 1604681595
transform 1 0 37076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 37260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_395
timestamp 1604681595
transform 1 0 37444 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_398
timestamp 1604681595
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1604681595
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1604681595
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1604681595
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_228
timestamp 1604681595
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp 1604681595
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_235
timestamp 1604681595
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_261
timestamp 1604681595
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_265
timestamp 1604681595
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_285
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1604681595
transform 1 0 27692 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_293
timestamp 1604681595
transform 1 0 28060 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_301
timestamp 1604681595
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_306
timestamp 1604681595
transform 1 0 29256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 29440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_315
timestamp 1604681595
transform 1 0 30084 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_311
timestamp 1604681595
transform 1 0 29716 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 29900 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 30268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 30452 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_322
timestamp 1604681595
transform 1 0 30728 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 30820 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_327
timestamp 1604681595
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 31924 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 31740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 31372 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 32936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_331
timestamp 1604681595
transform 1 0 31556 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_344
timestamp 1604681595
transform 1 0 32752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_348
timestamp 1604681595
transform 1 0 33120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 33304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 33488 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_356
timestamp 1604681595
transform 1 0 33856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 34040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_360
timestamp 1604681595
transform 1 0 34224 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_367
timestamp 1604681595
transform 1 0 34868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_365
timestamp 1604681595
transform 1 0 34684 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 35236 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 35420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 37076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_389
timestamp 1604681595
transform 1 0 36892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1604681595
transform 1 0 37260 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1604681595
transform 1 0 38364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1604681595
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1604681595
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 22172 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 24380 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1604681595
transform 1 0 23644 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_262
timestamp 1604681595
transform 1 0 25208 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 27048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 26680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604681595
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1604681595
transform 1 0 28520 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 29256 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_322
timestamp 1604681595
transform 1 0 30728 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 32108 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 34500 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 34316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_353
timestamp 1604681595
transform 1 0 33580 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 36064 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 35512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_372
timestamp 1604681595
transform 1 0 35328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_376
timestamp 1604681595
transform 1 0 35696 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_385
timestamp 1604681595
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_398
timestamp 1604681595
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1604681595
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_226
timestamp 1604681595
transform 1 0 21896 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_229
timestamp 1604681595
transform 1 0 22172 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_233
timestamp 1604681595
transform 1 0 22540 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_237
timestamp 1604681595
transform 1 0 22908 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_254
timestamp 1604681595
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604681595
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_262
timestamp 1604681595
transform 1 0 25208 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 26680 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 26496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_270
timestamp 1604681595
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_274
timestamp 1604681595
transform 1 0 26312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 28612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_294
timestamp 1604681595
transform 1 0 28152 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1604681595
transform 1 0 28520 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_301
timestamp 1604681595
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 29256 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 30912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_322
timestamp 1604681595
transform 1 0 30728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_326
timestamp 1604681595
transform 1 0 31096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 31464 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 32476 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 32292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 31924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_333
timestamp 1604681595
transform 1 0 31740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1604681595
transform 1 0 32108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 34868 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 34132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_357
timestamp 1604681595
transform 1 0 33948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_361
timestamp 1604681595
transform 1 0 34316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 36432 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 36984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 35880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 36248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_376
timestamp 1604681595
transform 1 0 35696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_380
timestamp 1604681595
transform 1 0 36064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_388
timestamp 1604681595
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_392
timestamp 1604681595
transform 1 0 37168 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_404
timestamp 1604681595
transform 1 0 38272 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1604681595
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_222
timestamp 1604681595
transform 1 0 21528 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_226
timestamp 1604681595
transform 1 0 21896 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1604681595
transform 1 0 25208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_243
timestamp 1604681595
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_247
timestamp 1604681595
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_260
timestamp 1604681595
transform 1 0 25024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 26772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 27140 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_264
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_272
timestamp 1604681595
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_281
timestamp 1604681595
transform 1 0 26956 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 27324 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 29072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_301
timestamp 1604681595
transform 1 0 28796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 29716 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 29440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1604681595
transform 1 0 29256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_310
timestamp 1604681595
transform 1 0 29624 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_327
timestamp 1604681595
transform 1 0 31188 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 32752 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 32476 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_333
timestamp 1604681595
transform 1 0 31740 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_337
timestamp 1604681595
transform 1 0 32108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_343
timestamp 1604681595
transform 1 0 32660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 34868 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 35236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1604681595
transform 1 0 34684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_369
timestamp 1604681595
transform 1 0 35052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 35420 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1604681595
transform 1 0 36892 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_398
timestamp 1604681595
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1604681595
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1604681595
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_216
timestamp 1604681595
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1604681595
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 21160 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 22724 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 22540 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_255
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1604681595
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_254
timestamp 1604681595
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_prog_clk
timestamp 1604681595
transform 1 0 25208 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 25024 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_265
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_275
timestamp 1604681595
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 26220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 26588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 26772 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 27048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_284
timestamp 1604681595
transform 1 0 27232 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_292
timestamp 1604681595
transform 1 0 27968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_288
timestamp 1604681595
transform 1 0 27600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 27784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 27324 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_300
timestamp 1604681595
transform 1 0 28704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_294
timestamp 1604681595
transform 1 0 28152 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_301
timestamp 1604681595
transform 1 0 28796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_296
timestamp 1604681595
transform 1 0 28336 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 28888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 28520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 28152 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 28612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 29072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1604681595
transform 1 0 29348 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_310
timestamp 1604681595
transform 1 0 29624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1604681595
transform 1 0 29256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 29716 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 29440 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_325
timestamp 1604681595
transform 1 0 31004 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_321
timestamp 1604681595
transform 1 0 30636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_317
timestamp 1604681595
transform 1 0 30268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 30820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 30452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 29900 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_20_337
timestamp 1604681595
transform 1 0 32108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1604681595
transform 1 0 31648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_329
timestamp 1604681595
transform 1 0 31372 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1604681595
transform 1 0 31832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1604681595
transform 1 0 31464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 32016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_344
timestamp 1604681595
transform 1 0 32752 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_341
timestamp 1604681595
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_338
timestamp 1604681595
transform 1 0 32200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32568 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32568 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_352
timestamp 1604681595
transform 1 0 33488 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_359
timestamp 1604681595
transform 1 0 34132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_355
timestamp 1604681595
transform 1 0 33764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_351
timestamp 1604681595
transform 1 0 33396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 33948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 33580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_369
timestamp 1604681595
transform 1 0 35052 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_363
timestamp 1604681595
transform 1 0 34500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 35236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 34868 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 33580 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 37076 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35788 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 36524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 36892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_383
timestamp 1604681595
transform 1 0 36340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_387
timestamp 1604681595
transform 1 0 36708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_373
timestamp 1604681595
transform 1 0 35420 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_386
timestamp 1604681595
transform 1 0 36616 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_398
timestamp 1604681595
transform 1 0 37720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_394
timestamp 1604681595
transform 1 0 37352 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_398
timestamp 1604681595
transform 1 0 37720 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_394
timestamp 1604681595
transform 1 0 37352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 37536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1604681595
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1604681595
transform 1 0 38456 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_216
timestamp 1604681595
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_261
timestamp 1604681595
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 27048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 25300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_265
timestamp 1604681595
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_278
timestamp 1604681595
transform 1 0 26680 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_284
timestamp 1604681595
transform 1 0 27232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 27416 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_290
timestamp 1604681595
transform 1 0 27784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 27968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_294
timestamp 1604681595
transform 1 0 28152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 28336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 28520 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_301
timestamp 1604681595
transform 1 0 28796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 29900 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 29716 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 30912 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1604681595
transform 1 0 29256 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_310
timestamp 1604681595
transform 1 0 29624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_322
timestamp 1604681595
transform 1 0 30728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_326
timestamp 1604681595
transform 1 0 31096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_337
timestamp 1604681595
transform 1 0 32108 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_333
timestamp 1604681595
transform 1 0 31740 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 31280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_prog_clk
timestamp 1604681595
transform 1 0 31464 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_344
timestamp 1604681595
transform 1 0 32752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_340
timestamp 1604681595
transform 1 0 32384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 32936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_348
timestamp 1604681595
transform 1 0 33120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 34868 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_360
timestamp 1604681595
transform 1 0 34224 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_370
timestamp 1604681595
transform 1 0 35144 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_382
timestamp 1604681595
transform 1 0 36248 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_394
timestamp 1604681595
transform 1 0 37352 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1604681595
transform 1 0 38456 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 21344 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1604681595
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_222
timestamp 1604681595
transform 1 0 21528 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1604681595
transform 1 0 22632 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_238
timestamp 1604681595
transform 1 0 23000 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_243
timestamp 1604681595
transform 1 0 23460 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_249
timestamp 1604681595
transform 1 0 24012 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 27048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 26680 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 25852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_267
timestamp 1604681595
transform 1 0 25668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1604681595
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_280
timestamp 1604681595
transform 1 0 26864 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 28612 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 28244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1604681595
transform 1 0 27876 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1604681595
transform 1 0 28428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_303
timestamp 1604681595
transform 1 0 28980 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 29716 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 30268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 29256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 30636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_308
timestamp 1604681595
transform 1 0 29440 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_315
timestamp 1604681595
transform 1 0 30084 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_319
timestamp 1604681595
transform 1 0 30452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_323
timestamp 1604681595
transform 1 0 30820 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32200 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_329
timestamp 1604681595
transform 1 0 31372 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_335
timestamp 1604681595
transform 1 0 31924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_337
timestamp 1604681595
transform 1 0 32108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_347
timestamp 1604681595
transform 1 0 33028 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 34868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 35236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 34408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_359
timestamp 1604681595
transform 1 0 34132 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_364
timestamp 1604681595
transform 1 0 34592 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_369
timestamp 1604681595
transform 1 0 35052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_373
timestamp 1604681595
transform 1 0 35420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_385
timestamp 1604681595
transform 1 0 36524 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_398
timestamp 1604681595
transform 1 0 37720 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1604681595
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_214
timestamp 1604681595
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1604681595
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_221
timestamp 1604681595
transform 1 0 21436 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_233
timestamp 1604681595
transform 1 0 22540 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_237
timestamp 1604681595
transform 1 0 22908 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 23828 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_256
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_260
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 25392 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 27048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_280
timestamp 1604681595
transform 1 0 26864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_288
timestamp 1604681595
transform 1 0 27600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_284
timestamp 1604681595
transform 1 0 27232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 27416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 27784 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_298
timestamp 1604681595
transform 1 0 28520 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_294
timestamp 1604681595
transform 1 0 28152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 28336 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_302
timestamp 1604681595
transform 1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 28704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1604681595
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_314
timestamp 1604681595
transform 1 0 29992 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_310
timestamp 1604681595
transform 1 0 29624 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 29808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 29256 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_323
timestamp 1604681595
transform 1 0 30820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_319
timestamp 1604681595
transform 1 0 30452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 30636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 31004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 30268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 31188 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 32844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 33212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_343
timestamp 1604681595
transform 1 0 32660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_347
timestamp 1604681595
transform 1 0 33028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 33396 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 34868 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1604681595
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 34224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 33856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_354
timestamp 1604681595
transform 1 0 33672 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_358
timestamp 1604681595
transform 1 0 34040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_362
timestamp 1604681595
transform 1 0 34408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_376
timestamp 1604681595
transform 1 0 35696 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_388
timestamp 1604681595
transform 1 0 36800 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_400
timestamp 1604681595
transform 1 0 37904 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1604681595
transform 1 0 38456 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 19964 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 20332 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_207
timestamp 1604681595
transform 1 0 20148 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1604681595
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_231
timestamp 1604681595
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_prog_clk
timestamp 1604681595
transform 1 0 23920 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1604681595
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_243
timestamp 1604681595
transform 1 0 23460 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_255
timestamp 1604681595
transform 1 0 24564 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_267
timestamp 1604681595
transform 1 0 25668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1604681595
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 28244 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 27508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_285
timestamp 1604681595
transform 1 0 27324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_289
timestamp 1604681595
transform 1 0 27692 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1604681595
transform 1 0 29072 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 30268 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 29532 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 29900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_308
timestamp 1604681595
transform 1 0 29440 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_311
timestamp 1604681595
transform 1 0 29716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_315
timestamp 1604681595
transform 1 0 30084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_326
timestamp 1604681595
transform 1 0 31096 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 32200 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1604681595
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 31832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31464 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_332
timestamp 1604681595
transform 1 0 31648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_337
timestamp 1604681595
transform 1 0 32108 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 34408 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1604681595
transform 1 0 33672 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 36616 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 36064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_378
timestamp 1604681595
transform 1 0 35880 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_382
timestamp 1604681595
transform 1 0 36248 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_389
timestamp 1604681595
transform 1 0 36892 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1604681595
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_398
timestamp 1604681595
transform 1 0 37720 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1604681595
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_192
timestamp 1604681595
transform 1 0 18768 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 19964 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_199
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1604681595
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1604681595
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1604681595
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_241
timestamp 1604681595
transform 1 0 23276 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_251
timestamp 1604681595
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_255
timestamp 1604681595
transform 1 0 24564 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_260
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 25484 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 26956 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 26772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 26036 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_264
timestamp 1604681595
transform 1 0 25392 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1604681595
transform 1 0 26220 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1604681595
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 28612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1604681595
transform 1 0 28428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_301
timestamp 1604681595
transform 1 0 28796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 29532 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_306
timestamp 1604681595
transform 1 0 29256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_325
timestamp 1604681595
transform 1 0 31004 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 32016 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 31832 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 31464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_329
timestamp 1604681595
transform 1 0 31372 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_332
timestamp 1604681595
transform 1 0 31648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1604681595
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 34132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 34500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 35236 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_357
timestamp 1604681595
transform 1 0 33948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1604681595
transform 1 0 34316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_365
timestamp 1604681595
transform 1 0 34684 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_367
timestamp 1604681595
transform 1 0 34868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 35420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 37076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_389
timestamp 1604681595
transform 1 0 36892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1604681595
transform 1 0 37260 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1604681595
transform 1 0 38364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_195
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1604681595
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1604681595
transform 1 0 18400 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_194
timestamp 1604681595
transform 1 0 18952 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_199
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_218
timestamp 1604681595
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 19688 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1604681595
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21896 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_235
timestamp 1604681595
transform 1 0 22724 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_235
timestamp 1604681595
transform 1 0 22724 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_231
timestamp 1604681595
transform 1 0 22356 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 22540 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22908 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_239
timestamp 1604681595
transform 1 0 23092 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_249
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_241
timestamp 1604681595
transform 1 0 23276 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_262
timestamp 1604681595
transform 1 0 25208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24380 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 23828 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_26_270
timestamp 1604681595
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_266
timestamp 1604681595
transform 1 0 25576 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 25392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_283
timestamp 1604681595
transform 1 0 27140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_279
timestamp 1604681595
transform 1 0 26772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_283
timestamp 1604681595
transform 1 0 27140 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_280
timestamp 1604681595
transform 1 0 26864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604681595
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 26956 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 25300 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_27_287
timestamp 1604681595
transform 1 0 27508 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1604681595
transform 1 0 27600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 27324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 27784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 27968 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 27232 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_301
timestamp 1604681595
transform 1 0 28796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1604681595
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 28980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 28612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1604681595
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 28336 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 30544 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 29256 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 31096 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 31004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_312
timestamp 1604681595
transform 1 0 29808 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_324
timestamp 1604681595
transform 1 0 30912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_315
timestamp 1604681595
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_323
timestamp 1604681595
transform 1 0 30820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_327
timestamp 1604681595
transform 1 0 31188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_337
timestamp 1604681595
transform 1 0 32108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_328
timestamp 1604681595
transform 1 0 31280 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 31832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 31372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1604681595
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_347
timestamp 1604681595
transform 1 0 33028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_341
timestamp 1604681595
transform 1 0 32476 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 33212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 32292 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 31556 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 32752 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_27_351
timestamp 1604681595
transform 1 0 33396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 33580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_358
timestamp 1604681595
transform 1 0 34040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604681595
transform 1 0 33764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_363
timestamp 1604681595
transform 1 0 34500 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 34316 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_367
timestamp 1604681595
transform 1 0 34868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1604681595
transform 1 0 34684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 34868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1604681595
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_369
timestamp 1604681595
transform 1 0 35052 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 35236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 35236 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 35420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 36432 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 36800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_389
timestamp 1604681595
transform 1 0 36892 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_382
timestamp 1604681595
transform 1 0 36248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_386
timestamp 1604681595
transform 1 0 36616 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_390
timestamp 1604681595
transform 1 0 36984 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1604681595
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_398
timestamp 1604681595
transform 1 0 37720 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1604681595
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_402
timestamp 1604681595
transform 1 0 38088 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_406
timestamp 1604681595
transform 1 0 38456 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_196
timestamp 1604681595
transform 1 0 19136 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604681595
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 22540 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 22908 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_231
timestamp 1604681595
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_235
timestamp 1604681595
transform 1 0 22724 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_243
timestamp 1604681595
transform 1 0 23460 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_247
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_292
timestamp 1604681595
transform 1 0 27968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_304
timestamp 1604681595
transform 1 0 29072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 30268 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 29256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 29624 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_308
timestamp 1604681595
transform 1 0 29440 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_312
timestamp 1604681595
transform 1 0 29808 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_316
timestamp 1604681595
transform 1 0 30176 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_320
timestamp 1604681595
transform 1 0 30544 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 32108 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1604681595
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 31556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_328
timestamp 1604681595
transform 1 0 31280 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_333
timestamp 1604681595
transform 1 0 31740 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_346
timestamp 1604681595
transform 1 0 32936 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 34316 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_358
timestamp 1604681595
transform 1 0 34040 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_370
timestamp 1604681595
transform 1 0 35144 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 35880 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 35420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_375
timestamp 1604681595
transform 1 0 35604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_382
timestamp 1604681595
transform 1 0 36248 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1604681595
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_394
timestamp 1604681595
transform 1 0 37352 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_398
timestamp 1604681595
transform 1 0 37720 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1604681595
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_188
timestamp 1604681595
transform 1 0 18400 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1604681595
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_195
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 19780 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 21988 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 23092 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1604681595
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_223
timestamp 1604681595
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_241
timestamp 1604681595
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1604681595
transform 1 0 24012 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_259
timestamp 1604681595
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_255
timestamp 1604681595
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1604681595
transform 1 0 25300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_267
timestamp 1604681595
transform 1 0 25668 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1604681595
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 28704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 28336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 27968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_290
timestamp 1604681595
transform 1 0 27784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_294
timestamp 1604681595
transform 1 0 28152 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_298
timestamp 1604681595
transform 1 0 28520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_302
timestamp 1604681595
transform 1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_310
timestamp 1604681595
transform 1 0 29624 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_306
timestamp 1604681595
transform 1 0 29256 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 29440 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_314
timestamp 1604681595
transform 1 0 29992 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 29808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_320
timestamp 1604681595
transform 1 0 30544 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 30360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_324
timestamp 1604681595
transform 1 0 30912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 30728 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 31096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32660 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 32108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1604681595
transform 1 0 31280 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_336
timestamp 1604681595
transform 1 0 32016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_339
timestamp 1604681595
transform 1 0 32292 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1604681595
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 34040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 34408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 33672 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_352
timestamp 1604681595
transform 1 0 33488 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_356
timestamp 1604681595
transform 1 0 33856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_360
timestamp 1604681595
transform 1 0 34224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_364
timestamp 1604681595
transform 1 0 34592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_367
timestamp 1604681595
transform 1 0 34868 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 35604 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 35972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 36340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_377
timestamp 1604681595
transform 1 0 35788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_381
timestamp 1604681595
transform 1 0 36156 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_385
timestamp 1604681595
transform 1 0 36524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_397
timestamp 1604681595
transform 1 0 37628 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1604681595
transform 1 0 38364 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1604681595
transform 1 0 14720 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1604681595
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_158
timestamp 1604681595
transform 1 0 15640 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_170
timestamp 1604681595
transform 1 0 16744 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_182
timestamp 1604681595
transform 1 0 17848 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_194
timestamp 1604681595
transform 1 0 18952 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 22540 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_231
timestamp 1604681595
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_235
timestamp 1604681595
transform 1 0 22724 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24748 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24472 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_248
timestamp 1604681595
transform 1 0 23920 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_252
timestamp 1604681595
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_256
timestamp 1604681595
transform 1 0 24656 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 1604681595
transform 1 0 25944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_266
timestamp 1604681595
transform 1 0 25576 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_272
timestamp 1604681595
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_280
timestamp 1604681595
transform 1 0 26864 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 28704 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 28060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_291
timestamp 1604681595
transform 1 0 27876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1604681595
transform 1 0 28244 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_299
timestamp 1604681595
transform 1 0 28612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 30360 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 29900 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1604681595
transform 1 0 29532 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_315
timestamp 1604681595
transform 1 0 30084 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_327
timestamp 1604681595
transform 1 0 31188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1604681595
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 33028 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 31372 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_331
timestamp 1604681595
transform 1 0 31556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_335
timestamp 1604681595
transform 1 0 31924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_337
timestamp 1604681595
transform 1 0 32108 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_345
timestamp 1604681595
transform 1 0 32844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_349
timestamp 1604681595
transform 1 0 33212 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 34040 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_357
timestamp 1604681595
transform 1 0 33948 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_367
timestamp 1604681595
transform 1 0 34868 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35604 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 35420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1604681595
transform 1 0 36432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1604681595
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_396
timestamp 1604681595
transform 1 0 37536 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_398
timestamp 1604681595
transform 1 0 37720 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1604681595
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 14536 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_143
timestamp 1604681595
transform 1 0 14260 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1604681595
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_170
timestamp 1604681595
transform 1 0 16744 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 17480 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 18216 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1604681595
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_192
timestamp 1604681595
transform 1 0 18768 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 19964 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_198
timestamp 1604681595
transform 1 0 19320 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_201
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 22172 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 21896 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_221
timestamp 1604681595
transform 1 0 21436 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1604681595
transform 1 0 21804 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_228
timestamp 1604681595
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp 1604681595
transform 1 0 22540 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_237
timestamp 1604681595
transform 1 0 22908 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24196 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25208 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_241
timestamp 1604681595
transform 1 0 23276 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_260
timestamp 1604681595
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 26864 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 25760 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_264
timestamp 1604681595
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_272
timestamp 1604681595
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1604681595
transform 1 0 26680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_284
timestamp 1604681595
transform 1 0 27232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 27416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_288
timestamp 1604681595
transform 1 0 27600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 27784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_292
timestamp 1604681595
transform 1 0 27968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 28152 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1604681595
transform 1 0 28428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 28612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_301
timestamp 1604681595
transform 1 0 28796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1604681595
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 29900 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 29716 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1604681595
transform 1 0 29256 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_310
timestamp 1604681595
transform 1 0 29624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 32936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 32568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_334
timestamp 1604681595
transform 1 0 31832 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_344
timestamp 1604681595
transform 1 0 32752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_348
timestamp 1604681595
transform 1 0 33120 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604681595
transform 1 0 33764 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1604681595
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 35236 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 33304 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_352
timestamp 1604681595
transform 1 0 33488 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_358
timestamp 1604681595
transform 1 0 34040 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_367
timestamp 1604681595
transform 1 0 34868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 35420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 37076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_389
timestamp 1604681595
transform 1 0 36892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1604681595
transform 1 0 37260 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1604681595
transform 1 0 38364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_137
timestamp 1604681595
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1604681595
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1604681595
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_198
timestamp 1604681595
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_210
timestamp 1604681595
transform 1 0 20424 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604681595
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 21896 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 21712 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_220
timestamp 1604681595
transform 1 0 21344 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_235
timestamp 1604681595
transform 1 0 22724 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23276 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_243
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_247
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1604681595
transform 1 0 24840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_262
timestamp 1604681595
transform 1 0 25208 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 26036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 27048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_270
timestamp 1604681595
transform 1 0 25944 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1604681595
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_280
timestamp 1604681595
transform 1 0 26864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 27600 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 27416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_284
timestamp 1604681595
transform 1 0 27232 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_304
timestamp 1604681595
transform 1 0 29072 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 29808 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 29256 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 29624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_308
timestamp 1604681595
transform 1 0 29440 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 32936 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1604681595
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 32752 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 32292 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_328
timestamp 1604681595
transform 1 0 31280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_337
timestamp 1604681595
transform 1 0 32108 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_341
timestamp 1604681595
transform 1 0 32476 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 35052 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_367
timestamp 1604681595
transform 1 0 34868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_371
timestamp 1604681595
transform 1 0 35236 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35604 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 35420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_384
timestamp 1604681595
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1604681595
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_396
timestamp 1604681595
transform 1 0 37536 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_398
timestamp 1604681595
transform 1 0 37720 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1604681595
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_131
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_127
timestamp 1604681595
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 13892 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 13340 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 15548 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_155
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_158
timestamp 1604681595
transform 1 0 15640 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 15824 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_162
timestamp 1604681595
transform 1 0 16008 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 16100 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1604681595
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 16192 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk
timestamp 1604681595
transform 1 0 18400 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 17480 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_176
timestamp 1604681595
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_180
timestamp 1604681595
transform 1 0 17664 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_186
timestamp 1604681595
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 19504 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 21160 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 20516 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_208
timestamp 1604681595
transform 1 0 20240 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1604681595
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_226
timestamp 1604681595
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_222
timestamp 1604681595
transform 1 0 21528 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_227
timestamp 1604681595
transform 1 0 21988 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 22264 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_34_246
timestamp 1604681595
transform 1 0 23736 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_255
timestamp 1604681595
transform 1 0 24564 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_260
timestamp 1604681595
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_267
timestamp 1604681595
transform 1 0 25668 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_268
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_264
timestamp 1604681595
transform 1 0 25392 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 26036 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 26036 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1604681595
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_280
timestamp 1604681595
transform 1 0 26864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 27048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 26772 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_284
timestamp 1604681595
transform 1 0 27232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 27416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 27600 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_301
timestamp 1604681595
transform 1 0 28796 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1604681595
transform 1 0 28244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_301
timestamp 1604681595
transform 1 0 28796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1604681595
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 28612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 28612 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_305
timestamp 1604681595
transform 1 0 29164 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1604681595
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 29256 0 1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 29624 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 29256 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_327
timestamp 1604681595
transform 1 0 31188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_308
timestamp 1604681595
transform 1 0 29440 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_326
timestamp 1604681595
transform 1 0 31096 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_332
timestamp 1604681595
transform 1 0 31648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_331
timestamp 1604681595
transform 1 0 31556 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 31464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 31740 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1604681595
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 32108 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_347
timestamp 1604681595
transform 1 0 33028 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_344
timestamp 1604681595
transform 1 0 32752 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_340
timestamp 1604681595
transform 1 0 32384 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 32844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 33212 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 31924 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_34_351
timestamp 1604681595
transform 1 0 33396 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_359
timestamp 1604681595
transform 1 0 34132 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_355
timestamp 1604681595
transform 1 0 33764 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_351
timestamp 1604681595
transform 1 0 33396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 33948 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 33580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_367
timestamp 1604681595
transform 1 0 34868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_363
timestamp 1604681595
transform 1 0 34500 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 34316 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1604681595
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 35052 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 33488 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 36156 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 37260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 35604 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 36708 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_385
timestamp 1604681595
transform 1 0 36524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_389
timestamp 1604681595
transform 1 0 36892 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_373
timestamp 1604681595
transform 1 0 35420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_377
timestamp 1604681595
transform 1 0 35788 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_384
timestamp 1604681595
transform 1 0 36432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1604681595
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_396
timestamp 1604681595
transform 1 0 37536 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_404
timestamp 1604681595
transform 1 0 38272 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_396
timestamp 1604681595
transform 1 0 37536 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_398
timestamp 1604681595
transform 1 0 37720 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1604681595
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 12972 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 12788 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_110
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 14628 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_145
timestamp 1604681595
transform 1 0 14444 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 15180 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 16744 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_162
timestamp 1604681595
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1604681595
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_174
timestamp 1604681595
transform 1 0 17112 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 17296 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_178
timestamp 1604681595
transform 1 0 17480 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1604681595
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_200
timestamp 1604681595
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_204
timestamp 1604681595
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_213
timestamp 1604681595
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_217
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1604681595
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 23828 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_258
timestamp 1604681595
transform 1 0 24840 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 25576 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_282
timestamp 1604681595
transform 1 0 27048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_286
timestamp 1604681595
transform 1 0 27416 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 27600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 27232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 27784 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_294
timestamp 1604681595
transform 1 0 28152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 28336 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_302
timestamp 1604681595
transform 1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 28704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1604681595
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 29256 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 30912 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_322
timestamp 1604681595
transform 1 0 30728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_326
timestamp 1604681595
transform 1 0 31096 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 31464 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 33212 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 33028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 31280 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_339
timestamp 1604681595
transform 1 0 32292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_345
timestamp 1604681595
transform 1 0 32844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 34960 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1604681595
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 34224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_358
timestamp 1604681595
transform 1 0 34040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_362
timestamp 1604681595
transform 1 0 34408 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_367
timestamp 1604681595
transform 1 0 34868 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 36616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_384
timestamp 1604681595
transform 1 0 36432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_388
timestamp 1604681595
transform 1 0 36800 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_400
timestamp 1604681595
transform 1 0 37904 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1604681595
transform 1 0 38456 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 12880 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_144
timestamp 1604681595
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_148
timestamp 1604681595
transform 1 0 14720 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 16836 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_163
timestamp 1604681595
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_167
timestamp 1604681595
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 18400 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_186
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 19780 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1604681595
transform 1 0 19228 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_201
timestamp 1604681595
transform 1 0 19596 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_205
timestamp 1604681595
transform 1 0 19964 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1604681595
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_231
timestamp 1604681595
transform 1 0 22356 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 23460 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25116 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_259
timestamp 1604681595
transform 1 0 24932 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_268
timestamp 1604681595
transform 1 0 25760 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1604681595
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_280
timestamp 1604681595
transform 1 0 26864 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 27600 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 28612 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 28428 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_291
timestamp 1604681595
transform 1 0 27876 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 30176 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 29624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 29992 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_308
timestamp 1604681595
transform 1 0 29440 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_312
timestamp 1604681595
transform 1 0 29808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_319
timestamp 1604681595
transform 1 0 30452 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_327
timestamp 1604681595
transform 1 0 31188 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 33212 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1604681595
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 31464 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 33028 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1604681595
transform 1 0 31648 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_337
timestamp 1604681595
transform 1 0 32108 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_345
timestamp 1604681595
transform 1 0 32844 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 34776 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 34224 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 34592 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_358
timestamp 1604681595
transform 1 0 34040 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1604681595
transform 1 0 34408 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_382
timestamp 1604681595
transform 1 0 36248 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1604681595
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_394
timestamp 1604681595
transform 1 0 37352 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_398
timestamp 1604681595
transform 1 0 37720 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1604681595
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_103
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_115
timestamp 1604681595
transform 1 0 11684 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1604681595
transform 1 0 12052 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_131
timestamp 1604681595
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13892 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1604681595
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_152
timestamp 1604681595
transform 1 0 15088 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15456 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16468 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_165
timestamp 1604681595
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1604681595
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_173
timestamp 1604681595
transform 1 0 17020 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 18308 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_181
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19964 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 20332 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20700 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_203
timestamp 1604681595
transform 1 0 19780 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_207
timestamp 1604681595
transform 1 0 20148 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_211
timestamp 1604681595
transform 1 0 20516 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_215
timestamp 1604681595
transform 1 0 20884 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_223
timestamp 1604681595
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_236
timestamp 1604681595
transform 1 0 22816 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1604681595
transform 1 0 24380 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1604681595
transform 1 0 24196 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_249
timestamp 1604681595
transform 1 0 24012 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 26864 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1604681595
transform 1 0 26220 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1604681595
transform 1 0 26772 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_288
timestamp 1604681595
transform 1 0 27600 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_284
timestamp 1604681595
transform 1 0 27232 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 27416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_292
timestamp 1604681595
transform 1 0 27968 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 28060 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_295
timestamp 1604681595
transform 1 0 28244 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_301
timestamp 1604681595
transform 1 0 28796 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 28612 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1604681595
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 29256 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_prog_clk
timestamp 1604681595
transform 1 0 31188 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 30268 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 30636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_315
timestamp 1604681595
transform 1 0 30084 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_319
timestamp 1604681595
transform 1 0 30452 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_323
timestamp 1604681595
transform 1 0 30820 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_334
timestamp 1604681595
transform 1 0 31832 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_330
timestamp 1604681595
transform 1 0 31464 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1604681595
transform 1 0 31648 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_345
timestamp 1604681595
transform 1 0 32844 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_341
timestamp 1604681595
transform 1 0 32476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_338
timestamp 1604681595
transform 1 0 32200 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 32292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 32660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 33028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 33212 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 34868 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1604681595
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 34224 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 34592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_358
timestamp 1604681595
transform 1 0 34040 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_362
timestamp 1604681595
transform 1 0 34408 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 36524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_383
timestamp 1604681595
transform 1 0 36340 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_387
timestamp 1604681595
transform 1 0 36708 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_399
timestamp 1604681595
transform 1 0 37812 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_104
timestamp 1604681595
transform 1 0 10672 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 12512 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_116
timestamp 1604681595
transform 1 0 11776 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1604681595
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1604681595
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16836 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_163
timestamp 1604681595
transform 1 0 16100 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_168
timestamp 1604681595
transform 1 0 16560 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19136 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 18308 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17848 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_180
timestamp 1604681595
transform 1 0 17664 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_184
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_189
timestamp 1604681595
transform 1 0 18492 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1604681595
transform 1 0 18860 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_212
timestamp 1604681595
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 1604681595
transform 1 0 21436 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1604681595
transform 1 0 21252 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1604681595
transform 1 0 21620 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_229
timestamp 1604681595
transform 1 0 22172 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 24656 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24288 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_241
timestamp 1604681595
transform 1 0 23276 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1604681595
transform 1 0 24012 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_254
timestamp 1604681595
transform 1 0 24472 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_272
timestamp 1604681595
transform 1 0 26128 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 28888 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 28060 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1604681595
transform 1 0 27600 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_292
timestamp 1604681595
transform 1 0 27968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_296
timestamp 1604681595
transform 1 0 28336 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 30544 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_318
timestamp 1604681595
transform 1 0 30360 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_322
timestamp 1604681595
transform 1 0 30728 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 33028 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1604681595
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_334
timestamp 1604681595
transform 1 0 31832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_337
timestamp 1604681595
transform 1 0 32108 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_345
timestamp 1604681595
transform 1 0 32844 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 34132 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 33580 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 33948 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_351
timestamp 1604681595
transform 1 0 33396 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_355
timestamp 1604681595
transform 1 0 33764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 36340 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 35788 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_375
timestamp 1604681595
transform 1 0 35604 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_379
timestamp 1604681595
transform 1 0 35972 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_386
timestamp 1604681595
transform 1 0 36616 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1604681595
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_394
timestamp 1604681595
transform 1 0 37352 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_398
timestamp 1604681595
transform 1 0 37720 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1604681595
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_64
timestamp 1604681595
transform 1 0 6992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_71
timestamp 1604681595
transform 1 0 7636 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_67
timestamp 1604681595
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_75
timestamp 1604681595
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_70
timestamp 1604681595
transform 1 0 7544 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 7820 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_82
timestamp 1604681595
transform 1 0 8648 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_79
timestamp 1604681595
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_83
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_97
timestamp 1604681595
transform 1 0 10028 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_90
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_95
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_100
timestamp 1604681595
transform 1 0 10304 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_109
timestamp 1604681595
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_105
timestamp 1604681595
transform 1 0 10764 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 10580 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_prog_clk
timestamp 1604681595
transform 1 0 11316 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_125
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_119
timestamp 1604681595
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_129
timestamp 1604681595
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_138
timestamp 1604681595
transform 1 0 13800 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_133
timestamp 1604681595
transform 1 0 13340 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_133
timestamp 1604681595
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_151
timestamp 1604681595
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 13708 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_39_157
timestamp 1604681595
transform 1 0 15548 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_153
timestamp 1604681595
transform 1 0 15180 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 15916 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_168
timestamp 1604681595
transform 1 0 16560 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_163
timestamp 1604681595
transform 1 0 16100 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_164
timestamp 1604681595
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_185
timestamp 1604681595
transform 1 0 18124 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_180
timestamp 1604681595
transform 1 0 17664 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_175
timestamp 1604681595
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_189
timestamp 1604681595
transform 1 0 18492 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_192
timestamp 1604681595
transform 1 0 18768 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_188
timestamp 1604681595
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_206
timestamp 1604681595
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_206
timestamp 1604681595
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_202
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 19228 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_40_210
timestamp 1604681595
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1604681595
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1604681595
transform 1 0 20792 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_39_234
timestamp 1604681595
transform 1 0 22632 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_224
timestamp 1604681595
transform 1 0 21712 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_236
timestamp 1604681595
transform 1 0 22816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1604681595
transform 1 0 23920 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_249
timestamp 1604681595
transform 1 0 24012 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_252
timestamp 1604681595
transform 1 0 24288 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_prog_clk
timestamp 1604681595
transform 1 0 24656 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24288 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_261
timestamp 1604681595
transform 1 0 25116 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_265
timestamp 1604681595
transform 1 0 25484 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_268
timestamp 1604681595
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 25944 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 25392 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_273
timestamp 1604681595
transform 1 0 26220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_276
timestamp 1604681595
transform 1 0 26496 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_272
timestamp 1604681595
transform 1 0 26128 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1604681595
transform 1 0 26312 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_294
timestamp 1604681595
transform 1 0 28152 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_286
timestamp 1604681595
transform 1 0 27416 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 27232 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 27232 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_303
timestamp 1604681595
transform 1 0 28980 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_299
timestamp 1604681595
transform 1 0 28612 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_298
timestamp 1604681595
transform 1 0 28520 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 29072 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 28336 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 28704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 28888 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1604681595
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_287
timestamp 1604681595
transform 1 0 27508 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 29900 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 29256 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 29440 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 30912 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_306
timestamp 1604681595
transform 1 0 29256 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_310
timestamp 1604681595
transform 1 0 29624 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_322
timestamp 1604681595
transform 1 0 30728 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_326
timestamp 1604681595
transform 1 0 31096 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_322
timestamp 1604681595
transform 1 0 30728 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_332
timestamp 1604681595
transform 1 0 31648 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_336
timestamp 1604681595
transform 1 0 32016 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1604681595
transform 1 0 31464 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1604681595
transform 1 0 31832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 31280 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 31464 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1604681595
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_341
timestamp 1604681595
transform 1 0 32476 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_339
timestamp 1604681595
transform 1 0 32292 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 32108 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 32108 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 32568 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_349
timestamp 1604681595
transform 1 0 33212 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_346
timestamp 1604681595
transform 1 0 32936 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 33120 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_357
timestamp 1604681595
transform 1 0 33948 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_353
timestamp 1604681595
transform 1 0 33580 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_358
timestamp 1604681595
transform 1 0 34040 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_350
timestamp 1604681595
transform 1 0 33304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 33764 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 33488 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 33396 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 34224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 33672 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_362
timestamp 1604681595
transform 1 0 34408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1604681595
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 34868 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 34224 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 36432 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 36432 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 35880 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_376
timestamp 1604681595
transform 1 0 35696 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_380
timestamp 1604681595
transform 1 0 36064 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_386
timestamp 1604681595
transform 1 0 36616 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_376
timestamp 1604681595
transform 1 0 35696 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_388
timestamp 1604681595
transform 1 0 36800 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1604681595
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_398
timestamp 1604681595
transform 1 0 37720 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1604681595
transform 1 0 38456 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_396
timestamp 1604681595
transform 1 0 37536 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_398
timestamp 1604681595
transform 1 0 37720 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1604681595
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 7360 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_84
timestamp 1604681595
transform 1 0 8832 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 9568 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_94
timestamp 1604681595
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 14812 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_138
timestamp 1604681595
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_142
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_146
timestamp 1604681595
transform 1 0 14536 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_prog_clk
timestamp 1604681595
transform 1 0 17020 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16468 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_165
timestamp 1604681595
transform 1 0 16284 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1604681595
transform 1 0 16652 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18308 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_176
timestamp 1604681595
transform 1 0 17296 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_180
timestamp 1604681595
transform 1 0 17664 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19872 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19688 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_200
timestamp 1604681595
transform 1 0 19504 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604681595
transform 1 0 22080 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 21528 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 21896 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_224
timestamp 1604681595
transform 1 0 21712 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_231
timestamp 1604681595
transform 1 0 22356 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_239
timestamp 1604681595
transform 1 0 23092 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 24472 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 24196 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23828 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_249
timestamp 1604681595
transform 1 0 24012 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_253
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_270
timestamp 1604681595
transform 1 0 25944 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_274
timestamp 1604681595
transform 1 0 26312 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 27416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_288
timestamp 1604681595
transform 1 0 27600 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 27784 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_292
timestamp 1604681595
transform 1 0 27968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 28152 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_296
timestamp 1604681595
transform 1 0 28336 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 28612 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_301
timestamp 1604681595
transform 1 0 28796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 28980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1604681595
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 29256 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 30912 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_322
timestamp 1604681595
transform 1 0 30728 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_326
timestamp 1604681595
transform 1 0 31096 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 31464 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 31280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 32476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 33120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_339
timestamp 1604681595
transform 1 0 32292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_343
timestamp 1604681595
transform 1 0 32660 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_347
timestamp 1604681595
transform 1 0 33028 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 33672 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 34868 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1604681595
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 34224 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 33488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_350
timestamp 1604681595
transform 1 0 33304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_358
timestamp 1604681595
transform 1 0 34040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_362
timestamp 1604681595
transform 1 0 34408 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 36432 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 36984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 35880 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 36248 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_376
timestamp 1604681595
transform 1 0 35696 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_380
timestamp 1604681595
transform 1 0 36064 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_388
timestamp 1604681595
transform 1 0 36800 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_392
timestamp 1604681595
transform 1 0 37168 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_404
timestamp 1604681595
transform 1 0 38272 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 7084 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_62
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_81
timestamp 1604681595
transform 1 0 8556 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10488 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_89
timestamp 1604681595
transform 1 0 9292 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_97
timestamp 1604681595
transform 1 0 10028 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_100
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12420 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_120
timestamp 1604681595
transform 1 0 12144 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_129
timestamp 1604681595
transform 1 0 12972 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_135
timestamp 1604681595
transform 1 0 13524 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_145
timestamp 1604681595
transform 1 0 14444 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 16928 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_170
timestamp 1604681595
transform 1 0 16744 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_174
timestamp 1604681595
transform 1 0 17112 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 18124 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 17296 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_178
timestamp 1604681595
transform 1 0 17480 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_184
timestamp 1604681595
transform 1 0 18032 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_189
timestamp 1604681595
transform 1 0 18492 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_193
timestamp 1604681595
transform 1 0 18860 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 20884 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1604681595
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20608 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_206
timestamp 1604681595
transform 1 0 20056 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_210
timestamp 1604681595
transform 1 0 20424 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 23184 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 21436 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21804 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_219
timestamp 1604681595
transform 1 0 21252 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_223
timestamp 1604681595
transform 1 0 21620 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1604681595
transform 1 0 21988 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_239
timestamp 1604681595
transform 1 0 23092 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 24196 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_243
timestamp 1604681595
transform 1 0 23460 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_247
timestamp 1604681595
transform 1 0 23828 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1604681595
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 26772 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 27140 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_267
timestamp 1604681595
transform 1 0 25668 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_276
timestamp 1604681595
transform 1 0 26496 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_281
timestamp 1604681595
transform 1 0 26956 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 27784 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 27508 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 29164 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_285
timestamp 1604681595
transform 1 0 27324 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_289
timestamp 1604681595
transform 1 0 27692 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_299
timestamp 1604681595
transform 1 0 28612 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 29348 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_323
timestamp 1604681595
transform 1 0 30820 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 32292 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1604681595
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_prog_clk
timestamp 1604681595
transform 1 0 31556 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 32844 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 33212 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_334
timestamp 1604681595
transform 1 0 31832 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_337
timestamp 1604681595
transform 1 0 32108 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_343
timestamp 1604681595
transform 1 0 32660 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_347
timestamp 1604681595
transform 1 0 33028 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 33396 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 34960 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 34408 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 34776 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_360
timestamp 1604681595
transform 1 0 34224 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_364
timestamp 1604681595
transform 1 0 34592 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_384
timestamp 1604681595
transform 1 0 36432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1604681595
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_396
timestamp 1604681595
transform 1 0 37536 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_398
timestamp 1604681595
transform 1 0 37720 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1604681595
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604681595
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1604681595
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1604681595
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1604681595
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1604681595
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 6900 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1604681595
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1604681595
transform 1 0 5796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1604681595
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_62
timestamp 1604681595
transform 1 0 6808 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_79
timestamp 1604681595
transform 1 0 8372 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_83
timestamp 1604681595
transform 1 0 8740 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 10120 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 9936 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 9568 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_91
timestamp 1604681595
transform 1 0 9476 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_94
timestamp 1604681595
transform 1 0 9752 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1604681595
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 11776 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_114
timestamp 1604681595
transform 1 0 11592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_118
timestamp 1604681595
transform 1 0 11960 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15088 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14352 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 13984 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_132
timestamp 1604681595
transform 1 0 13248 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_142
timestamp 1604681595
transform 1 0 14168 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_146
timestamp 1604681595
transform 1 0 14536 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_150
timestamp 1604681595
transform 1 0 14904 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 17020 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_170
timestamp 1604681595
transform 1 0 16744 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 18032 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 19136 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1604681595
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 18584 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 18952 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_175
timestamp 1604681595
transform 1 0 17204 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_188
timestamp 1604681595
transform 1 0 18400 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_192
timestamp 1604681595
transform 1 0 18768 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 20792 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 20608 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 20240 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19688 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_200
timestamp 1604681595
transform 1 0 19504 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1604681595
transform 1 0 19872 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_210
timestamp 1604681595
transform 1 0 20424 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_235
timestamp 1604681595
transform 1 0 22724 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 24104 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1604681595
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 23920 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_241
timestamp 1604681595
transform 1 0 23276 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_245
timestamp 1604681595
transform 1 0 23644 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 26772 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 26496 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_271
timestamp 1604681595
transform 1 0 26036 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_275
timestamp 1604681595
transform 1 0 26404 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_278
timestamp 1604681595
transform 1 0 26680 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1604681595
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 27784 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 28152 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 28980 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 28612 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_288
timestamp 1604681595
transform 1 0 27600 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_292
timestamp 1604681595
transform 1 0 27968 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_296
timestamp 1604681595
transform 1 0 28336 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_301
timestamp 1604681595
transform 1 0 28796 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 29440 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 31096 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_306
timestamp 1604681595
transform 1 0 29256 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_324
timestamp 1604681595
transform 1 0 30912 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 32752 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 31648 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 32200 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 32568 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 31464 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_328
timestamp 1604681595
transform 1 0 31280 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_336
timestamp 1604681595
transform 1 0 32016 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_340
timestamp 1604681595
transform 1 0 32384 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1604681595
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 35236 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 34592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 33764 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 34132 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_353
timestamp 1604681595
transform 1 0 33580 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_357
timestamp 1604681595
transform 1 0 33948 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_361
timestamp 1604681595
transform 1 0 34316 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_367
timestamp 1604681595
transform 1 0 34868 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 36616 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 35420 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 36064 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 37168 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 36432 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_378
timestamp 1604681595
transform 1 0 35880 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_382
timestamp 1604681595
transform 1 0 36248 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1604681595
transform 1 0 36984 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604681595
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_394
timestamp 1604681595
transform 1 0 37352 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1604681595
transform 1 0 38456 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604681595
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604681595
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1604681595
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1604681595
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604681595
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1604681595
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 6900 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1604681595
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_56
timestamp 1604681595
transform 1 0 6256 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_62
timestamp 1604681595
transform 1 0 6808 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8556 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_79
timestamp 1604681595
transform 1 0 8372 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_83
timestamp 1604681595
transform 1 0 8740 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11040 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1604681595
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10304 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_91
timestamp 1604681595
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_93
timestamp 1604681595
transform 1 0 9660 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_99
timestamp 1604681595
transform 1 0 10212 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_102
timestamp 1604681595
transform 1 0 10488 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_106
timestamp 1604681595
transform 1 0 10856 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12696 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_124
timestamp 1604681595
transform 1 0 12512 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_128
timestamp 1604681595
transform 1 0 12880 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_140
timestamp 1604681595
transform 1 0 13984 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_148
timestamp 1604681595
transform 1 0 14720 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 17020 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1604681595
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_154
timestamp 1604681595
transform 1 0 15272 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_165
timestamp 1604681595
transform 1 0 16284 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18676 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1604681595
transform 1 0 17388 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_189
timestamp 1604681595
transform 1 0 18492 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_193
timestamp 1604681595
transform 1 0 18860 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1604681595
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20424 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1604681595
transform 1 0 20056 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_212
timestamp 1604681595
transform 1 0 20608 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_231
timestamp 1604681595
transform 1 0 22356 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 24104 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23736 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_243
timestamp 1604681595
transform 1 0 23460 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_248
timestamp 1604681595
transform 1 0 23920 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_252
timestamp 1604681595
transform 1 0 24288 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 26496 0 -1 26656
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1604681595
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25852 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_267
timestamp 1604681595
transform 1 0 25668 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_271
timestamp 1604681595
transform 1 0 26036 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 28888 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_297
timestamp 1604681595
transform 1 0 28428 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_301
timestamp 1604681595
transform 1 0 28796 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_304
timestamp 1604681595
transform 1 0 29072 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 29440 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 29256 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_324
timestamp 1604681595
transform 1 0 30912 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 32108 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1604681595
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 31648 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 33120 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 31280 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_330
timestamp 1604681595
transform 1 0 31464 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_334
timestamp 1604681595
transform 1 0 31832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_346
timestamp 1604681595
transform 1 0 32936 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 33672 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 35236 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 34868 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 33488 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_350
timestamp 1604681595
transform 1 0 33304 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_363
timestamp 1604681595
transform 1 0 34500 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_369
timestamp 1604681595
transform 1 0 35052 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 36892 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_387
timestamp 1604681595
transform 1 0 36708 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_391
timestamp 1604681595
transform 1 0 37076 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604681595
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1604681595
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_398
timestamp 1604681595
transform 1 0 37720 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1604681595
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604681595
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 1564 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 1932 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1604681595
transform 1 0 1380 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_7
timestamp 1604681595
transform 1 0 1748 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_11
timestamp 1604681595
transform 1 0 2116 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_23
timestamp 1604681595
transform 1 0 3220 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_35
timestamp 1604681595
transform 1 0 4324 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1604681595
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_47
timestamp 1604681595
transform 1 0 5428 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_62
timestamp 1604681595
transform 1 0 6808 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8188 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 7176 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_68
timestamp 1604681595
transform 1 0 7360 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_73
timestamp 1604681595
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_86
timestamp 1604681595
transform 1 0 9016 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 9936 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9568 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_94
timestamp 1604681595
transform 1 0 9752 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_98
timestamp 1604681595
transform 1 0 10120 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1604681595
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11684 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1604681595
transform 1 0 11500 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_117
timestamp 1604681595
transform 1 0 11868 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 14168 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 13432 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14628 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_132
timestamp 1604681595
transform 1 0 13248 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_136
timestamp 1604681595
transform 1 0 13616 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_145
timestamp 1604681595
transform 1 0 14444 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1604681595
transform 1 0 14812 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15364 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 17020 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15180 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_171
timestamp 1604681595
transform 1 0 16836 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1604681595
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_175
timestamp 1604681595
transform 1 0 17204 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_184
timestamp 1604681595
transform 1 0 18032 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_192
timestamp 1604681595
transform 1 0 18768 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_195
timestamp 1604681595
transform 1 0 19044 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1604681595
transform 1 0 19412 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20424 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19872 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_202
timestamp 1604681595
transform 1 0 19688 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_206
timestamp 1604681595
transform 1 0 20056 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22448 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22816 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22080 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23184 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_226
timestamp 1604681595
transform 1 0 21896 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_230
timestamp 1604681595
transform 1 0 22264 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_234
timestamp 1604681595
transform 1 0 22632 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_238
timestamp 1604681595
transform 1 0 23000 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1604681595
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_242
timestamp 1604681595
transform 1 0 23368 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_245
timestamp 1604681595
transform 1 0 23644 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_258
timestamp 1604681595
transform 1 0 24840 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_262
timestamp 1604681595
transform 1 0 25208 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 25576 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_282
timestamp 1604681595
transform 1 0 27048 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1604681595
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_prog_clk
timestamp 1604681595
transform 1 0 27784 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1604681595
transform 1 0 28244 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 28612 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_293
timestamp 1604681595
transform 1 0 28060 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1604681595
transform 1 0 28428 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_301
timestamp 1604681595
transform 1 0 28796 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 29440 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 31096 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_306
timestamp 1604681595
transform 1 0 29256 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_324
timestamp 1604681595
transform 1 0 30912 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 31648 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 33212 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 31464 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 33028 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 32660 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_328
timestamp 1604681595
transform 1 0 31280 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_341
timestamp 1604681595
transform 1 0 32476 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_345
timestamp 1604681595
transform 1 0 32844 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 34868 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1604681595
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 34224 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_358
timestamp 1604681595
transform 1 0 34040 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_362
timestamp 1604681595
transform 1 0 34408 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 36432 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 35880 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 36248 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_376
timestamp 1604681595
transform 1 0 35696 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_380
timestamp 1604681595
transform 1 0 36064 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1604681595
transform 1 0 37260 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604681595
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 37444 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_397
timestamp 1604681595
transform 1 0 37628 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1604681595
transform 1 0 38364 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604681595
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604681595
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 1748 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 2116 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_19
timestamp 1604681595
transform 1 0 2852 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1604681595
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_9
timestamp 1604681595
transform 1 0 1932 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_13
timestamp 1604681595
transform 1 0 2300 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1604681595
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 4048 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1604681595
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_25
timestamp 1604681595
transform 1 0 3404 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_31
timestamp 1604681595
transform 1 0 3956 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_34
timestamp 1604681595
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_38
timestamp 1604681595
transform 1 0 4600 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1604681595
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1604681595
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_56
timestamp 1604681595
transform 1 0 6256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_64
timestamp 1604681595
transform 1 0 6992 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_50
timestamp 1604681595
transform 1 0 5704 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_58
timestamp 1604681595
transform 1 0 6440 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1604681595
transform 1 0 6808 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_68
timestamp 1604681595
transform 1 0 7360 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 7176 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 7544 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 7728 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_85
timestamp 1604681595
transform 1 0 8924 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_81
timestamp 1604681595
transform 1 0 8556 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_82
timestamp 1604681595
transform 1 0 8648 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 9108 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 8740 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 7176 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_47_97
timestamp 1604681595
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_89
timestamp 1604681595
transform 1 0 9292 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1604681595
transform 1 0 9660 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 9476 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1604681595
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 9936 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 9660 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_101
timestamp 1604681595
transform 1 0 10396 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_107
timestamp 1604681595
transform 1 0 10948 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_104
timestamp 1604681595
transform 1 0 10672 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_100
timestamp 1604681595
transform 1 0 10304 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 10212 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11040 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1604681595
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12696 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_124
timestamp 1604681595
transform 1 0 12512 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_128
timestamp 1604681595
transform 1 0 12880 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_114
timestamp 1604681595
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_118
timestamp 1604681595
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_136
timestamp 1604681595
transform 1 0 13616 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_132
timestamp 1604681595
transform 1 0 13248 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 13432 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 13248 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_152
timestamp 1604681595
transform 1 0 15088 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_148
timestamp 1604681595
transform 1 0 14720 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_144
timestamp 1604681595
transform 1 0 14352 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_152
timestamp 1604681595
transform 1 0 15088 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_148
timestamp 1604681595
transform 1 0 14720 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14536 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14904 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_136
timestamp 1604681595
transform 1 0 13616 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_162
timestamp 1604681595
transform 1 0 16008 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_158
timestamp 1604681595
transform 1 0 15640 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_154
timestamp 1604681595
transform 1 0 15272 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1604681595
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_165
timestamp 1604681595
transform 1 0 16284 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_166
timestamp 1604681595
transform 1 0 16376 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16192 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 16468 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1604681595
transform 1 0 16652 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_171
timestamp 1604681595
transform 1 0 16836 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1604681595
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18860 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_183
timestamp 1604681595
transform 1 0 17940 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_195
timestamp 1604681595
transform 1 0 19044 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_181
timestamp 1604681595
transform 1 0 17756 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_184
timestamp 1604681595
transform 1 0 18032 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_192
timestamp 1604681595
transform 1 0 18768 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_195
timestamp 1604681595
transform 1 0 19044 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_204
timestamp 1604681595
transform 1 0 19872 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_199
timestamp 1604681595
transform 1 0 19412 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_206
timestamp 1604681595
transform 1 0 20056 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20056 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1604681595
transform 1 0 19596 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_208
timestamp 1604681595
transform 1 0 20240 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_210
timestamp 1604681595
transform 1 0 20424 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20516 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1604681595
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20700 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 22356 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_224
timestamp 1604681595
transform 1 0 21712 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1604681595
transform 1 0 22080 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_229
timestamp 1604681595
transform 1 0 22172 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_233
timestamp 1604681595
transform 1 0 22540 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1604681595
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_241
timestamp 1604681595
transform 1 0 23276 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_241
timestamp 1604681595
transform 1 0 23276 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_245
timestamp 1604681595
transform 1 0 23644 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_247
timestamp 1604681595
transform 1 0 23828 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_258
timestamp 1604681595
transform 1 0 24840 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_255
timestamp 1604681595
transform 1 0 24564 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_251
timestamp 1604681595
transform 1 0 24196 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24656 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_262
timestamp 1604681595
transform 1 0 25208 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 25024 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1604681595
transform 1 0 26036 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_267
timestamp 1604681595
transform 1 0 25668 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 25392 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_282
timestamp 1604681595
transform 1 0 27048 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_279
timestamp 1604681595
transform 1 0 26772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 26956 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1604681595
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 26496 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_283
timestamp 1604681595
transform 1 0 27140 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 25576 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1604681595
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 27232 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_295
timestamp 1604681595
transform 1 0 28244 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1604681595
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_298
timestamp 1604681595
transform 1 0 28520 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_302
timestamp 1604681595
transform 1 0 28888 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 29624 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 30084 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 29900 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 29532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 29440 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1604681595
transform 1 0 29348 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_326
timestamp 1604681595
transform 1 0 31096 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_306
timestamp 1604681595
transform 1 0 29256 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_311
timestamp 1604681595
transform 1 0 29716 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_335
timestamp 1604681595
transform 1 0 31924 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_331
timestamp 1604681595
transform 1 0 31556 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_332
timestamp 1604681595
transform 1 0 31648 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 31464 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 31832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 31740 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 32108 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1604681595
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 32108 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_46_346
timestamp 1604681595
transform 1 0 32936 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 32292 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_348
timestamp 1604681595
transform 1 0 33120 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 33212 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_360
timestamp 1604681595
transform 1 0 34224 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_356
timestamp 1604681595
transform 1 0 33856 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_352
timestamp 1604681595
transform 1 0 33488 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_357
timestamp 1604681595
transform 1 0 33948 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_351
timestamp 1604681595
transform 1 0 33396 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 34040 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 33672 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 33304 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 34040 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_367
timestamp 1604681595
transform 1 0 34868 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_366
timestamp 1604681595
transform 1 0 34776 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1604681595
transform 1 0 34408 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 34592 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 34960 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 34592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1604681595
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 35144 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 34960 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 36800 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 36616 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_386
timestamp 1604681595
transform 1 0 36616 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_390
timestamp 1604681595
transform 1 0 36984 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_384
timestamp 1604681595
transform 1 0 36432 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_388
timestamp 1604681595
transform 1 0 36800 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604681595
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604681595
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1604681595
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_396
timestamp 1604681595
transform 1 0 37536 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_398
timestamp 1604681595
transform 1 0 37720 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1604681595
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_400
timestamp 1604681595
transform 1 0 37904 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1604681595
transform 1 0 38456 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1748 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604681595
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1604681595
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4048 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1604681595
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_23
timestamp 1604681595
transform 1 0 3220 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1604681595
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5704 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_48
timestamp 1604681595
transform 1 0 5520 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_52
timestamp 1604681595
transform 1 0 5888 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_64
timestamp 1604681595
transform 1 0 6992 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 8004 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 7728 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 7360 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_70
timestamp 1604681595
transform 1 0 7544 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_74
timestamp 1604681595
transform 1 0 7912 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_84
timestamp 1604681595
transform 1 0 8832 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 9660 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1604681595
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10212 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10580 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_97
timestamp 1604681595
transform 1 0 10028 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_101
timestamp 1604681595
transform 1 0 10396 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_105
timestamp 1604681595
transform 1 0 10764 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 13156 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12972 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_123
timestamp 1604681595
transform 1 0 12420 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_127
timestamp 1604681595
transform 1 0 12788 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14352 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 1604681595
transform 1 0 13524 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1604681595
transform 1 0 13892 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_142
timestamp 1604681595
transform 1 0 14168 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_146
timestamp 1604681595
transform 1 0 14536 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_150
timestamp 1604681595
transform 1 0 14904 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604681595
transform 1 0 16836 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1604681595
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 16284 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_163
timestamp 1604681595
transform 1 0 16100 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_167
timestamp 1604681595
transform 1 0 16468 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_174
timestamp 1604681595
transform 1 0 17112 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_186
timestamp 1604681595
transform 1 0 18216 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_190
timestamp 1604681595
transform 1 0 18584 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_193
timestamp 1604681595
transform 1 0 18860 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1604681595
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_206
timestamp 1604681595
transform 1 0 20056 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_210
timestamp 1604681595
transform 1 0 20424 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 23184 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_231
timestamp 1604681595
transform 1 0 22356 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_239
timestamp 1604681595
transform 1 0 23092 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 24196 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_243
timestamp 1604681595
transform 1 0 23460 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_247
timestamp 1604681595
transform 1 0 23828 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 26496 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1604681595
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_267
timestamp 1604681595
transform 1 0 25668 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1604681595
transform 1 0 26036 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_292
timestamp 1604681595
transform 1 0 27968 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_304
timestamp 1604681595
transform 1 0 29072 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 29808 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 29624 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 32384 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1604681595
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 31464 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_328
timestamp 1604681595
transform 1 0 31280 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_332
timestamp 1604681595
transform 1 0 31648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_337
timestamp 1604681595
transform 1 0 32108 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 34592 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 34408 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_356
timestamp 1604681595
transform 1 0 33856 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_380
timestamp 1604681595
transform 1 0 36064 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_392
timestamp 1604681595
transform 1 0 37168 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604681595
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1604681595
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_396
timestamp 1604681595
transform 1 0 37536 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_398
timestamp 1604681595
transform 1 0 37720 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1604681595
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2668 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604681595
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2024 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1656 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp 1604681595
transform 1 0 1380 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_8
timestamp 1604681595
transform 1 0 1840 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_12
timestamp 1604681595
transform 1 0 2208 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_16
timestamp 1604681595
transform 1 0 2576 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 4324 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_33
timestamp 1604681595
transform 1 0 4140 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_37
timestamp 1604681595
transform 1 0 4508 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_41
timestamp 1604681595
transform 1 0 4876 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1604681595
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 6440 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 6992 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_53
timestamp 1604681595
transform 1 0 5980 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_57
timestamp 1604681595
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_60
timestamp 1604681595
transform 1 0 6624 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_62
timestamp 1604681595
transform 1 0 6808 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 7728 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 7544 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_66
timestamp 1604681595
transform 1 0 7176 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9936 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 9660 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10948 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_88
timestamp 1604681595
transform 1 0 9200 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_92
timestamp 1604681595
transform 1 0 9568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_95
timestamp 1604681595
transform 1 0 9844 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_105
timestamp 1604681595
transform 1 0 10764 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_109
timestamp 1604681595
transform 1 0 11132 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1604681595
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11316 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1604681595
transform 1 0 11500 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_118
timestamp 1604681595
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 15088 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13432 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_132
timestamp 1604681595
transform 1 0 13248 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_136
timestamp 1604681595
transform 1 0 13616 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_149
timestamp 1604681595
transform 1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15640 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 15456 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_154
timestamp 1604681595
transform 1 0 15272 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_174
timestamp 1604681595
transform 1 0 17112 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_178
timestamp 1604681595
transform 1 0 17480 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17296 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_184
timestamp 1604681595
transform 1 0 18032 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1604681595
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 18400 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_194
timestamp 1604681595
transform 1 0 18952 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_190
timestamp 1604681595
transform 1 0 18584 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18768 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 19136 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 19320 0 1 28832
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1604681595
transform 1 0 21988 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21436 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21804 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_219
timestamp 1604681595
transform 1 0 21252 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_223
timestamp 1604681595
transform 1 0 21620 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_230
timestamp 1604681595
transform 1 0 22264 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 23644 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 24748 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1604681595
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24564 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24196 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_249
timestamp 1604681595
transform 1 0 24012 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_253
timestamp 1604681595
transform 1 0 24380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 26956 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 26772 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 26404 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_273
timestamp 1604681595
transform 1 0 26220 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_277
timestamp 1604681595
transform 1 0 26588 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1604681595
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_290
timestamp 1604681595
transform 1 0 27784 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_302
timestamp 1604681595
transform 1 0 28888 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_306
timestamp 1604681595
transform 1 0 29256 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_318
timestamp 1604681595
transform 1 0 30360 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_326
timestamp 1604681595
transform 1 0 31096 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 31464 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 31280 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_346
timestamp 1604681595
transform 1 0 32936 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 34868 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1604681595
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 33488 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 34224 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 33856 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_354
timestamp 1604681595
transform 1 0 33672 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_358
timestamp 1604681595
transform 1 0 34040 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_362
timestamp 1604681595
transform 1 0 34408 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 35880 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_376
timestamp 1604681595
transform 1 0 35696 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_380
timestamp 1604681595
transform 1 0 36064 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_392
timestamp 1604681595
transform 1 0 37168 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604681595
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_404
timestamp 1604681595
transform 1 0 38272 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604681595
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1604681595
transform 1 0 1380 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_11
timestamp 1604681595
transform 1 0 2116 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 4232 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1604681595
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_23
timestamp 1604681595
transform 1 0 3220 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_32
timestamp 1604681595
transform 1 0 4048 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 6440 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5888 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 6256 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_50
timestamp 1604681595
transform 1 0 5704 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_54
timestamp 1604681595
transform 1 0 6072 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 8464 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_74
timestamp 1604681595
transform 1 0 7912 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_78
timestamp 1604681595
transform 1 0 8280 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1604681595
transform 1 0 8648 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_86
timestamp 1604681595
transform 1 0 9016 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 9660 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1604681595
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_109
timestamp 1604681595
transform 1 0 11132 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11316 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12052 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_113
timestamp 1604681595
transform 1 0 11500 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_121
timestamp 1604681595
transform 1 0 12236 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_125
timestamp 1604681595
transform 1 0 12604 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 14444 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_143
timestamp 1604681595
transform 1 0 14260 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_147
timestamp 1604681595
transform 1 0 14628 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_151
timestamp 1604681595
transform 1 0 14996 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 15640 0 -1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1604681595
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_154
timestamp 1604681595
transform 1 0 15272 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 18032 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 18400 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_179
timestamp 1604681595
transform 1 0 17572 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1604681595
transform 1 0 17940 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_186
timestamp 1604681595
transform 1 0 18216 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_190
timestamp 1604681595
transform 1 0 18584 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_194
timestamp 1604681595
transform 1 0 18952 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1604681595
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_206
timestamp 1604681595
transform 1 0 20056 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_231
timestamp 1604681595
transform 1 0 22356 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24564 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 24380 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_243
timestamp 1604681595
transform 1 0 23460 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_251
timestamp 1604681595
transform 1 0 24196 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1604681595
transform 1 0 26496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1604681595
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 26956 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25576 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1604681595
transform 1 0 25392 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_268
timestamp 1604681595
transform 1 0 25760 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_274
timestamp 1604681595
transform 1 0 26312 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_279
timestamp 1604681595
transform 1 0 26772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_283
timestamp 1604681595
transform 1 0 27140 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_295
timestamp 1604681595
transform 1 0 28244 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_307
timestamp 1604681595
transform 1 0 29348 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_319
timestamp 1604681595
transform 1 0 30452 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1604681595
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 32384 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_331
timestamp 1604681595
transform 1 0 31556 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_335
timestamp 1604681595
transform 1 0 31924 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_337
timestamp 1604681595
transform 1 0 32108 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_342
timestamp 1604681595
transform 1 0 32568 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 33488 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 35144 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_350
timestamp 1604681595
transform 1 0 33304 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_368
timestamp 1604681595
transform 1 0 34960 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 35696 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_372
timestamp 1604681595
transform 1 0 35328 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_380
timestamp 1604681595
transform 1 0 36064 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_392
timestamp 1604681595
transform 1 0 37168 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604681595
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1604681595
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_396
timestamp 1604681595
transform 1 0 37536 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_398
timestamp 1604681595
transform 1 0 37720 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1604681595
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2944 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604681595
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2760 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2392 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 1564 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1604681595
transform 1 0 1380 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_7
timestamp 1604681595
transform 1 0 1748 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_13
timestamp 1604681595
transform 1 0 2300 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_16
timestamp 1604681595
transform 1 0 2576 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 4508 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 4324 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 3956 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_29
timestamp 1604681595
transform 1 0 3772 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_33
timestamp 1604681595
transform 1 0 4140 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1604681595
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_53
timestamp 1604681595
transform 1 0 5980 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1604681595
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 8464 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 7820 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 8280 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_71
timestamp 1604681595
transform 1 0 7636 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_75
timestamp 1604681595
transform 1 0 8004 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 10580 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_96
timestamp 1604681595
transform 1 0 9936 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_101
timestamp 1604681595
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12604 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1604681595
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_114
timestamp 1604681595
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_118
timestamp 1604681595
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_123
timestamp 1604681595
transform 1 0 12420 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14168 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 13616 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 13984 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_134
timestamp 1604681595
transform 1 0 13432 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_138
timestamp 1604681595
transform 1 0 13800 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15824 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_158
timestamp 1604681595
transform 1 0 15640 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_162
timestamp 1604681595
transform 1 0 16008 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1604681595
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_175
timestamp 1604681595
transform 1 0 17204 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_179
timestamp 1604681595
transform 1 0 17572 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20700 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20516 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20148 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_205
timestamp 1604681595
transform 1 0 19964 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_209
timestamp 1604681595
transform 1 0 20332 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 22540 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_229
timestamp 1604681595
transform 1 0 22172 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_235
timestamp 1604681595
transform 1 0 22724 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 23644 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 24748 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1604681595
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 24564 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 24196 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23368 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1604681595
transform 1 0 23276 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_249
timestamp 1604681595
transform 1 0 24012 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_253
timestamp 1604681595
transform 1 0 24380 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 26956 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 26496 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_273
timestamp 1604681595
transform 1 0 26220 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_278
timestamp 1604681595
transform 1 0 26680 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1604681595
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 27508 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_285
timestamp 1604681595
transform 1 0 27324 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_289
timestamp 1604681595
transform 1 0 27692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_301
timestamp 1604681595
transform 1 0 28796 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_306
timestamp 1604681595
transform 1 0 29256 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_318
timestamp 1604681595
transform 1 0 30360 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 32384 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 32200 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_330
timestamp 1604681595
transform 1 0 31464 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1604681595
transform 1 0 33212 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1604681595
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 35236 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_361
timestamp 1604681595
transform 1 0 34316 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_365
timestamp 1604681595
transform 1 0 34684 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_367
timestamp 1604681595
transform 1 0 34868 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 35420 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 35972 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_377
timestamp 1604681595
transform 1 0 35788 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_381
timestamp 1604681595
transform 1 0 36156 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1604681595
transform 1 0 37260 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604681595
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1604681595
transform 1 0 38364 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_7
timestamp 1604681595
transform 1 0 1748 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1604681595
transform 1 0 1380 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 1932 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 1564 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604681595
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604681595
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_19
timestamp 1604681595
transform 1 0 2852 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_19
timestamp 1604681595
transform 1 0 2852 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1604681595
transform 1 0 2484 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_11
timestamp 1604681595
transform 1 0 2116 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2944 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 1380 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_53_23
timestamp 1604681595
transform 1 0 3220 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1604681595
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_26
timestamp 1604681595
transform 1 0 3496 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_22
timestamp 1604681595
transform 1 0 3128 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 3404 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1604681595
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_40
timestamp 1604681595
transform 1 0 4784 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_36
timestamp 1604681595
transform 1 0 4416 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_38
timestamp 1604681595
transform 1 0 4600 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_32
timestamp 1604681595
transform 1 0 4048 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 4784 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 4600 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 4232 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_42
timestamp 1604681595
transform 1 0 4968 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_53
timestamp 1604681595
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1604681595
transform 1 0 6348 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_62
timestamp 1604681595
transform 1 0 6808 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 6992 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1604681595
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 6808 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 5336 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_53_70
timestamp 1604681595
transform 1 0 7544 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_66
timestamp 1604681595
transform 1 0 7176 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 8096 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_86
timestamp 1604681595
transform 1 0 9016 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_82
timestamp 1604681595
transform 1 0 8648 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_78
timestamp 1604681595
transform 1 0 8280 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_83
timestamp 1604681595
transform 1 0 8740 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_78
timestamp 1604681595
transform 1 0 8280 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 8464 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_prog_clk
timestamp 1604681595
transform 1 0 8464 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1604681595
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_97
timestamp 1604681595
transform 1 0 10028 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_89
timestamp 1604681595
transform 1 0 9292 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 9200 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1604681595
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 9660 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 9384 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_103
timestamp 1604681595
transform 1 0 10580 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_99
timestamp 1604681595
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_101
timestamp 1604681595
transform 1 0 10396 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 10580 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 10212 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10764 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 10948 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 10764 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_53_114
timestamp 1604681595
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 11224 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_118
timestamp 1604681595
transform 1 0 11960 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1604681595
transform 1 0 12236 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1604681595
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 12420 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_131
timestamp 1604681595
transform 1 0 13156 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_127
timestamp 1604681595
transform 1 0 12788 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_127
timestamp 1604681595
transform 1 0 12788 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12972 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 12972 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 13156 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_52_136
timestamp 1604681595
transform 1 0 13616 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 13524 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_143
timestamp 1604681595
transform 1 0 14260 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_139
timestamp 1604681595
transform 1 0 13892 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14168 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 14076 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 14352 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_151
timestamp 1604681595
transform 1 0 14996 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_147
timestamp 1604681595
transform 1 0 14628 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_147
timestamp 1604681595
transform 1 0 14628 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 14720 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_160
timestamp 1604681595
transform 1 0 15824 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_155
timestamp 1604681595
transform 1 0 15364 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_154
timestamp 1604681595
transform 1 0 15272 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 15180 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 16008 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1604681595
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 15456 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_168
timestamp 1604681595
transform 1 0 16560 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_164
timestamp 1604681595
transform 1 0 16192 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_173
timestamp 1604681595
transform 1 0 17020 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 16836 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16376 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_prog_clk
timestamp 1604681595
transform 1 0 17020 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15548 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_53_184
timestamp 1604681595
transform 1 0 18032 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_180
timestamp 1604681595
transform 1 0 17664 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_176
timestamp 1604681595
transform 1 0 17296 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_177
timestamp 1604681595
transform 1 0 17388 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17572 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1604681595
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_188
timestamp 1604681595
transform 1 0 18400 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_190
timestamp 1604681595
transform 1 0 18584 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18768 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18584 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_192
timestamp 1604681595
transform 1 0 18768 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_194
timestamp 1604681595
transform 1 0 18952 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1604681595
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21068 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20700 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_206
timestamp 1604681595
transform 1 0 20056 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_215
timestamp 1604681595
transform 1 0 20884 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_204
timestamp 1604681595
transform 1 0 19872 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_212
timestamp 1604681595
transform 1 0 20608 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_215
timestamp 1604681595
transform 1 0 20884 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_219
timestamp 1604681595
transform 1 0 21252 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_227
timestamp 1604681595
transform 1 0 21988 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_223
timestamp 1604681595
transform 1 0 21620 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_219
timestamp 1604681595
transform 1 0 21252 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21804 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21436 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_53_238
timestamp 1604681595
transform 1 0 23000 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_230
timestamp 1604681595
transform 1 0 22264 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 22540 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_237
timestamp 1604681595
transform 1 0 22908 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_245
timestamp 1604681595
transform 1 0 23644 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_243
timestamp 1604681595
transform 1 0 23460 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_249
timestamp 1604681595
transform 1 0 24012 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 23276 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24012 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1604681595
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_251
timestamp 1604681595
transform 1 0 24196 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 24196 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 24380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 24564 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24380 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_260
timestamp 1604681595
transform 1 0 25024 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_262
timestamp 1604681595
transform 1 0 25208 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 25208 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_272
timestamp 1604681595
transform 1 0 26128 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_268
timestamp 1604681595
transform 1 0 25760 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1604681595
transform 1 0 25392 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_266
timestamp 1604681595
transform 1 0 25576 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 25392 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25576 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_275
timestamp 1604681595
transform 1 0 26404 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_280
timestamp 1604681595
transform 1 0 26864 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_274
timestamp 1604681595
transform 1 0 26312 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 27048 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 26220 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 26588 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1604681595
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 26496 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 26772 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1604681595
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 27416 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_284
timestamp 1604681595
transform 1 0 27232 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_288
timestamp 1604681595
transform 1 0 27600 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_300
timestamp 1604681595
transform 1 0 28704 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_295
timestamp 1604681595
transform 1 0 28244 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_303
timestamp 1604681595
transform 1 0 28980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_312
timestamp 1604681595
transform 1 0 29808 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_324
timestamp 1604681595
transform 1 0 30912 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_306
timestamp 1604681595
transform 1 0 29256 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_318
timestamp 1604681595
transform 1 0 30360 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1604681595
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 32384 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_337
timestamp 1604681595
transform 1 0 32108 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_342
timestamp 1604681595
transform 1 0 32568 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_330
timestamp 1604681595
transform 1 0 31464 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_342
timestamp 1604681595
transform 1 0 32568 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1604681595
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_354
timestamp 1604681595
transform 1 0 33672 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_366
timestamp 1604681595
transform 1 0 34776 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_354
timestamp 1604681595
transform 1 0 33672 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_367
timestamp 1604681595
transform 1 0 34868 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 35420 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 35420 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_372
timestamp 1604681595
transform 1 0 35328 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1604681595
transform 1 0 35788 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_389
timestamp 1604681595
transform 1 0 36892 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_375
timestamp 1604681595
transform 1 0 35604 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_387
timestamp 1604681595
transform 1 0 36708 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604681595
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604681595
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1604681595
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_398
timestamp 1604681595
transform 1 0 37720 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1604681595
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_399
timestamp 1604681595
transform 1 0 37812 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 1380 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604681595
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_19
timestamp 1604681595
transform 1 0 2852 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 4048 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1604681595
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 3220 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_25
timestamp 1604681595
transform 1 0 3404 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1604681595
transform 1 0 3772 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_41
timestamp 1604681595
transform 1 0 4876 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 5612 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6440 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_46
timestamp 1604681595
transform 1 0 5336 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_53
timestamp 1604681595
transform 1 0 5980 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_57
timestamp 1604681595
transform 1 0 6348 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_60
timestamp 1604681595
transform 1 0 6624 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_64
timestamp 1604681595
transform 1 0 6992 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 8464 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7176 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 9016 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7544 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_68
timestamp 1604681595
transform 1 0 7360 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_72
timestamp 1604681595
transform 1 0 7728 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_84
timestamp 1604681595
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1604681595
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_88
timestamp 1604681595
transform 1 0 9200 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1604681595
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_105
timestamp 1604681595
transform 1 0 10764 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_123
timestamp 1604681595
transform 1 0 12420 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14352 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_135
timestamp 1604681595
transform 1 0 13524 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_138
timestamp 1604681595
transform 1 0 13800 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_146
timestamp 1604681595
transform 1 0 14536 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_150
timestamp 1604681595
transform 1 0 14904 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604681595
transform 1 0 15272 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1604681595
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 15732 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16100 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_157
timestamp 1604681595
transform 1 0 15548 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_161
timestamp 1604681595
transform 1 0 15916 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1604681595
transform 1 0 16284 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18768 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_177
timestamp 1604681595
transform 1 0 17388 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_190
timestamp 1604681595
transform 1 0 18584 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_194
timestamp 1604681595
transform 1 0 18952 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21068 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1604681595
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_206
timestamp 1604681595
transform 1 0 20056 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_215
timestamp 1604681595
transform 1 0 20884 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23092 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_233
timestamp 1604681595
transform 1 0 22540 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 23276 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 24656 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24196 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_245
timestamp 1604681595
transform 1 0 23644 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_249
timestamp 1604681595
transform 1 0 24012 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_253
timestamp 1604681595
transform 1 0 24380 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 27048 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1604681595
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 26772 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 25852 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_267
timestamp 1604681595
transform 1 0 25668 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_271
timestamp 1604681595
transform 1 0 26036 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_276
timestamp 1604681595
transform 1 0 26496 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_281
timestamp 1604681595
transform 1 0 26956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_298
timestamp 1604681595
transform 1 0 28520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_310
timestamp 1604681595
transform 1 0 29624 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_322
timestamp 1604681595
transform 1 0 30728 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1604681595
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_334
timestamp 1604681595
transform 1 0 31832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_337
timestamp 1604681595
transform 1 0 32108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1604681595
transform 1 0 33212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_361
timestamp 1604681595
transform 1 0 34316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 35420 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1604681595
transform 1 0 35788 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_389
timestamp 1604681595
transform 1 0 36892 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604681595
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1604681595
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_398
timestamp 1604681595
transform 1 0 37720 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1604681595
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 1840 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604681595
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 1656 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp 1604681595
transform 1 0 1380 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4048 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 3864 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 3496 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_24
timestamp 1604681595
transform 1 0 3312 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_28
timestamp 1604681595
transform 1 0 3680 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_41
timestamp 1604681595
transform 1 0 4876 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 5612 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1604681595
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 5428 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_45
timestamp 1604681595
transform 1 0 5244 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_53
timestamp 1604681595
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1604681595
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_71
timestamp 1604681595
transform 1 0 7636 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_75
timestamp 1604681595
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 9660 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_88
timestamp 1604681595
transform 1 0 9200 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_92
timestamp 1604681595
transform 1 0 9568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_95
timestamp 1604681595
transform 1 0 9844 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_107
timestamp 1604681595
transform 1 0 10948 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1604681595
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12604 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_115
timestamp 1604681595
transform 1 0 11684 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_119
timestamp 1604681595
transform 1 0 12052 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_123
timestamp 1604681595
transform 1 0 12420 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_127
timestamp 1604681595
transform 1 0 12788 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_131
timestamp 1604681595
transform 1 0 13156 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_134
timestamp 1604681595
transform 1 0 13432 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_138
timestamp 1604681595
transform 1 0 13800 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_153
timestamp 1604681595
transform 1 0 15180 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 15364 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_157
timestamp 1604681595
transform 1 0 15548 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 15732 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_161
timestamp 1604681595
transform 1 0 15916 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_prog_clk
timestamp 1604681595
transform 1 0 16192 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_167
timestamp 1604681595
transform 1 0 16468 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_171
timestamp 1604681595
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 16652 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604681595
transform 1 0 16928 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1604681595
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_175
timestamp 1604681595
transform 1 0 17204 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_179
timestamp 1604681595
transform 1 0 17572 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 21068 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 20884 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 20516 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19688 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 20148 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_200
timestamp 1604681595
transform 1 0 19504 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_204
timestamp 1604681595
transform 1 0 19872 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_209
timestamp 1604681595
transform 1 0 20332 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_213
timestamp 1604681595
transform 1 0 20700 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23092 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22724 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_233
timestamp 1604681595
transform 1 0 22540 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_237
timestamp 1604681595
transform 1 0 22908 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 25208 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1604681595
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 25024 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 24656 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_241
timestamp 1604681595
transform 1 0 23276 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_254
timestamp 1604681595
transform 1 0 24472 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_258
timestamp 1604681595
transform 1 0 24840 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 26772 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 26588 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26220 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_271
timestamp 1604681595
transform 1 0 26036 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_275
timestamp 1604681595
transform 1 0 26404 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1604681595
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 27784 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 28152 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 28520 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_288
timestamp 1604681595
transform 1 0 27600 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_292
timestamp 1604681595
transform 1 0 27968 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_296
timestamp 1604681595
transform 1 0 28336 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_300
timestamp 1604681595
transform 1 0 28704 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_304
timestamp 1604681595
transform 1 0 29072 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 29440 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_306
timestamp 1604681595
transform 1 0 29256 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_310
timestamp 1604681595
transform 1 0 29624 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1604681595
transform 1 0 30728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_334
timestamp 1604681595
transform 1 0 31832 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_346
timestamp 1604681595
transform 1 0 32936 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1604681595
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_358
timestamp 1604681595
transform 1 0 34040 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1604681595
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1604681595
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_391
timestamp 1604681595
transform 1 0 37076 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604681595
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1604681595
transform 1 0 38180 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 1748 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604681595
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 1564 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1604681595
transform 1 0 1380 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 4048 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1604681595
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 3772 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3404 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_23
timestamp 1604681595
transform 1 0 3220 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1604681595
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6532 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 6348 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_48
timestamp 1604681595
transform 1 0 5520 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_52
timestamp 1604681595
transform 1 0 5888 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_55
timestamp 1604681595
transform 1 0 6164 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 8464 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 7544 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_68
timestamp 1604681595
transform 1 0 7360 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_72
timestamp 1604681595
transform 1 0 7728 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_84
timestamp 1604681595
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_88
timestamp 1604681595
transform 1 0 9200 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1604681595
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_97
timestamp 1604681595
transform 1 0 10028 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 9660 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_101
timestamp 1604681595
transform 1 0 10396 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_107
timestamp 1604681595
transform 1 0 10948 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11868 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12880 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_111
timestamp 1604681595
transform 1 0 11316 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_126
timestamp 1604681595
transform 1 0 12696 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_130
timestamp 1604681595
transform 1 0 13064 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 14996 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14628 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_145
timestamp 1604681595
transform 1 0 14444 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_149
timestamp 1604681595
transform 1 0 14812 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 33184
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1604681595
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17940 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17756 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_175
timestamp 1604681595
transform 1 0 17204 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 20884 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1604681595
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_199
timestamp 1604681595
transform 1 0 19412 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_211
timestamp 1604681595
transform 1 0 20516 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23092 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_231
timestamp 1604681595
transform 1 0 22356 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24840 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24656 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_248
timestamp 1604681595
transform 1 0 23920 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_252
timestamp 1604681595
transform 1 0 24288 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 27140 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1604681595
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 26956 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_267
timestamp 1604681595
transform 1 0 25668 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_276
timestamp 1604681595
transform 1 0 26496 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_280
timestamp 1604681595
transform 1 0 26864 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_299
timestamp 1604681595
transform 1 0 28612 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 29348 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_311
timestamp 1604681595
transform 1 0 29716 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_323
timestamp 1604681595
transform 1 0 30820 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1604681595
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_335
timestamp 1604681595
transform 1 0 31924 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_337
timestamp 1604681595
transform 1 0 32108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_349
timestamp 1604681595
transform 1 0 33212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_361
timestamp 1604681595
transform 1 0 34316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_373
timestamp 1604681595
transform 1 0 35420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1604681595
transform 1 0 36524 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604681595
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1604681595
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_398
timestamp 1604681595
transform 1 0 37720 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1604681595
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 2852 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604681595
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 2668 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 2300 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 1748 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1604681595
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_9
timestamp 1604681595
transform 1 0 1932 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_15
timestamp 1604681595
transform 1 0 2484 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 4416 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1604681595
transform 1 0 4232 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 3864 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_28
timestamp 1604681595
transform 1 0 3680 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_32
timestamp 1604681595
transform 1 0 4048 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 6808 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1604681595
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 6072 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1604681595
transform 1 0 6440 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_52
timestamp 1604681595
transform 1 0 5888 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_56
timestamp 1604681595
transform 1 0 6256 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_60
timestamp 1604681595
transform 1 0 6624 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8372 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_71
timestamp 1604681595
transform 1 0 7636 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_75
timestamp 1604681595
transform 1 0 8004 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10212 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_97
timestamp 1604681595
transform 1 0 10028 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_101
timestamp 1604681595
transform 1 0 10396 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1604681595
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_114
timestamp 1604681595
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_118
timestamp 1604681595
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604681595
transform 1 0 14168 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 14996 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 14628 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13984 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_132
timestamp 1604681595
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_136
timestamp 1604681595
transform 1 0 13616 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_145
timestamp 1604681595
transform 1 0 14444 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_149
timestamp 1604681595
transform 1 0 14812 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 15180 0 1 33184
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_57_174
timestamp 1604681595
transform 1 0 17112 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1604681595
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_179
timestamp 1604681595
transform 1 0 17572 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1604681595
transform 1 0 20608 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
timestamp 1604681595
transform 1 0 20424 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
timestamp 1604681595
transform 1 0 20056 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19688 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_200
timestamp 1604681595
transform 1 0 19504 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_204
timestamp 1604681595
transform 1 0 19872 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_208
timestamp 1604681595
transform 1 0 20240 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
timestamp 1604681595
transform 1 0 22264 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
timestamp 1604681595
transform 1 0 22632 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_228
timestamp 1604681595
transform 1 0 22080 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_232
timestamp 1604681595
transform 1 0 22448 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_236
timestamp 1604681595
transform 1 0 22816 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_240
timestamp 1604681595
transform 1 0 23184 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1604681595
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
timestamp 1604681595
transform 1 0 23368 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 25208 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_254
timestamp 1604681595
transform 1 0 24472 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_258
timestamp 1604681595
transform 1 0 24840 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 25392 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1604681595
transform 1 0 26956 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
timestamp 1604681595
transform 1 0 26772 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
timestamp 1604681595
transform 1 0 26404 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_273
timestamp 1604681595
transform 1 0 26220 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_277
timestamp 1604681595
transform 1 0 26588 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1604681595
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 28612 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_297
timestamp 1604681595
transform 1 0 28428 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_301
timestamp 1604681595
transform 1 0 28796 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_306
timestamp 1604681595
transform 1 0 29256 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_318
timestamp 1604681595
transform 1 0 30360 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_330
timestamp 1604681595
transform 1 0 31464 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_342
timestamp 1604681595
transform 1 0 32568 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1604681595
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 35236 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_354
timestamp 1604681595
transform 1 0 33672 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_367
timestamp 1604681595
transform 1 0 34868 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 35420 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 35972 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_377
timestamp 1604681595
transform 1 0 35788 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_381
timestamp 1604681595
transform 1 0 36156 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1604681595
transform 1 0 37260 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604681595
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1604681595
transform 1 0 38364 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604681595
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 1564 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 2852 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1604681595
transform 1 0 1380 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1604681595
transform 1 0 1748 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_21
timestamp 1604681595
transform 1 0 3036 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 4508 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1604681595
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 4324 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_32
timestamp 1604681595
transform 1 0 4048 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1604681595
transform 1 0 6072 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5520 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5888 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_46
timestamp 1604681595
transform 1 0 5336 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_50
timestamp 1604681595
transform 1 0 5704 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 8464 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 9016 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_70
timestamp 1604681595
transform 1 0 7544 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_78
timestamp 1604681595
transform 1 0 8280 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_84
timestamp 1604681595
transform 1 0 8832 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1604681595
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_88
timestamp 1604681595
transform 1 0 9200 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_109
timestamp 1604681595
transform 1 0 11132 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11868 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_115
timestamp 1604681595
transform 1 0 11684 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604681595
transform 1 0 14076 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14720 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1604681595
transform 1 0 13340 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_144
timestamp 1604681595
transform 1 0 14352 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_150
timestamp 1604681595
transform 1 0 14904 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1604681595
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16928 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_170
timestamp 1604681595
transform 1 0 16744 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_174
timestamp 1604681595
transform 1 0 17112 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17756 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17296 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_178
timestamp 1604681595
transform 1 0 17480 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1604681595
transform 1 0 20884 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1604681595
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19596 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19964 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_197
timestamp 1604681595
transform 1 0 19228 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_203
timestamp 1604681595
transform 1 0 19780 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_207
timestamp 1604681595
transform 1 0 20148 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_213
timestamp 1604681595
transform 1 0 20700 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
timestamp 1604681595
transform 1 0 22540 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_231
timestamp 1604681595
transform 1 0 22356 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_235
timestamp 1604681595
transform 1 0 22724 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1604681595
transform 1 0 23644 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23460 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_261
timestamp 1604681595
transform 1 0 25116 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1604681595
transform 1 0 26864 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1604681595
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 25392 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 25760 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
timestamp 1604681595
transform 1 0 26680 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_266
timestamp 1604681595
transform 1 0 25576 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_270
timestamp 1604681595
transform 1 0 25944 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_274
timestamp 1604681595
transform 1 0 26312 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_276
timestamp 1604681595
transform 1 0 26496 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_296
timestamp 1604681595
transform 1 0 28336 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_308
timestamp 1604681595
transform 1 0 29440 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_320
timestamp 1604681595
transform 1 0 30544 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1604681595
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_332
timestamp 1604681595
transform 1 0 31648 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_337
timestamp 1604681595
transform 1 0 32108 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1604681595
transform 1 0 33212 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_361
timestamp 1604681595
transform 1 0 34316 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 35420 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1604681595
transform 1 0 35788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_389
timestamp 1604681595
transform 1 0 36892 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604681595
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1604681595
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_398
timestamp 1604681595
transform 1 0 37720 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1604681595
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_7
timestamp 1604681595
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604681595
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604681595
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_19
timestamp 1604681595
transform 1 0 2852 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_11
timestamp 1604681595
transform 1 0 2116 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 3036 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 2484 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_19
timestamp 1604681595
transform 1 0 2852 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1604681595
transform 1 0 1748 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_23
timestamp 1604681595
transform 1 0 3220 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 3588 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_37
timestamp 1604681595
transform 1 0 4508 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_32
timestamp 1604681595
transform 1 0 4048 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_39
timestamp 1604681595
transform 1 0 4692 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_35
timestamp 1604681595
transform 1 0 4324 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_31
timestamp 1604681595
transform 1 0 3956 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 4508 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 4140 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1604681595
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 4140 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
timestamp 1604681595
transform 1 0 4968 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_53
timestamp 1604681595
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_61
timestamp 1604681595
transform 1 0 6716 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_62
timestamp 1604681595
transform 1 0 6808 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1604681595
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
timestamp 1604681595
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 7084 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1604681595
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1604681595
transform 1 0 5244 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_60_71
timestamp 1604681595
transform 1 0 7636 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_67
timestamp 1604681595
transform 1 0 7268 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
timestamp 1604681595
transform 1 0 7452 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1604681595
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_82
timestamp 1604681595
transform 1 0 8648 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_77
timestamp 1604681595
transform 1 0 8188 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_84
timestamp 1604681595
transform 1 0 8832 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 9016 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 8280 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1604681595
transform 1 0 7360 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_60_90
timestamp 1604681595
transform 1 0 9384 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_88
timestamp 1604681595
transform 1 0 9200 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 9384 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1604681595
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9568 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_60_102
timestamp 1604681595
transform 1 0 10488 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_98
timestamp 1604681595
transform 1 0 10120 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_105
timestamp 1604681595
transform 1 0 10764 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_101
timestamp 1604681595
transform 1 0 10396 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 10580 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604681595
transform 1 0 11132 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_110
timestamp 1604681595
transform 1 0 11224 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_116
timestamp 1604681595
transform 1 0 11776 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_112
timestamp 1604681595
transform 1 0 11408 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_129
timestamp 1604681595
transform 1 0 12972 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_123
timestamp 1604681595
transform 1 0 12420 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1604681595
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12512 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_60_141
timestamp 1604681595
transform 1 0 14076 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_133
timestamp 1604681595
transform 1 0 13340 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_140
timestamp 1604681595
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 13708 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_150
timestamp 1604681595
transform 1 0 14904 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_147
timestamp 1604681595
transform 1 0 14628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_144
timestamp 1604681595
transform 1 0 14352 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 14168 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14720 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604681595
transform 1 0 16928 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1604681595
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_164
timestamp 1604681595
transform 1 0 16192 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_168
timestamp 1604681595
transform 1 0 16560 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_163
timestamp 1604681595
transform 1 0 16100 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_180
timestamp 1604681595
transform 1 0 17664 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_179
timestamp 1604681595
transform 1 0 17572 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_175
timestamp 1604681595
transform 1 0 17204 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1604681595
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_60_192
timestamp 1604681595
transform 1 0 18768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_186
timestamp 1604681595
transform 1 0 18216 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_193
timestamp 1604681595
transform 1 0 18860 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 18400 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 19044 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_203
timestamp 1604681595
transform 1 0 19780 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_200
timestamp 1604681595
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_197
timestamp 1604681595
transform 1 0 19228 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19596 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_60_215
timestamp 1604681595
transform 1 0 20884 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_211
timestamp 1604681595
transform 1 0 20516 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_214
timestamp 1604681595
transform 1 0 20792 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_210
timestamp 1604681595
transform 1 0 20424 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
timestamp 1604681595
transform 1 0 20608 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 20976 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1604681595
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 20976 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1604681595
transform 1 0 21160 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1604681595
transform 1 0 22080 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
timestamp 1604681595
transform 1 0 22816 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
timestamp 1604681595
transform 1 0 21528 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_234
timestamp 1604681595
transform 1 0 22632 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_238
timestamp 1604681595
transform 1 0 23000 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_220
timestamp 1604681595
transform 1 0 21344 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1604681595
transform 1 0 21712 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1604681595
transform 1 0 24104 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_244
timestamp 1604681595
transform 1 0 23552 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_249
timestamp 1604681595
transform 1 0 24012 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_245
timestamp 1604681595
transform 1 0 23644 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
timestamp 1604681595
transform 1 0 23920 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 23828 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
timestamp 1604681595
transform 1 0 24196 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1604681595
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_254
timestamp 1604681595
transform 1 0 24472 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24288 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 24656 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24840 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1604681595
transform 1 0 24380 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1604681595
transform 1 0 26496 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1604681595
transform 1 0 26588 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1604681595
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1604681595
transform 1 0 26404 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
timestamp 1604681595
transform 1 0 26036 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_269
timestamp 1604681595
transform 1 0 25852 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_273
timestamp 1604681595
transform 1 0 26220 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_267
timestamp 1604681595
transform 1 0 25668 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1604681595
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
timestamp 1604681595
transform 1 0 28244 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_293
timestamp 1604681595
transform 1 0 28060 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_297
timestamp 1604681595
transform 1 0 28428 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_292
timestamp 1604681595
transform 1 0 27968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_304
timestamp 1604681595
transform 1 0 29072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_306
timestamp 1604681595
transform 1 0 29256 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_318
timestamp 1604681595
transform 1 0 30360 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_316
timestamp 1604681595
transform 1 0 30176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1604681595
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_330
timestamp 1604681595
transform 1 0 31464 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_342
timestamp 1604681595
transform 1 0 32568 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_328
timestamp 1604681595
transform 1 0 31280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_337
timestamp 1604681595
transform 1 0 32108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_349
timestamp 1604681595
transform 1 0 33212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1604681595
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 35236 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_354
timestamp 1604681595
transform 1 0 33672 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1604681595
transform 1 0 34868 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_361
timestamp 1604681595
transform 1 0 34316 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_369
timestamp 1604681595
transform 1 0 35052 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_381
timestamp 1604681595
transform 1 0 36156 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_377
timestamp 1604681595
transform 1 0 35788 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 35972 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 35420 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 35328 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_388
timestamp 1604681595
transform 1 0 36800 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_389
timestamp 1604681595
transform 1 0 36892 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 37076 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 36524 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_376
timestamp 1604681595
transform 1 0 35696 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1604681595
transform 1 0 37260 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604681595
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604681595
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1604681595
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1604681595
transform 1 0 38364 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_396
timestamp 1604681595
transform 1 0 37536 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1604681595
transform 1 0 37720 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1604681595
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604681595
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604681595
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604681595
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1604681595
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_39
timestamp 1604681595
transform 1 0 4692 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 5428 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 7084 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1604681595
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 5980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_51
timestamp 1604681595
transform 1 0 5796 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_55
timestamp 1604681595
transform 1 0 6164 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_61_62
timestamp 1604681595
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 8188 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 7636 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 8740 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_69
timestamp 1604681595
transform 1 0 7452 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_73
timestamp 1604681595
transform 1 0 7820 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_81
timestamp 1604681595
transform 1 0 8556 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_85
timestamp 1604681595
transform 1 0 8924 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_97
timestamp 1604681595
transform 1 0 10028 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_109
timestamp 1604681595
transform 1 0 11132 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604681595
transform 1 0 12420 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1604681595
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_121
timestamp 1604681595
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_126
timestamp 1604681595
transform 1 0 12696 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13892 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13708 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_134
timestamp 1604681595
transform 1 0 13432 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16284 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_155
timestamp 1604681595
transform 1 0 15364 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_159
timestamp 1604681595
transform 1 0 15732 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_163
timestamp 1604681595
transform 1 0 16100 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_167
timestamp 1604681595
transform 1 0 16468 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1604681595
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_179
timestamp 1604681595
transform 1 0 17572 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1604681595
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1604681595
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21160 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20792 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_208
timestamp 1604681595
transform 1 0 20240 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_216
timestamp 1604681595
transform 1 0 20976 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21344 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 22356 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 22724 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 23092 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_229
timestamp 1604681595
transform 1 0 22172 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_233
timestamp 1604681595
transform 1 0 22540 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_237
timestamp 1604681595
transform 1 0 22908 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 24932 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 23644 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1604681595
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 24196 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 24564 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_241
timestamp 1604681595
transform 1 0 23276 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_249
timestamp 1604681595
transform 1 0 24012 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_253
timestamp 1604681595
transform 1 0 24380 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_257
timestamp 1604681595
transform 1 0 24748 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 26312 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 26128 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 25760 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_263
timestamp 1604681595
transform 1 0 25300 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_267
timestamp 1604681595
transform 1 0 25668 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_270
timestamp 1604681595
transform 1 0 25944 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_283
timestamp 1604681595
transform 1 0 27140 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1604681595
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_295
timestamp 1604681595
transform 1 0 28244 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_303
timestamp 1604681595
transform 1 0 28980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_306
timestamp 1604681595
transform 1 0 29256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1604681595
transform 1 0 30360 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_330
timestamp 1604681595
transform 1 0 31464 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_342
timestamp 1604681595
transform 1 0 32568 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1604681595
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_354
timestamp 1604681595
transform 1 0 33672 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_367
timestamp 1604681595
transform 1 0 34868 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 35420 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 35972 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_377
timestamp 1604681595
transform 1 0 35788 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_381
timestamp 1604681595
transform 1 0 36156 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1604681595
transform 1 0 37260 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604681595
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1604681595
transform 1 0 38364 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604681595
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604681595
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604681595
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1604681595
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604681595
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1604681595
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 6808 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1604681595
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_56
timestamp 1604681595
transform 1 0 6256 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_66
timestamp 1604681595
transform 1 0 7176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_78
timestamp 1604681595
transform 1 0 8280 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1604681595
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_90
timestamp 1604681595
transform 1 0 9384 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604681595
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604681595
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604681595
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_129
timestamp 1604681595
transform 1 0 12972 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_137
timestamp 1604681595
transform 1 0 13708 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1604681595
transform 1 0 14076 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1604681595
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_163
timestamp 1604681595
transform 1 0 16100 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_175
timestamp 1604681595
transform 1 0 17204 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_187
timestamp 1604681595
transform 1 0 18308 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1604681595
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_199
timestamp 1604681595
transform 1 0 19412 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_211
timestamp 1604681595
transform 1 0 20516 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_215
timestamp 1604681595
transform 1 0 20884 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 22264 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21344 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_219
timestamp 1604681595
transform 1 0 21252 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_222
timestamp 1604681595
transform 1 0 21528 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_239
timestamp 1604681595
transform 1 0 23092 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 23828 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 24932 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_251
timestamp 1604681595
transform 1 0 24196 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_261
timestamp 1604681595
transform 1 0 25116 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1604681595
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 26680 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_273
timestamp 1604681595
transform 1 0 26220 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_276
timestamp 1604681595
transform 1 0 26496 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_280
timestamp 1604681595
transform 1 0 26864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_292
timestamp 1604681595
transform 1 0 27968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_304
timestamp 1604681595
transform 1 0 29072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_316
timestamp 1604681595
transform 1 0 30176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1604681595
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_328
timestamp 1604681595
transform 1 0 31280 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1604681595
transform 1 0 32108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1604681595
transform 1 0 33212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_361
timestamp 1604681595
transform 1 0 34316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_373
timestamp 1604681595
transform 1 0 35420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_385
timestamp 1604681595
transform 1 0 36524 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604681595
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1604681595
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_398
timestamp 1604681595
transform 1 0 37720 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1604681595
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604681595
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604681595
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604681595
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604681595
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604681595
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 6808 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1604681595
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604681595
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604681595
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 7360 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_66
timestamp 1604681595
transform 1 0 7176 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_70
timestamp 1604681595
transform 1 0 7544 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_82
timestamp 1604681595
transform 1 0 8648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1604681595
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_106
timestamp 1604681595
transform 1 0 10856 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1604681595
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1604681595
transform 1 0 11960 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604681595
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_135
timestamp 1604681595
transform 1 0 13524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_147
timestamp 1604681595
transform 1 0 14628 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_159
timestamp 1604681595
transform 1 0 15732 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_171
timestamp 1604681595
transform 1 0 16836 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1604681595
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1604681595
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1604681595
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1604681595
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_220
timestamp 1604681595
transform 1 0 21344 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_232
timestamp 1604681595
transform 1 0 22448 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1604681595
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1604681595
transform 1 0 23644 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_257
timestamp 1604681595
transform 1 0 24748 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_269
timestamp 1604681595
transform 1 0 25852 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1604681595
transform 1 0 26956 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1604681595
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1604681595
transform 1 0 28060 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1604681595
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1604681595
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_330
timestamp 1604681595
transform 1 0 31464 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_342
timestamp 1604681595
transform 1 0 32568 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1604681595
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_354
timestamp 1604681595
transform 1 0 33672 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1604681595
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1604681595
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1604681595
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604681595
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1604681595
transform 1 0 38180 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604681595
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604681595
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604681595
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1604681595
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604681595
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604681595
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1604681595
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604681595
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604681595
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604681595
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604681595
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604681595
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1604681595
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604681595
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604681595
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1604681595
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604681595
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604681595
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_137
timestamp 1604681595
transform 1 0 13708 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_149
timestamp 1604681595
transform 1 0 14812 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1604681595
transform 1 0 15364 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_156
timestamp 1604681595
transform 1 0 15456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_168
timestamp 1604681595
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1604681595
transform 1 0 18216 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_180
timestamp 1604681595
transform 1 0 17664 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_187
timestamp 1604681595
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1604681595
transform 1 0 21068 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_199
timestamp 1604681595
transform 1 0 19412 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_211
timestamp 1604681595
transform 1 0 20516 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_218
timestamp 1604681595
transform 1 0 21160 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_230
timestamp 1604681595
transform 1 0 22264 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1604681595
transform 1 0 23920 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_242
timestamp 1604681595
transform 1 0 23368 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_249
timestamp 1604681595
transform 1 0 24012 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_261
timestamp 1604681595
transform 1 0 25116 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1604681595
transform 1 0 26772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1604681595
transform 1 0 26220 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_280
timestamp 1604681595
transform 1 0 26864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_292
timestamp 1604681595
transform 1 0 27968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_304
timestamp 1604681595
transform 1 0 29072 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1604681595
transform 1 0 29624 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_311
timestamp 1604681595
transform 1 0 29716 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_323
timestamp 1604681595
transform 1 0 30820 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1604681595
transform 1 0 32476 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_335
timestamp 1604681595
transform 1 0 31924 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_342
timestamp 1604681595
transform 1 0 32568 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_354
timestamp 1604681595
transform 1 0 33672 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_366
timestamp 1604681595
transform 1 0 34776 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1604681595
transform 1 0 35328 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_373
timestamp 1604681595
transform 1 0 35420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_385
timestamp 1604681595
transform 1 0 36524 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604681595
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1604681595
transform 1 0 38180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_397
timestamp 1604681595
transform 1 0 37628 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_404
timestamp 1604681595
transform 1 0 38272 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal2 s 30010 0 30066 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 38290 39520 38346 40000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 36634 0 36690 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 39394 39520 39450 40000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 Test_en
port 4 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_width_0_height_0__pin_50_
port 5 nsew default tristate
rlabel metal2 s 9954 0 10010 480 6 bottom_width_0_height_0__pin_51_
port 6 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 ccff_head
port 7 nsew default input
rlabel metal3 s 39520 10208 40000 10328 6 ccff_tail
port 8 nsew default tristate
rlabel metal2 s 23294 0 23350 480 6 clk
port 9 nsew default input
rlabel metal3 s 0 33328 480 33448 6 left_width_0_height_0__pin_52_
port 10 nsew default input
rlabel metal3 s 0 6672 480 6792 6 prog_clk
port 11 nsew default input
rlabel metal3 s 39520 11432 40000 11552 6 right_width_0_height_0__pin_16_
port 12 nsew default input
rlabel metal3 s 39520 12656 40000 12776 6 right_width_0_height_0__pin_17_
port 13 nsew default input
rlabel metal3 s 39520 13880 40000 14000 6 right_width_0_height_0__pin_18_
port 14 nsew default input
rlabel metal3 s 39520 14968 40000 15088 6 right_width_0_height_0__pin_19_
port 15 nsew default input
rlabel metal3 s 39520 16192 40000 16312 6 right_width_0_height_0__pin_20_
port 16 nsew default input
rlabel metal3 s 39520 17416 40000 17536 6 right_width_0_height_0__pin_21_
port 17 nsew default input
rlabel metal3 s 39520 18640 40000 18760 6 right_width_0_height_0__pin_22_
port 18 nsew default input
rlabel metal3 s 39520 19864 40000 19984 6 right_width_0_height_0__pin_23_
port 19 nsew default input
rlabel metal3 s 39520 21088 40000 21208 6 right_width_0_height_0__pin_24_
port 20 nsew default input
rlabel metal3 s 39520 22312 40000 22432 6 right_width_0_height_0__pin_25_
port 21 nsew default input
rlabel metal3 s 39520 23536 40000 23656 6 right_width_0_height_0__pin_26_
port 22 nsew default input
rlabel metal3 s 39520 24760 40000 24880 6 right_width_0_height_0__pin_27_
port 23 nsew default input
rlabel metal3 s 39520 25984 40000 26104 6 right_width_0_height_0__pin_28_
port 24 nsew default input
rlabel metal3 s 39520 27208 40000 27328 6 right_width_0_height_0__pin_29_
port 25 nsew default input
rlabel metal3 s 39520 28296 40000 28416 6 right_width_0_height_0__pin_30_
port 26 nsew default input
rlabel metal3 s 39520 29520 40000 29640 6 right_width_0_height_0__pin_31_
port 27 nsew default input
rlabel metal3 s 39520 552 40000 672 6 right_width_0_height_0__pin_42_lower
port 28 nsew default tristate
rlabel metal3 s 39520 30744 40000 30864 6 right_width_0_height_0__pin_42_upper
port 29 nsew default tristate
rlabel metal3 s 39520 1640 40000 1760 6 right_width_0_height_0__pin_43_lower
port 30 nsew default tristate
rlabel metal3 s 39520 31968 40000 32088 6 right_width_0_height_0__pin_43_upper
port 31 nsew default tristate
rlabel metal3 s 39520 2864 40000 2984 6 right_width_0_height_0__pin_44_lower
port 32 nsew default tristate
rlabel metal3 s 39520 33192 40000 33312 6 right_width_0_height_0__pin_44_upper
port 33 nsew default tristate
rlabel metal3 s 39520 4088 40000 4208 6 right_width_0_height_0__pin_45_lower
port 34 nsew default tristate
rlabel metal3 s 39520 34416 40000 34536 6 right_width_0_height_0__pin_45_upper
port 35 nsew default tristate
rlabel metal3 s 39520 5312 40000 5432 6 right_width_0_height_0__pin_46_lower
port 36 nsew default tristate
rlabel metal3 s 39520 35640 40000 35760 6 right_width_0_height_0__pin_46_upper
port 37 nsew default tristate
rlabel metal3 s 39520 6536 40000 6656 6 right_width_0_height_0__pin_47_lower
port 38 nsew default tristate
rlabel metal3 s 39520 36864 40000 36984 6 right_width_0_height_0__pin_47_upper
port 39 nsew default tristate
rlabel metal3 s 39520 7760 40000 7880 6 right_width_0_height_0__pin_48_lower
port 40 nsew default tristate
rlabel metal3 s 39520 38088 40000 38208 6 right_width_0_height_0__pin_48_upper
port 41 nsew default tristate
rlabel metal3 s 39520 8984 40000 9104 6 right_width_0_height_0__pin_49_lower
port 42 nsew default tristate
rlabel metal3 s 39520 39312 40000 39432 6 right_width_0_height_0__pin_49_upper
port 43 nsew default tristate
rlabel metal2 s 9402 39520 9458 40000 6 top_width_0_height_0__pin_0_
port 44 nsew default input
rlabel metal2 s 20534 39520 20590 40000 6 top_width_0_height_0__pin_10_
port 45 nsew default input
rlabel metal2 s 21638 39520 21694 40000 6 top_width_0_height_0__pin_11_
port 46 nsew default input
rlabel metal2 s 22742 39520 22798 40000 6 top_width_0_height_0__pin_12_
port 47 nsew default input
rlabel metal2 s 23846 39520 23902 40000 6 top_width_0_height_0__pin_13_
port 48 nsew default input
rlabel metal2 s 24950 39520 25006 40000 6 top_width_0_height_0__pin_14_
port 49 nsew default input
rlabel metal2 s 26054 39520 26110 40000 6 top_width_0_height_0__pin_15_
port 50 nsew default input
rlabel metal2 s 10506 39520 10562 40000 6 top_width_0_height_0__pin_1_
port 51 nsew default input
rlabel metal2 s 11610 39520 11666 40000 6 top_width_0_height_0__pin_2_
port 52 nsew default input
rlabel metal2 s 27250 39520 27306 40000 6 top_width_0_height_0__pin_32_
port 53 nsew default input
rlabel metal2 s 28354 39520 28410 40000 6 top_width_0_height_0__pin_33_
port 54 nsew default input
rlabel metal2 s 29458 39520 29514 40000 6 top_width_0_height_0__pin_34_lower
port 55 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 top_width_0_height_0__pin_34_upper
port 56 nsew default tristate
rlabel metal2 s 30562 39520 30618 40000 6 top_width_0_height_0__pin_35_lower
port 57 nsew default tristate
rlabel metal2 s 1674 39520 1730 40000 6 top_width_0_height_0__pin_35_upper
port 58 nsew default tristate
rlabel metal2 s 31666 39520 31722 40000 6 top_width_0_height_0__pin_36_lower
port 59 nsew default tristate
rlabel metal2 s 2778 39520 2834 40000 6 top_width_0_height_0__pin_36_upper
port 60 nsew default tristate
rlabel metal2 s 32770 39520 32826 40000 6 top_width_0_height_0__pin_37_lower
port 61 nsew default tristate
rlabel metal2 s 3882 39520 3938 40000 6 top_width_0_height_0__pin_37_upper
port 62 nsew default tristate
rlabel metal2 s 33874 39520 33930 40000 6 top_width_0_height_0__pin_38_lower
port 63 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 top_width_0_height_0__pin_38_upper
port 64 nsew default tristate
rlabel metal2 s 34978 39520 35034 40000 6 top_width_0_height_0__pin_39_lower
port 65 nsew default tristate
rlabel metal2 s 6090 39520 6146 40000 6 top_width_0_height_0__pin_39_upper
port 66 nsew default tristate
rlabel metal2 s 12714 39520 12770 40000 6 top_width_0_height_0__pin_3_
port 67 nsew default input
rlabel metal2 s 36082 39520 36138 40000 6 top_width_0_height_0__pin_40_lower
port 68 nsew default tristate
rlabel metal2 s 7194 39520 7250 40000 6 top_width_0_height_0__pin_40_upper
port 69 nsew default tristate
rlabel metal2 s 37186 39520 37242 40000 6 top_width_0_height_0__pin_41_lower
port 70 nsew default tristate
rlabel metal2 s 8298 39520 8354 40000 6 top_width_0_height_0__pin_41_upper
port 71 nsew default tristate
rlabel metal2 s 13910 39520 13966 40000 6 top_width_0_height_0__pin_4_
port 72 nsew default input
rlabel metal2 s 15014 39520 15070 40000 6 top_width_0_height_0__pin_5_
port 73 nsew default input
rlabel metal2 s 16118 39520 16174 40000 6 top_width_0_height_0__pin_6_
port 74 nsew default input
rlabel metal2 s 17222 39520 17278 40000 6 top_width_0_height_0__pin_7_
port 75 nsew default input
rlabel metal2 s 18326 39520 18382 40000 6 top_width_0_height_0__pin_8_
port 76 nsew default input
rlabel metal2 s 19430 39520 19486 40000 6 top_width_0_height_0__pin_9_
port 77 nsew default input
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 78 nsew default input
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 79 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
