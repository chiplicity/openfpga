magic
tech EFS8A
magscale 1 2
timestamp 1602209602
<< locali >>
rect 2789 4063 2823 4165
<< viali >>
rect 17969 21097 18003 21131
rect 17049 21029 17083 21063
rect 21649 21029 21683 21063
rect 16313 20961 16347 20995
rect 16773 20961 16807 20995
rect 18153 20961 18187 20995
rect 18429 20961 18463 20995
rect 20913 20961 20947 20995
rect 21465 20961 21499 20995
rect 19257 20757 19291 20791
rect 14657 20485 14691 20519
rect 20361 20485 20395 20519
rect 20729 20485 20763 20519
rect 4537 20417 4571 20451
rect 8401 20417 8435 20451
rect 11529 20417 11563 20451
rect 13185 20417 13219 20451
rect 15761 20417 15795 20451
rect 18705 20417 18739 20451
rect 19901 20417 19935 20451
rect 21649 20417 21683 20451
rect 3525 20349 3559 20383
rect 4169 20349 4203 20383
rect 4445 20349 4479 20383
rect 7757 20349 7791 20383
rect 8125 20349 8159 20383
rect 8309 20349 8343 20383
rect 10793 20349 10827 20383
rect 11253 20349 11287 20383
rect 12449 20349 12483 20383
rect 12909 20349 12943 20383
rect 15209 20349 15243 20383
rect 15669 20349 15703 20383
rect 19441 20349 19475 20383
rect 19625 20349 19659 20383
rect 20913 20349 20947 20383
rect 21465 20349 21499 20383
rect 3893 20281 3927 20315
rect 15117 20281 15151 20315
rect 16681 20281 16715 20315
rect 21925 20281 21959 20315
rect 10609 20213 10643 20247
rect 12265 20213 12299 20247
rect 16405 20213 16439 20247
rect 18337 20213 18371 20247
rect 18981 20213 19015 20247
rect 22293 20213 22327 20247
rect 5273 19941 5307 19975
rect 8769 19941 8803 19975
rect 16681 19941 16715 19975
rect 19257 19941 19291 19975
rect 21649 19941 21683 19975
rect 4813 19873 4847 19907
rect 4997 19873 5031 19907
rect 8033 19873 8067 19907
rect 8493 19873 8527 19907
rect 16221 19873 16255 19907
rect 16497 19873 16531 19907
rect 18521 19873 18555 19907
rect 18981 19873 19015 19907
rect 20913 19873 20947 19907
rect 21465 19873 21499 19907
rect 7941 19805 7975 19839
rect 10885 19669 10919 19703
rect 12449 19669 12483 19703
rect 8033 19465 8067 19499
rect 21281 19465 21315 19499
rect 21005 19397 21039 19431
rect 16405 19329 16439 19363
rect 19625 19329 19659 19363
rect 18889 19261 18923 19295
rect 19349 19261 19383 19295
rect 4629 19193 4663 19227
rect 16037 19193 16071 19227
rect 4997 19125 5031 19159
rect 8493 19125 8527 19159
rect 18521 19125 18555 19159
rect 1593 18921 1627 18955
rect 21649 18853 21683 18887
rect 1501 18785 1535 18819
rect 1961 18785 1995 18819
rect 20913 18785 20947 18819
rect 21373 18785 21407 18819
rect 18521 18717 18555 18751
rect 19257 18717 19291 18751
rect 18889 18649 18923 18683
rect 1961 18377 1995 18411
rect 20913 18173 20947 18207
rect 21373 18173 21407 18207
rect 21649 18173 21683 18207
rect 20361 18105 20395 18139
rect 20729 18105 20763 18139
rect 1685 18037 1719 18071
rect 19993 18037 20027 18071
rect 1685 17833 1719 17867
rect 21097 17493 21131 17527
rect 1593 17085 1627 17119
rect 1869 17085 1903 17119
rect 1501 16949 1535 16983
rect 19441 16745 19475 16779
rect 1685 16405 1719 16439
rect 14565 16065 14599 16099
rect 15393 16065 15427 16099
rect 20085 16065 20119 16099
rect 14749 15997 14783 16031
rect 15117 15997 15151 16031
rect 19533 15997 19567 16031
rect 19809 15997 19843 16031
rect 19165 15861 19199 15895
rect 1501 15657 1535 15691
rect 19993 15589 20027 15623
rect 1685 15521 1719 15555
rect 1961 15521 1995 15555
rect 19257 15521 19291 15555
rect 19717 15521 19751 15555
rect 14749 15317 14783 15351
rect 19257 15113 19291 15147
rect 19625 15113 19659 15147
rect 14197 14977 14231 15011
rect 1685 14909 1719 14943
rect 13461 14909 13495 14943
rect 13921 14909 13955 14943
rect 2053 14773 2087 14807
rect 13277 14773 13311 14807
rect 1593 14569 1627 14603
rect 13553 14569 13587 14603
rect 20637 13889 20671 13923
rect 1593 13821 1627 13855
rect 1961 13821 1995 13855
rect 19809 13821 19843 13855
rect 20177 13821 20211 13855
rect 20361 13821 20395 13855
rect 1501 13685 1535 13719
rect 1685 13481 1719 13515
rect 19901 13481 19935 13515
rect 10057 12937 10091 12971
rect 19349 12937 19383 12971
rect 20269 12801 20303 12835
rect 10241 12733 10275 12767
rect 10793 12733 10827 12767
rect 19533 12733 19567 12767
rect 19993 12733 20027 12767
rect 10333 12597 10367 12631
rect 1501 12393 1535 12427
rect 19625 12393 19659 12427
rect 21649 12325 21683 12359
rect 1685 12257 1719 12291
rect 1961 12257 1995 12291
rect 20913 12257 20947 12291
rect 21373 12257 21407 12291
rect 10333 12053 10367 12087
rect 2053 11849 2087 11883
rect 20913 11849 20947 11883
rect 1685 11645 1719 11679
rect 21281 11509 21315 11543
rect 1593 11305 1627 11339
rect 20729 10761 20763 10795
rect 21649 10625 21683 10659
rect 1593 10557 1627 10591
rect 1961 10557 1995 10591
rect 20913 10557 20947 10591
rect 21373 10557 21407 10591
rect 1501 10421 1535 10455
rect 20361 10421 20395 10455
rect 1685 10217 1719 10251
rect 21189 10081 21223 10115
rect 21465 10081 21499 10115
rect 21649 10081 21683 10115
rect 18337 9469 18371 9503
rect 20821 9469 20855 9503
rect 21005 9469 21039 9503
rect 18981 9401 19015 9435
rect 20453 9401 20487 9435
rect 17877 9333 17911 9367
rect 20821 9333 20855 9367
rect 21557 9333 21591 9367
rect 1501 9129 1535 9163
rect 6837 9129 6871 9163
rect 18981 9129 19015 9163
rect 1593 8993 1627 9027
rect 1961 8993 1995 9027
rect 6561 8993 6595 9027
rect 7113 8993 7147 9027
rect 18245 8993 18279 9027
rect 18337 8993 18371 9027
rect 19349 8993 19383 9027
rect 17877 8925 17911 8959
rect 18705 8925 18739 8959
rect 18613 8857 18647 8891
rect 20637 8857 20671 8891
rect 18475 8789 18509 8823
rect 21097 8789 21131 8823
rect 1685 8585 1719 8619
rect 1961 8585 1995 8619
rect 6561 8585 6595 8619
rect 17785 8585 17819 8619
rect 18337 8585 18371 8619
rect 19073 8585 19107 8619
rect 18751 8517 18785 8551
rect 18889 8517 18923 8551
rect 18981 8449 19015 8483
rect 20177 8449 20211 8483
rect 18613 8381 18647 8415
rect 20085 8381 20119 8415
rect 20269 8381 20303 8415
rect 17509 8313 17543 8347
rect 7113 8245 7147 8279
rect 19717 8245 19751 8279
rect 1593 8041 1627 8075
rect 18337 8041 18371 8075
rect 19073 8041 19107 8075
rect 18429 7973 18463 8007
rect 21649 7973 21683 8007
rect 21189 7905 21223 7939
rect 21465 7905 21499 7939
rect 18797 7837 18831 7871
rect 18705 7769 18739 7803
rect 17877 7701 17911 7735
rect 18567 7701 18601 7735
rect 19441 7701 19475 7735
rect 20361 7701 20395 7735
rect 17877 7497 17911 7531
rect 19441 7497 19475 7531
rect 20821 7497 20855 7531
rect 18521 7429 18555 7463
rect 18935 7429 18969 7463
rect 19073 7429 19107 7463
rect 20499 7429 20533 7463
rect 19165 7361 19199 7395
rect 1685 7293 1719 7327
rect 1869 7293 1903 7327
rect 19809 7293 19843 7327
rect 20591 7293 20625 7327
rect 20700 7293 20734 7327
rect 18797 7225 18831 7259
rect 20361 7225 20395 7259
rect 21373 7225 21407 7259
rect 21741 7225 21775 7259
rect 1501 7157 1535 7191
rect 17509 7157 17543 7191
rect 20269 7157 20303 7191
rect 22109 7157 22143 7191
rect 1685 6953 1719 6987
rect 18889 6953 18923 6987
rect 20085 6953 20119 6987
rect 18245 6885 18279 6919
rect 21649 6885 21683 6919
rect 16681 6817 16715 6851
rect 17020 6817 17054 6851
rect 19257 6817 19291 6851
rect 20913 6817 20947 6851
rect 21465 6817 21499 6851
rect 17141 6749 17175 6783
rect 18153 6749 18187 6783
rect 18613 6749 18647 6783
rect 18521 6681 18555 6715
rect 16497 6613 16531 6647
rect 16819 6613 16853 6647
rect 16957 6613 16991 6647
rect 17693 6613 17727 6647
rect 18383 6613 18417 6647
rect 19717 6613 19751 6647
rect 20453 6613 20487 6647
rect 7573 6409 7607 6443
rect 10609 6409 10643 6443
rect 15577 6409 15611 6443
rect 16681 6409 16715 6443
rect 20729 6409 20763 6443
rect 22293 6409 22327 6443
rect 17417 6341 17451 6375
rect 19349 6341 19383 6375
rect 15945 6273 15979 6307
rect 16773 6273 16807 6307
rect 19441 6273 19475 6307
rect 7757 6205 7791 6239
rect 8217 6205 8251 6239
rect 10885 6205 10919 6239
rect 11253 6205 11287 6239
rect 16405 6205 16439 6239
rect 16552 6205 16586 6239
rect 17877 6205 17911 6239
rect 19073 6205 19107 6239
rect 19220 6205 19254 6239
rect 19809 6205 19843 6239
rect 21189 6205 21223 6239
rect 21373 6205 21407 6239
rect 21649 6205 21683 6239
rect 8493 6137 8527 6171
rect 18245 6137 18279 6171
rect 21925 6137 21959 6171
rect 10793 6069 10827 6103
rect 16313 6069 16347 6103
rect 17049 6069 17083 6103
rect 18797 6069 18831 6103
rect 20177 6069 20211 6103
rect 2145 5865 2179 5899
rect 15393 5865 15427 5899
rect 20637 5865 20671 5899
rect 21557 5865 21591 5899
rect 18613 5797 18647 5831
rect 19533 5797 19567 5831
rect 2605 5729 2639 5763
rect 2789 5729 2823 5763
rect 15301 5729 15335 5763
rect 15853 5729 15887 5763
rect 17325 5729 17359 5763
rect 17969 5729 18003 5763
rect 18797 5729 18831 5763
rect 19809 5729 19843 5763
rect 20913 5729 20947 5763
rect 2881 5661 2915 5695
rect 19165 5661 19199 5695
rect 21281 5661 21315 5695
rect 19073 5593 19107 5627
rect 7849 5525 7883 5559
rect 10793 5525 10827 5559
rect 16405 5525 16439 5559
rect 16865 5525 16899 5559
rect 18935 5525 18969 5559
rect 20177 5525 20211 5559
rect 21051 5525 21085 5559
rect 21189 5525 21223 5559
rect 3525 5321 3559 5355
rect 15393 5321 15427 5355
rect 16773 5321 16807 5355
rect 18981 5321 19015 5355
rect 22293 5321 22327 5355
rect 17877 5253 17911 5287
rect 18659 5253 18693 5287
rect 18797 5253 18831 5287
rect 19533 5253 19567 5287
rect 20361 5253 20395 5287
rect 2053 5185 2087 5219
rect 18429 5185 18463 5219
rect 18889 5185 18923 5219
rect 20729 5185 20763 5219
rect 21925 5185 21959 5219
rect 2145 5117 2179 5151
rect 2697 5117 2731 5151
rect 18521 5117 18555 5151
rect 20913 5117 20947 5151
rect 21373 5117 21407 5151
rect 21649 5117 21683 5151
rect 3249 5049 3283 5083
rect 15761 5049 15795 5083
rect 1593 4981 1627 5015
rect 2237 4981 2271 5015
rect 17325 4981 17359 5015
rect 19993 4981 20027 5015
rect 17969 4777 18003 4811
rect 18337 4777 18371 4811
rect 19809 4777 19843 4811
rect 20637 4777 20671 4811
rect 18429 4709 18463 4743
rect 1593 4641 1627 4675
rect 11161 4641 11195 4675
rect 11437 4641 11471 4675
rect 12541 4641 12575 4675
rect 13001 4641 13035 4675
rect 15761 4641 15795 4675
rect 16313 4641 16347 4675
rect 20913 4641 20947 4675
rect 21373 4641 21407 4675
rect 2145 4573 2179 4607
rect 11621 4573 11655 4607
rect 13277 4573 13311 4607
rect 16497 4573 16531 4607
rect 18797 4573 18831 4607
rect 21649 4573 21683 4607
rect 18889 4505 18923 4539
rect 2513 4437 2547 4471
rect 2881 4437 2915 4471
rect 18567 4437 18601 4471
rect 18705 4437 18739 4471
rect 19441 4437 19475 4471
rect 4445 4233 4479 4267
rect 10977 4233 11011 4267
rect 12633 4233 12667 4267
rect 15853 4233 15887 4267
rect 16313 4233 16347 4267
rect 17877 4233 17911 4267
rect 18521 4233 18555 4267
rect 18889 4233 18923 4267
rect 2789 4165 2823 4199
rect 2881 4165 2915 4199
rect 19349 4165 19383 4199
rect 19717 4165 19751 4199
rect 1593 4097 1627 4131
rect 3065 4097 3099 4131
rect 4629 4097 4663 4131
rect 19441 4097 19475 4131
rect 21833 4097 21867 4131
rect 22201 4097 22235 4131
rect 1501 4029 1535 4063
rect 1777 4029 1811 4063
rect 2789 4029 2823 4063
rect 3157 4029 3191 4063
rect 4721 4029 4755 4063
rect 9229 4029 9263 4063
rect 9321 4029 9355 4063
rect 9781 4029 9815 4063
rect 11345 4029 11379 4063
rect 16497 4029 16531 4063
rect 19220 4029 19254 4063
rect 20821 4029 20855 4063
rect 21281 4029 21315 4063
rect 2237 3961 2271 3995
rect 10057 3961 10091 3995
rect 17141 3961 17175 3995
rect 19073 3961 19107 3995
rect 21557 3961 21591 3995
rect 2513 3893 2547 3927
rect 13093 3893 13127 3927
rect 15485 3893 15519 3927
rect 20269 3893 20303 3927
rect 20637 3893 20671 3927
rect 4169 3689 4203 3723
rect 9413 3689 9447 3723
rect 19625 3689 19659 3723
rect 1593 3621 1627 3655
rect 19993 3621 20027 3655
rect 2145 3553 2179 3587
rect 2237 3553 2271 3587
rect 2421 3553 2455 3587
rect 3893 3553 3927 3587
rect 4077 3553 4111 3587
rect 4537 3553 4571 3587
rect 17049 3553 17083 3587
rect 18613 3553 18647 3587
rect 20913 3553 20947 3587
rect 21373 3553 21407 3587
rect 2881 3485 2915 3519
rect 17417 3485 17451 3519
rect 18061 3485 18095 3519
rect 18981 3485 19015 3519
rect 21649 3485 21683 3519
rect 18429 3417 18463 3451
rect 18751 3417 18785 3451
rect 18889 3417 18923 3451
rect 1961 3349 1995 3383
rect 3249 3349 3283 3383
rect 17187 3349 17221 3383
rect 17325 3349 17359 3383
rect 17509 3349 17543 3383
rect 19073 3349 19107 3383
rect 2513 3145 2547 3179
rect 2881 3145 2915 3179
rect 3341 3145 3375 3179
rect 5641 3145 5675 3179
rect 16773 3145 16807 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 18337 3145 18371 3179
rect 21557 3145 21591 3179
rect 1593 3077 1627 3111
rect 17141 3077 17175 3111
rect 18705 3077 18739 3111
rect 1961 3009 1995 3043
rect 4169 3009 4203 3043
rect 20085 3009 20119 3043
rect 20361 3009 20395 3043
rect 1501 2941 1535 2975
rect 1777 2941 1811 2975
rect 4813 2941 4847 2975
rect 5089 2941 5123 2975
rect 19257 2941 19291 2975
rect 19441 2941 19475 2975
rect 19717 2941 19751 2975
rect 20821 2941 20855 2975
rect 21005 2941 21039 2975
rect 5273 2873 5307 2907
rect 21281 2873 21315 2907
rect 3801 2805 3835 2839
rect 1961 2601 1995 2635
rect 2881 2601 2915 2635
rect 3249 2601 3283 2635
rect 3801 2601 3835 2635
rect 4169 2601 4203 2635
rect 5181 2601 5215 2635
rect 7021 2601 7055 2635
rect 17141 2601 17175 2635
rect 18429 2601 18463 2635
rect 19717 2601 19751 2635
rect 20637 2601 20671 2635
rect 2513 2533 2547 2567
rect 6745 2533 6779 2567
rect 18153 2533 18187 2567
rect 1501 2465 1535 2499
rect 1593 2465 1627 2499
rect 1777 2465 1811 2499
rect 4353 2465 4387 2499
rect 4629 2465 4663 2499
rect 6377 2465 6411 2499
rect 7205 2465 7239 2499
rect 7389 2465 7423 2499
rect 17785 2465 17819 2499
rect 18337 2465 18371 2499
rect 18797 2465 18831 2499
rect 20913 2397 20947 2431
rect 19441 2261 19475 2295
<< metal1 >>
rect 842 23196 848 23248
rect 900 23236 906 23248
rect 1762 23236 1768 23248
rect 900 23208 1768 23236
rect 900 23196 906 23208
rect 1762 23196 1768 23208
rect 1820 23196 1826 23248
rect 20714 22652 20720 22704
rect 20772 22692 20778 22704
rect 21726 22692 21732 22704
rect 20772 22664 21732 22692
rect 20772 22652 20778 22664
rect 21726 22652 21732 22664
rect 21784 22652 21790 22704
rect 106 22040 112 22092
rect 164 22080 170 22092
rect 17954 22080 17960 22092
rect 164 22052 17960 22080
rect 164 22040 170 22052
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 17954 21128 17960 21140
rect 17915 21100 17960 21128
rect 17954 21088 17960 21100
rect 18012 21088 18018 21140
rect 18322 21088 18328 21140
rect 18380 21088 18386 21140
rect 17037 21063 17095 21069
rect 17037 21029 17049 21063
rect 17083 21060 17095 21063
rect 18340 21060 18368 21088
rect 17083 21032 18368 21060
rect 21637 21063 21695 21069
rect 17083 21029 17095 21032
rect 17037 21023 17095 21029
rect 21637 21029 21649 21063
rect 21683 21060 21695 21063
rect 23014 21060 23020 21072
rect 21683 21032 23020 21060
rect 21683 21029 21695 21032
rect 21637 21023 21695 21029
rect 23014 21020 23020 21032
rect 23072 21020 23078 21072
rect 16298 20992 16304 21004
rect 16259 20964 16304 20992
rect 16298 20952 16304 20964
rect 16356 20952 16362 21004
rect 16482 20952 16488 21004
rect 16540 20992 16546 21004
rect 16761 20995 16819 21001
rect 16761 20992 16773 20995
rect 16540 20964 16773 20992
rect 16540 20952 16546 20964
rect 16761 20961 16773 20964
rect 16807 20961 16819 20995
rect 16761 20955 16819 20961
rect 18141 20995 18199 21001
rect 18141 20961 18153 20995
rect 18187 20961 18199 20995
rect 18414 20992 18420 21004
rect 18375 20964 18420 20992
rect 18141 20955 18199 20961
rect 18156 20924 18184 20955
rect 18414 20952 18420 20964
rect 18472 20952 18478 21004
rect 20622 20952 20628 21004
rect 20680 20992 20686 21004
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 20680 20964 20913 20992
rect 20680 20952 20686 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 21450 20992 21456 21004
rect 21411 20964 21456 20992
rect 20901 20955 20959 20961
rect 21450 20952 21456 20964
rect 21508 20952 21514 21004
rect 18156 20896 19288 20924
rect 19260 20797 19288 20896
rect 19245 20791 19303 20797
rect 19245 20757 19257 20791
rect 19291 20788 19303 20791
rect 19426 20788 19432 20800
rect 19291 20760 19432 20788
rect 19291 20757 19303 20760
rect 19245 20751 19303 20757
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 106 20544 112 20596
rect 164 20584 170 20596
rect 164 20556 15792 20584
rect 164 20544 170 20556
rect 14645 20519 14703 20525
rect 14645 20516 14657 20519
rect 10796 20488 14657 20516
rect 4522 20448 4528 20460
rect 4483 20420 4528 20448
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 8386 20448 8392 20460
rect 8347 20420 8392 20448
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 1486 20340 1492 20392
rect 1544 20380 1550 20392
rect 3513 20383 3571 20389
rect 3513 20380 3525 20383
rect 1544 20352 3525 20380
rect 1544 20340 1550 20352
rect 3513 20349 3525 20352
rect 3559 20380 3571 20383
rect 4154 20380 4160 20392
rect 3559 20352 4160 20380
rect 3559 20349 3571 20352
rect 3513 20343 3571 20349
rect 4154 20340 4160 20352
rect 4212 20380 4218 20392
rect 4433 20383 4491 20389
rect 4212 20352 4305 20380
rect 4212 20340 4218 20352
rect 4433 20349 4445 20383
rect 4479 20380 4491 20383
rect 4982 20380 4988 20392
rect 4479 20352 4988 20380
rect 4479 20349 4491 20352
rect 4433 20343 4491 20349
rect 3881 20315 3939 20321
rect 3881 20281 3893 20315
rect 3927 20312 3939 20315
rect 4062 20312 4068 20324
rect 3927 20284 4068 20312
rect 3927 20281 3939 20284
rect 3881 20275 3939 20281
rect 4062 20272 4068 20284
rect 4120 20312 4126 20324
rect 4448 20312 4476 20343
rect 4982 20340 4988 20352
rect 5040 20340 5046 20392
rect 7745 20383 7803 20389
rect 7745 20349 7757 20383
rect 7791 20380 7803 20383
rect 8110 20380 8116 20392
rect 7791 20352 8116 20380
rect 7791 20349 7803 20352
rect 7745 20343 7803 20349
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 8297 20383 8355 20389
rect 8297 20349 8309 20383
rect 8343 20380 8355 20383
rect 8478 20380 8484 20392
rect 8343 20352 8484 20380
rect 8343 20349 8355 20352
rect 8297 20343 8355 20349
rect 8478 20340 8484 20352
rect 8536 20340 8542 20392
rect 10796 20389 10824 20488
rect 14645 20485 14657 20488
rect 14691 20485 14703 20519
rect 14645 20479 14703 20485
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20448 11575 20451
rect 11606 20448 11612 20460
rect 11563 20420 11612 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20448 13231 20451
rect 13262 20448 13268 20460
rect 13219 20420 13268 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 10781 20383 10839 20389
rect 10781 20349 10793 20383
rect 10827 20349 10839 20383
rect 10781 20343 10839 20349
rect 4120 20284 4476 20312
rect 4120 20272 4126 20284
rect 8018 20204 8024 20256
rect 8076 20244 8082 20256
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 8076 20216 10609 20244
rect 8076 20204 8082 20216
rect 10597 20213 10609 20216
rect 10643 20244 10655 20247
rect 10796 20244 10824 20343
rect 10870 20340 10876 20392
rect 10928 20380 10934 20392
rect 11241 20383 11299 20389
rect 11241 20380 11253 20383
rect 10928 20352 11253 20380
rect 10928 20340 10934 20352
rect 11241 20349 11253 20352
rect 11287 20349 11299 20383
rect 11241 20343 11299 20349
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20349 12495 20383
rect 12437 20343 12495 20349
rect 10643 20216 10824 20244
rect 12253 20247 12311 20253
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 12253 20213 12265 20247
rect 12299 20244 12311 20247
rect 12452 20244 12480 20343
rect 12802 20340 12808 20392
rect 12860 20380 12866 20392
rect 12897 20383 12955 20389
rect 12897 20380 12909 20383
rect 12860 20352 12909 20380
rect 12860 20340 12866 20352
rect 12897 20349 12909 20352
rect 12943 20349 12955 20383
rect 14660 20380 14688 20479
rect 15764 20457 15792 20556
rect 18414 20476 18420 20528
rect 18472 20516 18478 20528
rect 20349 20519 20407 20525
rect 20349 20516 20361 20519
rect 18472 20488 20361 20516
rect 18472 20476 18478 20488
rect 20349 20485 20361 20488
rect 20395 20516 20407 20519
rect 20717 20519 20775 20525
rect 20717 20516 20729 20519
rect 20395 20488 20729 20516
rect 20395 20485 20407 20488
rect 20349 20479 20407 20485
rect 20717 20485 20729 20488
rect 20763 20516 20775 20519
rect 20763 20488 21496 20516
rect 20763 20485 20775 20488
rect 20717 20479 20775 20485
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 19889 20451 19947 20457
rect 18739 20420 19472 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 19444 20392 19472 20420
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 20438 20448 20444 20460
rect 19935 20420 20444 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 21468 20392 21496 20488
rect 21634 20448 21640 20460
rect 21595 20420 21640 20448
rect 21634 20408 21640 20420
rect 21692 20408 21698 20460
rect 15194 20380 15200 20392
rect 14660 20352 15200 20380
rect 12897 20343 12955 20349
rect 15194 20340 15200 20352
rect 15252 20340 15258 20392
rect 15657 20383 15715 20389
rect 15657 20349 15669 20383
rect 15703 20380 15715 20383
rect 19426 20380 19432 20392
rect 15703 20352 19012 20380
rect 19387 20352 19432 20380
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 15105 20315 15163 20321
rect 15105 20281 15117 20315
rect 15151 20312 15163 20315
rect 15672 20312 15700 20343
rect 16298 20312 16304 20324
rect 15151 20284 15700 20312
rect 16211 20284 16304 20312
rect 15151 20281 15163 20284
rect 15105 20275 15163 20281
rect 16298 20272 16304 20284
rect 16356 20312 16362 20324
rect 16669 20315 16727 20321
rect 16669 20312 16681 20315
rect 16356 20284 16681 20312
rect 16356 20272 16362 20284
rect 16669 20281 16681 20284
rect 16715 20281 16727 20315
rect 16669 20275 16727 20281
rect 18984 20312 19012 20352
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20349 19671 20383
rect 20898 20380 20904 20392
rect 20859 20352 20904 20380
rect 19613 20343 19671 20349
rect 19628 20312 19656 20343
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 21450 20340 21456 20392
rect 21508 20380 21514 20392
rect 21508 20352 21601 20380
rect 21508 20340 21514 20352
rect 18984 20284 19656 20312
rect 20916 20312 20944 20340
rect 21913 20315 21971 20321
rect 21913 20312 21925 20315
rect 20916 20284 21925 20312
rect 13538 20244 13544 20256
rect 12299 20216 13544 20244
rect 12299 20213 12311 20216
rect 12253 20207 12311 20213
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 14734 20204 14740 20256
rect 14792 20244 14798 20256
rect 16316 20244 16344 20272
rect 18984 20256 19012 20284
rect 21913 20281 21925 20284
rect 21959 20281 21971 20315
rect 21913 20275 21971 20281
rect 14792 20216 16344 20244
rect 16393 20247 16451 20253
rect 14792 20204 14798 20216
rect 16393 20213 16405 20247
rect 16439 20244 16451 20247
rect 16482 20244 16488 20256
rect 16439 20216 16488 20244
rect 16439 20213 16451 20216
rect 16393 20207 16451 20213
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 18325 20247 18383 20253
rect 18325 20213 18337 20247
rect 18371 20244 18383 20247
rect 18414 20244 18420 20256
rect 18371 20216 18420 20244
rect 18371 20213 18383 20216
rect 18325 20207 18383 20213
rect 18414 20204 18420 20216
rect 18472 20204 18478 20256
rect 18966 20244 18972 20256
rect 18927 20216 18972 20244
rect 18966 20204 18972 20216
rect 19024 20204 19030 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 22281 20247 22339 20253
rect 22281 20244 22293 20247
rect 20680 20216 22293 20244
rect 20680 20204 20686 20216
rect 22281 20213 22293 20216
rect 22327 20213 22339 20247
rect 22281 20207 22339 20213
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4212 20012 8064 20040
rect 4212 20000 4218 20012
rect 5261 19975 5319 19981
rect 5261 19941 5273 19975
rect 5307 19972 5319 19975
rect 5626 19972 5632 19984
rect 5307 19944 5632 19972
rect 5307 19941 5319 19944
rect 5261 19935 5319 19941
rect 5626 19932 5632 19944
rect 5684 19932 5690 19984
rect 8036 19916 8064 20012
rect 8757 19975 8815 19981
rect 8757 19941 8769 19975
rect 8803 19972 8815 19975
rect 9490 19972 9496 19984
rect 8803 19944 9496 19972
rect 8803 19941 8815 19944
rect 8757 19935 8815 19941
rect 9490 19932 9496 19944
rect 9548 19932 9554 19984
rect 16666 19972 16672 19984
rect 16627 19944 16672 19972
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 19242 19972 19248 19984
rect 18524 19944 19104 19972
rect 19203 19944 19248 19972
rect 18524 19916 18552 19944
rect 4798 19904 4804 19916
rect 4759 19876 4804 19904
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 4982 19904 4988 19916
rect 4943 19876 4988 19904
rect 4982 19864 4988 19876
rect 5040 19864 5046 19916
rect 8018 19904 8024 19916
rect 7931 19876 8024 19904
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8478 19904 8484 19916
rect 8439 19876 8484 19904
rect 8478 19864 8484 19876
rect 8536 19864 8542 19916
rect 16206 19904 16212 19916
rect 16167 19876 16212 19904
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 16482 19904 16488 19916
rect 16443 19876 16488 19904
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 18506 19904 18512 19916
rect 18467 19876 18512 19904
rect 18506 19864 18512 19876
rect 18564 19864 18570 19916
rect 18966 19904 18972 19916
rect 18879 19876 18972 19904
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 19076 19904 19104 19944
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 21637 19975 21695 19981
rect 21637 19941 21649 19975
rect 21683 19972 21695 19975
rect 23566 19972 23572 19984
rect 21683 19944 23572 19972
rect 21683 19941 21695 19944
rect 21637 19935 21695 19941
rect 23566 19932 23572 19944
rect 23624 19932 23630 19984
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 19076 19876 20913 19904
rect 20901 19873 20913 19876
rect 20947 19904 20959 19907
rect 21266 19904 21272 19916
rect 20947 19876 21272 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 21450 19904 21456 19916
rect 21411 19876 21456 19904
rect 21450 19864 21456 19876
rect 21508 19864 21514 19916
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 8496 19836 8524 19864
rect 7975 19808 8524 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 18322 19796 18328 19848
rect 18380 19836 18386 19848
rect 18984 19836 19012 19864
rect 18380 19808 19012 19836
rect 18380 19796 18386 19808
rect 10870 19700 10876 19712
rect 10831 19672 10876 19700
rect 10870 19660 10876 19672
rect 10928 19700 10934 19712
rect 12437 19703 12495 19709
rect 12437 19700 12449 19703
rect 10928 19672 12449 19700
rect 10928 19660 10934 19672
rect 12437 19669 12449 19672
rect 12483 19700 12495 19703
rect 12802 19700 12808 19712
rect 12483 19672 12808 19700
rect 12483 19669 12495 19672
rect 12437 19663 12495 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 8018 19496 8024 19508
rect 7979 19468 8024 19496
rect 8018 19456 8024 19468
rect 8076 19456 8082 19508
rect 21266 19496 21272 19508
rect 21227 19468 21272 19496
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 20993 19431 21051 19437
rect 20993 19397 21005 19431
rect 21039 19428 21051 19431
rect 21450 19428 21456 19440
rect 21039 19400 21456 19428
rect 21039 19397 21051 19400
rect 20993 19391 21051 19397
rect 21450 19388 21456 19400
rect 21508 19388 21514 19440
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16393 19363 16451 19369
rect 16393 19360 16405 19363
rect 16264 19332 16405 19360
rect 16264 19320 16270 19332
rect 16393 19329 16405 19332
rect 16439 19360 16451 19363
rect 19426 19360 19432 19372
rect 16439 19332 19432 19360
rect 16439 19329 16451 19332
rect 16393 19323 16451 19329
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 19610 19360 19616 19372
rect 19571 19332 19616 19360
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 16224 19292 16252 19320
rect 15948 19264 16252 19292
rect 4062 19184 4068 19236
rect 4120 19224 4126 19236
rect 4617 19227 4675 19233
rect 4617 19224 4629 19227
rect 4120 19196 4629 19224
rect 4120 19184 4126 19196
rect 4617 19193 4629 19196
rect 4663 19224 4675 19227
rect 5442 19224 5448 19236
rect 4663 19196 5448 19224
rect 4663 19193 4675 19196
rect 4617 19187 4675 19193
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 13538 19184 13544 19236
rect 13596 19224 13602 19236
rect 15948 19224 15976 19264
rect 18506 19252 18512 19304
rect 18564 19292 18570 19304
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18564 19264 18889 19292
rect 18564 19252 18570 19264
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 19334 19292 19340 19304
rect 19295 19264 19340 19292
rect 18877 19255 18935 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 13596 19196 15976 19224
rect 16025 19227 16083 19233
rect 13596 19184 13602 19196
rect 16025 19193 16037 19227
rect 16071 19224 16083 19227
rect 16482 19224 16488 19236
rect 16071 19196 16488 19224
rect 16071 19193 16083 19196
rect 16025 19187 16083 19193
rect 16482 19184 16488 19196
rect 16540 19224 16546 19236
rect 18138 19224 18144 19236
rect 16540 19196 18144 19224
rect 16540 19184 16546 19196
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 4985 19159 5043 19165
rect 4985 19156 4997 19159
rect 4856 19128 4997 19156
rect 4856 19116 4862 19128
rect 4985 19125 4997 19128
rect 5031 19156 5043 19159
rect 5810 19156 5816 19168
rect 5031 19128 5816 19156
rect 5031 19125 5043 19128
rect 4985 19119 5043 19125
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 8478 19156 8484 19168
rect 8391 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19156 8542 19168
rect 9306 19156 9312 19168
rect 8536 19128 9312 19156
rect 8536 19116 8542 19128
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 18509 19159 18567 19165
rect 18509 19156 18521 19159
rect 18380 19128 18521 19156
rect 18380 19116 18386 19128
rect 18509 19125 18521 19128
rect 18555 19125 18567 19159
rect 18509 19119 18567 19125
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 21637 18887 21695 18893
rect 21637 18853 21649 18887
rect 21683 18884 21695 18887
rect 23566 18884 23572 18896
rect 21683 18856 23572 18884
rect 21683 18853 21695 18856
rect 21637 18847 21695 18853
rect 23566 18844 23572 18856
rect 23624 18844 23630 18896
rect 1486 18816 1492 18828
rect 1447 18788 1492 18816
rect 1486 18776 1492 18788
rect 1544 18776 1550 18828
rect 1670 18776 1676 18828
rect 1728 18816 1734 18828
rect 1949 18819 2007 18825
rect 1949 18816 1961 18819
rect 1728 18788 1961 18816
rect 1728 18776 1734 18788
rect 1949 18785 1961 18788
rect 1995 18785 2007 18819
rect 1949 18779 2007 18785
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20622 18816 20628 18828
rect 20036 18788 20628 18816
rect 20036 18776 20042 18788
rect 20622 18776 20628 18788
rect 20680 18816 20686 18828
rect 20901 18819 20959 18825
rect 20901 18816 20913 18819
rect 20680 18788 20913 18816
rect 20680 18776 20686 18788
rect 20901 18785 20913 18788
rect 20947 18785 20959 18819
rect 21358 18816 21364 18828
rect 21319 18788 21364 18816
rect 20901 18779 20959 18785
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 18506 18748 18512 18760
rect 18467 18720 18512 18748
rect 18506 18708 18512 18720
rect 18564 18748 18570 18760
rect 18966 18748 18972 18760
rect 18564 18720 18972 18748
rect 18564 18708 18570 18720
rect 18966 18708 18972 18720
rect 19024 18748 19030 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19024 18720 19257 18748
rect 19024 18708 19030 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 18138 18640 18144 18692
rect 18196 18680 18202 18692
rect 18877 18683 18935 18689
rect 18877 18680 18889 18683
rect 18196 18652 18889 18680
rect 18196 18640 18202 18652
rect 18877 18649 18889 18652
rect 18923 18680 18935 18683
rect 19334 18680 19340 18692
rect 18923 18652 19340 18680
rect 18923 18649 18935 18652
rect 18877 18643 18935 18649
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 1486 18368 1492 18420
rect 1544 18408 1550 18420
rect 1949 18411 2007 18417
rect 1949 18408 1961 18411
rect 1544 18380 1961 18408
rect 1544 18368 1550 18380
rect 1949 18377 1961 18380
rect 1995 18377 2007 18411
rect 1949 18371 2007 18377
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 20806 18204 20812 18216
rect 19484 18176 20812 18204
rect 19484 18164 19490 18176
rect 20806 18164 20812 18176
rect 20864 18204 20870 18216
rect 20901 18207 20959 18213
rect 20901 18204 20913 18207
rect 20864 18176 20913 18204
rect 20864 18164 20870 18176
rect 20901 18173 20913 18176
rect 20947 18173 20959 18207
rect 21358 18204 21364 18216
rect 21271 18176 21364 18204
rect 20901 18167 20959 18173
rect 21358 18164 21364 18176
rect 21416 18164 21422 18216
rect 21634 18204 21640 18216
rect 21595 18176 21640 18204
rect 21634 18164 21640 18176
rect 21692 18164 21698 18216
rect 17862 18096 17868 18148
rect 17920 18136 17926 18148
rect 20349 18139 20407 18145
rect 20349 18136 20361 18139
rect 17920 18108 20361 18136
rect 17920 18096 17926 18108
rect 20349 18105 20361 18108
rect 20395 18136 20407 18139
rect 20717 18139 20775 18145
rect 20717 18136 20729 18139
rect 20395 18108 20729 18136
rect 20395 18105 20407 18108
rect 20349 18099 20407 18105
rect 20717 18105 20729 18108
rect 20763 18136 20775 18139
rect 21376 18136 21404 18164
rect 20763 18108 21404 18136
rect 20763 18105 20775 18108
rect 20717 18099 20775 18105
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 19978 18068 19984 18080
rect 14792 18040 19984 18068
rect 14792 18028 14798 18040
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 1578 17824 1584 17876
rect 1636 17864 1642 17876
rect 1673 17867 1731 17873
rect 1673 17864 1685 17867
rect 1636 17836 1685 17864
rect 1636 17824 1642 17836
rect 1673 17833 1685 17836
rect 1719 17864 1731 17867
rect 8110 17864 8116 17876
rect 1719 17836 8116 17864
rect 1719 17833 1731 17836
rect 1673 17827 1731 17833
rect 8110 17824 8116 17836
rect 8168 17824 8174 17876
rect 20806 17484 20812 17536
rect 20864 17524 20870 17536
rect 21085 17527 21143 17533
rect 21085 17524 21097 17527
rect 20864 17496 21097 17524
rect 20864 17484 20870 17496
rect 21085 17493 21097 17496
rect 21131 17493 21143 17527
rect 21085 17487 21143 17493
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 1670 17076 1676 17128
rect 1728 17116 1734 17128
rect 1857 17119 1915 17125
rect 1857 17116 1869 17119
rect 1728 17088 1869 17116
rect 1728 17076 1734 17088
rect 1857 17085 1869 17088
rect 1903 17085 1915 17119
rect 1857 17079 1915 17085
rect 106 16940 112 16992
rect 164 16980 170 16992
rect 1489 16983 1547 16989
rect 1489 16980 1501 16983
rect 164 16952 1501 16980
rect 164 16940 170 16952
rect 1489 16949 1501 16952
rect 1535 16949 1547 16983
rect 1489 16943 1547 16949
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 19429 16779 19487 16785
rect 19429 16745 19441 16779
rect 19475 16776 19487 16779
rect 19518 16776 19524 16788
rect 19475 16748 19524 16776
rect 19475 16745 19487 16748
rect 19429 16739 19487 16745
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16096 14611 16099
rect 15378 16096 15384 16108
rect 14599 16068 15148 16096
rect 15339 16068 15384 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 14734 16028 14740 16040
rect 14695 16000 14740 16028
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 15120 16037 15148 16068
rect 15378 16056 15384 16068
rect 15436 16056 15442 16108
rect 20070 16096 20076 16108
rect 20031 16068 20076 16096
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 16028 15163 16031
rect 19242 16028 19248 16040
rect 15151 16000 19248 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 19518 16028 19524 16040
rect 19479 16000 19524 16028
rect 19518 15988 19524 16000
rect 19576 15988 19582 16040
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 19812 15960 19840 15991
rect 19168 15932 19840 15960
rect 19168 15904 19196 15932
rect 19150 15892 19156 15904
rect 19111 15864 19156 15892
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1489 15691 1547 15697
rect 1489 15688 1501 15691
rect 1452 15660 1501 15688
rect 1452 15648 1458 15660
rect 1489 15657 1501 15660
rect 1535 15657 1547 15691
rect 1489 15651 1547 15657
rect 19518 15620 19524 15632
rect 19260 15592 19524 15620
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15521 1731 15555
rect 1946 15552 1952 15564
rect 1907 15524 1952 15552
rect 1673 15515 1731 15521
rect 1688 15484 1716 15515
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 19260 15561 19288 15592
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 19981 15623 20039 15629
rect 19981 15589 19993 15623
rect 20027 15620 20039 15623
rect 23566 15620 23572 15632
rect 20027 15592 23572 15620
rect 20027 15589 20039 15592
rect 19981 15583 20039 15589
rect 23566 15580 23572 15592
rect 23624 15580 23630 15632
rect 19245 15555 19303 15561
rect 19245 15521 19257 15555
rect 19291 15521 19303 15555
rect 19245 15515 19303 15521
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19705 15555 19763 15561
rect 19705 15552 19717 15555
rect 19392 15524 19717 15552
rect 19392 15512 19398 15524
rect 19705 15521 19717 15524
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 2038 15484 2044 15496
rect 1688 15456 2044 15484
rect 2038 15444 2044 15456
rect 2096 15444 2102 15496
rect 14734 15348 14740 15360
rect 14695 15320 14740 15348
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 19242 15144 19248 15156
rect 18932 15116 19248 15144
rect 18932 15104 18938 15116
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 19576 15116 19625 15144
rect 19576 15104 19582 15116
rect 19613 15113 19625 15116
rect 19659 15113 19671 15147
rect 19613 15107 19671 15113
rect 11882 14968 11888 15020
rect 11940 15008 11946 15020
rect 13538 15008 13544 15020
rect 11940 14980 13544 15008
rect 11940 14968 11946 14980
rect 13538 14968 13544 14980
rect 13596 15008 13602 15020
rect 14182 15008 14188 15020
rect 13596 14980 13814 15008
rect 14143 14980 14188 15008
rect 13596 14968 13602 14980
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 1946 14940 1952 14952
rect 1719 14912 1952 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13280 14912 13461 14940
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 13280 14813 13308 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13786 14940 13814 14980
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13786 14912 13921 14940
rect 13449 14903 13507 14909
rect 13909 14909 13921 14912
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 12492 14776 13277 14804
rect 12492 14764 12498 14776
rect 13265 14773 13277 14776
rect 13311 14773 13323 14807
rect 13265 14767 13323 14773
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 19518 13880 19524 13932
rect 19576 13920 19582 13932
rect 20625 13923 20683 13929
rect 19576 13892 20392 13920
rect 19576 13880 19582 13892
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 19797 13855 19855 13861
rect 19797 13852 19809 13855
rect 12492 13824 19809 13852
rect 12492 13812 12498 13824
rect 19797 13821 19809 13824
rect 19843 13852 19855 13855
rect 20162 13852 20168 13864
rect 19843 13824 20168 13852
rect 19843 13821 19855 13824
rect 19797 13815 19855 13821
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20364 13861 20392 13892
rect 20625 13889 20637 13923
rect 20671 13920 20683 13923
rect 23566 13920 23572 13932
rect 20671 13892 23572 13920
rect 20671 13889 20683 13892
rect 20625 13883 20683 13889
rect 23566 13880 23572 13892
rect 23624 13880 23630 13932
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20438 13852 20444 13864
rect 20395 13824 20444 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 106 13676 112 13728
rect 164 13716 170 13728
rect 1489 13719 1547 13725
rect 1489 13716 1501 13719
rect 164 13688 1501 13716
rect 164 13676 170 13688
rect 1489 13685 1501 13688
rect 1535 13685 1547 13719
rect 19886 13716 19892 13728
rect 19799 13688 19892 13716
rect 1489 13679 1547 13685
rect 19886 13676 19892 13688
rect 19944 13716 19950 13728
rect 20438 13716 20444 13728
rect 19944 13688 20444 13716
rect 19944 13676 19950 13688
rect 20438 13676 20444 13688
rect 20496 13676 20502 13728
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 1946 13512 1952 13524
rect 1719 13484 1952 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 19886 13512 19892 13524
rect 19847 13484 19892 13512
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 5810 12928 5816 12980
rect 5868 12968 5874 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 5868 12940 10057 12968
rect 5868 12928 5874 12940
rect 10045 12937 10057 12940
rect 10091 12937 10103 12971
rect 10045 12931 10103 12937
rect 10060 12832 10088 12931
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 19337 12971 19395 12977
rect 19337 12968 19349 12971
rect 19024 12940 19349 12968
rect 19024 12928 19030 12940
rect 19337 12937 19349 12940
rect 19383 12937 19395 12971
rect 19337 12931 19395 12937
rect 11146 12832 11152 12844
rect 10060 12804 11152 12832
rect 10060 12764 10088 12804
rect 11146 12792 11152 12804
rect 11204 12832 11210 12844
rect 14734 12832 14740 12844
rect 11204 12804 14740 12832
rect 11204 12792 11210 12804
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 10229 12767 10287 12773
rect 10229 12764 10241 12767
rect 10060 12736 10241 12764
rect 10229 12733 10241 12736
rect 10275 12733 10287 12767
rect 10778 12764 10784 12776
rect 10739 12736 10784 12764
rect 10229 12727 10287 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 19352 12764 19380 12931
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 19518 12764 19524 12776
rect 19352 12736 19524 12764
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 19610 12724 19616 12776
rect 19668 12764 19674 12776
rect 19981 12767 20039 12773
rect 19981 12764 19993 12767
rect 19668 12736 19993 12764
rect 19668 12724 19674 12736
rect 19981 12733 19993 12736
rect 20027 12733 20039 12767
rect 19981 12727 20039 12733
rect 10318 12628 10324 12640
rect 10279 12600 10324 12628
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 1489 12427 1547 12433
rect 1489 12393 1501 12427
rect 1535 12393 1547 12427
rect 19610 12424 19616 12436
rect 19571 12396 19616 12424
rect 1489 12387 1547 12393
rect 1302 12316 1308 12368
rect 1360 12356 1366 12368
rect 1504 12356 1532 12387
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 2038 12356 2044 12368
rect 1360 12328 1532 12356
rect 1688 12328 2044 12356
rect 1360 12316 1366 12328
rect 1688 12297 1716 12328
rect 2038 12316 2044 12328
rect 2096 12316 2102 12368
rect 21637 12359 21695 12365
rect 21637 12325 21649 12359
rect 21683 12356 21695 12359
rect 23566 12356 23572 12368
rect 21683 12328 23572 12356
rect 21683 12325 21695 12328
rect 21637 12319 21695 12325
rect 23566 12316 23572 12328
rect 23624 12316 23630 12368
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12257 1731 12291
rect 1946 12288 1952 12300
rect 1907 12260 1952 12288
rect 1673 12251 1731 12257
rect 1946 12248 1952 12260
rect 2004 12248 2010 12300
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20864 12260 20913 12288
rect 20864 12248 20870 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 21266 12248 21272 12300
rect 21324 12288 21330 12300
rect 21361 12291 21419 12297
rect 21361 12288 21373 12291
rect 21324 12260 21373 12288
rect 21324 12248 21330 12260
rect 21361 12257 21373 12260
rect 21407 12257 21419 12291
rect 21361 12251 21419 12257
rect 10321 12087 10379 12093
rect 10321 12053 10333 12087
rect 10367 12084 10379 12087
rect 10778 12084 10784 12096
rect 10367 12056 10784 12084
rect 10367 12053 10379 12056
rect 10321 12047 10379 12053
rect 10778 12044 10784 12056
rect 10836 12084 10842 12096
rect 11422 12084 11428 12096
rect 10836 12056 11428 12084
rect 10836 12044 10842 12056
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20864 11852 20913 11880
rect 20864 11840 20870 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 1946 11676 1952 11688
rect 1719 11648 1952 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 21266 11540 21272 11552
rect 21227 11512 21272 11540
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 20717 10795 20775 10801
rect 20717 10792 20729 10795
rect 19576 10764 20729 10792
rect 19576 10752 19582 10764
rect 20717 10761 20729 10764
rect 20763 10761 20775 10795
rect 20717 10755 20775 10761
rect 1578 10588 1584 10600
rect 1539 10560 1584 10588
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 20732 10588 20760 10755
rect 21634 10656 21640 10668
rect 21595 10628 21640 10656
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 20901 10591 20959 10597
rect 20901 10588 20913 10591
rect 20680 10560 20913 10588
rect 20680 10548 20686 10560
rect 20901 10557 20913 10560
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 21266 10520 21272 10532
rect 20364 10492 21272 10520
rect 106 10412 112 10464
rect 164 10452 170 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 164 10424 1501 10452
rect 164 10412 170 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 19702 10412 19708 10464
rect 19760 10452 19766 10464
rect 20364 10461 20392 10492
rect 21266 10480 21272 10492
rect 21324 10520 21330 10532
rect 21376 10520 21404 10551
rect 21324 10492 21404 10520
rect 21324 10480 21330 10492
rect 20349 10455 20407 10461
rect 20349 10452 20361 10455
rect 19760 10424 20361 10452
rect 19760 10412 19766 10424
rect 20349 10421 20361 10424
rect 20395 10421 20407 10455
rect 20349 10415 20407 10421
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1946 10248 1952 10260
rect 1719 10220 1952 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 21177 10115 21235 10121
rect 21177 10081 21189 10115
rect 21223 10112 21235 10115
rect 21266 10112 21272 10124
rect 21223 10084 21272 10112
rect 21223 10081 21235 10084
rect 21177 10075 21235 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21450 10112 21456 10124
rect 21411 10084 21456 10112
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 21637 10115 21695 10121
rect 21637 10081 21649 10115
rect 21683 10112 21695 10115
rect 23566 10112 23572 10124
rect 21683 10084 23572 10112
rect 21683 10081 21695 10084
rect 21637 10075 21695 10081
rect 23566 10072 23572 10084
rect 23624 10072 23630 10124
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 13722 9908 13728 9920
rect 10928 9880 13728 9908
rect 10928 9868 10934 9880
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 19610 9568 19616 9580
rect 13780 9540 19616 9568
rect 13780 9528 13786 9540
rect 19610 9528 19616 9540
rect 19668 9528 19674 9580
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 18248 9472 18337 9500
rect 18248 9376 18276 9472
rect 18325 9469 18337 9472
rect 18371 9469 18383 9503
rect 20806 9500 20812 9512
rect 20767 9472 20812 9500
rect 18325 9463 18383 9469
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 20916 9472 21005 9500
rect 18969 9435 19027 9441
rect 18969 9401 18981 9435
rect 19015 9432 19027 9435
rect 19426 9432 19432 9444
rect 19015 9404 19432 9432
rect 19015 9401 19027 9404
rect 18969 9395 19027 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 19576 9404 20453 9432
rect 19576 9392 19582 9404
rect 20441 9401 20453 9404
rect 20487 9432 20499 9435
rect 20916 9432 20944 9472
rect 20993 9469 21005 9472
rect 21039 9469 21051 9503
rect 20993 9463 21051 9469
rect 20487 9404 20944 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 17865 9367 17923 9373
rect 17865 9333 17877 9367
rect 17911 9364 17923 9367
rect 18230 9364 18236 9376
rect 17911 9336 18236 9364
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 20714 9324 20720 9376
rect 20772 9364 20778 9376
rect 20809 9367 20867 9373
rect 20809 9364 20821 9367
rect 20772 9336 20821 9364
rect 20772 9324 20778 9336
rect 20809 9333 20821 9336
rect 20855 9333 20867 9367
rect 20809 9327 20867 9333
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 21545 9367 21603 9373
rect 21545 9364 21557 9367
rect 21416 9336 21557 9364
rect 21416 9324 21422 9336
rect 21545 9333 21557 9336
rect 21591 9333 21603 9367
rect 21545 9327 21603 9333
rect 1104 9274 22816 9296
rect 106 9188 112 9240
rect 164 9228 170 9240
rect 164 9200 980 9228
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 164 9188 170 9200
rect 952 9160 980 9200
rect 1489 9163 1547 9169
rect 1489 9160 1501 9163
rect 952 9132 1501 9160
rect 1489 9129 1501 9132
rect 1535 9129 1547 9163
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 1489 9123 1547 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 18969 9163 19027 9169
rect 18969 9160 18981 9163
rect 17920 9132 18981 9160
rect 17920 9120 17926 9132
rect 18969 9129 18981 9132
rect 19015 9129 19027 9163
rect 18969 9123 19027 9129
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 18690 9092 18696 9104
rect 17828 9064 18696 9092
rect 17828 9052 17834 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 8993 1639 9027
rect 1946 9024 1952 9036
rect 1907 8996 1952 9024
rect 1581 8987 1639 8993
rect 1596 8956 1624 8987
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 6546 9024 6552 9036
rect 6507 8996 6552 9024
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 7098 9024 7104 9036
rect 7059 8996 7104 9024
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 18233 9027 18291 9033
rect 18233 8993 18245 9027
rect 18279 9024 18291 9027
rect 18325 9027 18383 9033
rect 18325 9024 18337 9027
rect 18279 8996 18337 9024
rect 18279 8993 18291 8996
rect 18233 8987 18291 8993
rect 18325 8993 18337 8996
rect 18371 9024 18383 9027
rect 18598 9024 18604 9036
rect 18371 8996 18604 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 18598 8984 18604 8996
rect 18656 9024 18662 9036
rect 19337 9027 19395 9033
rect 19337 9024 19349 9027
rect 18656 8996 19349 9024
rect 18656 8984 18662 8996
rect 19337 8993 19349 8996
rect 19383 8993 19395 9027
rect 19337 8987 19395 8993
rect 1670 8956 1676 8968
rect 1596 8928 1676 8956
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8956 17923 8959
rect 18506 8956 18512 8968
rect 17911 8928 18512 8956
rect 17911 8925 17923 8928
rect 17865 8919 17923 8925
rect 18506 8916 18512 8928
rect 18564 8956 18570 8968
rect 18564 8928 18644 8956
rect 18564 8916 18570 8928
rect 18616 8897 18644 8928
rect 18690 8916 18696 8968
rect 18748 8956 18754 8968
rect 18966 8956 18972 8968
rect 18748 8928 18972 8956
rect 18748 8916 18754 8928
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8857 18659 8891
rect 18601 8851 18659 8857
rect 20625 8891 20683 8897
rect 20625 8857 20637 8891
rect 20671 8888 20683 8891
rect 20806 8888 20812 8900
rect 20671 8860 20812 8888
rect 20671 8857 20683 8860
rect 20625 8851 20683 8857
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 18230 8780 18236 8832
rect 18288 8820 18294 8832
rect 18463 8823 18521 8829
rect 18463 8820 18475 8823
rect 18288 8792 18475 8820
rect 18288 8780 18294 8792
rect 18463 8789 18475 8792
rect 18509 8789 18521 8823
rect 18463 8783 18521 8789
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21085 8823 21143 8829
rect 21085 8820 21097 8823
rect 20772 8792 21097 8820
rect 20772 8780 20778 8792
rect 21085 8789 21097 8792
rect 21131 8820 21143 8823
rect 21450 8820 21456 8832
rect 21131 8792 21456 8820
rect 21131 8789 21143 8792
rect 21085 8783 21143 8789
rect 21450 8780 21456 8792
rect 21508 8780 21514 8832
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8616 2010 8628
rect 2590 8616 2596 8628
rect 2004 8588 2596 8616
rect 2004 8576 2010 8588
rect 2590 8576 2596 8588
rect 2648 8616 2654 8628
rect 6546 8616 6552 8628
rect 2648 8588 6552 8616
rect 2648 8576 2654 8588
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 17770 8616 17776 8628
rect 17731 8588 17776 8616
rect 17770 8576 17776 8588
rect 17828 8616 17834 8628
rect 18325 8619 18383 8625
rect 18325 8616 18337 8619
rect 17828 8588 18337 8616
rect 17828 8576 17834 8588
rect 18325 8585 18337 8588
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 18472 8588 19073 8616
rect 18472 8576 18478 8588
rect 19061 8585 19073 8588
rect 19107 8585 19119 8619
rect 19061 8579 19119 8585
rect 18739 8551 18797 8557
rect 18739 8548 18751 8551
rect 18432 8520 18751 8548
rect 17497 8347 17555 8353
rect 17497 8313 17509 8347
rect 17543 8344 17555 8347
rect 18230 8344 18236 8356
rect 17543 8316 18236 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 18432 8344 18460 8520
rect 18739 8517 18751 8520
rect 18785 8517 18797 8551
rect 18739 8511 18797 8517
rect 18877 8551 18935 8557
rect 18877 8517 18889 8551
rect 18923 8548 18935 8551
rect 18923 8520 20208 8548
rect 18923 8517 18935 8520
rect 18877 8511 18935 8517
rect 18506 8440 18512 8492
rect 18564 8480 18570 8492
rect 18892 8480 18920 8511
rect 18564 8452 18920 8480
rect 18564 8440 18570 8452
rect 18966 8440 18972 8492
rect 19024 8480 19030 8492
rect 20180 8489 20208 8520
rect 20165 8483 20223 8489
rect 19024 8452 19069 8480
rect 19024 8440 19030 8452
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 18598 8412 18604 8424
rect 18559 8384 18604 8412
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19116 8384 20085 8412
rect 19116 8372 19122 8384
rect 20073 8381 20085 8384
rect 20119 8412 20131 8415
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 20119 8384 20269 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 20257 8375 20315 8381
rect 18432 8316 19472 8344
rect 19444 8288 19472 8316
rect 7098 8276 7104 8288
rect 7011 8248 7104 8276
rect 7098 8236 7104 8248
rect 7156 8276 7162 8288
rect 7834 8276 7840 8288
rect 7156 8248 7840 8276
rect 7156 8236 7162 8248
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 19705 8279 19763 8285
rect 19705 8276 19717 8279
rect 19484 8248 19717 8276
rect 19484 8236 19490 8248
rect 19705 8245 19717 8248
rect 19751 8245 19763 8279
rect 19705 8239 19763 8245
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 18325 8075 18383 8081
rect 18325 8041 18337 8075
rect 18371 8072 18383 8075
rect 18598 8072 18604 8084
rect 18371 8044 18604 8072
rect 18371 8041 18383 8044
rect 18325 8035 18383 8041
rect 18432 8013 18460 8044
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19061 8075 19119 8081
rect 19061 8072 19073 8075
rect 18932 8044 19073 8072
rect 18932 8032 18938 8044
rect 19061 8041 19073 8044
rect 19107 8041 19119 8075
rect 19061 8035 19119 8041
rect 18417 8007 18475 8013
rect 18417 8004 18429 8007
rect 18395 7976 18429 8004
rect 18417 7973 18429 7976
rect 18463 7973 18475 8007
rect 18417 7967 18475 7973
rect 21637 8007 21695 8013
rect 21637 7973 21649 8007
rect 21683 8004 21695 8007
rect 23566 8004 23572 8016
rect 21683 7976 23572 8004
rect 21683 7973 21695 7976
rect 21637 7967 21695 7973
rect 23566 7964 23572 7976
rect 23624 7964 23630 8016
rect 20806 7896 20812 7948
rect 20864 7936 20870 7948
rect 21177 7939 21235 7945
rect 21177 7936 21189 7939
rect 20864 7908 21189 7936
rect 20864 7896 20870 7908
rect 21177 7905 21189 7908
rect 21223 7905 21235 7939
rect 21450 7936 21456 7948
rect 21411 7908 21456 7936
rect 21177 7899 21235 7905
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18966 7868 18972 7880
rect 18831 7840 18972 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 21192 7868 21220 7899
rect 21450 7896 21456 7908
rect 21508 7896 21514 7948
rect 21726 7868 21732 7880
rect 21192 7840 21732 7868
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 18690 7800 18696 7812
rect 18603 7772 18696 7800
rect 18690 7760 18696 7772
rect 18748 7800 18754 7812
rect 19058 7800 19064 7812
rect 18748 7772 19064 7800
rect 18748 7760 18754 7772
rect 19058 7760 19064 7772
rect 19116 7760 19122 7812
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 17552 7704 17877 7732
rect 17552 7692 17558 7704
rect 17865 7701 17877 7704
rect 17911 7701 17923 7735
rect 17865 7695 17923 7701
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 18555 7735 18613 7741
rect 18555 7732 18567 7735
rect 18288 7704 18567 7732
rect 18288 7692 18294 7704
rect 18555 7701 18567 7704
rect 18601 7701 18613 7735
rect 18555 7695 18613 7701
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19392 7704 19441 7732
rect 19392 7692 19398 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 20346 7732 20352 7744
rect 20307 7704 20352 7732
rect 19429 7695 19487 7701
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 17865 7531 17923 7537
rect 17865 7497 17877 7531
rect 17911 7528 17923 7531
rect 18414 7528 18420 7540
rect 17911 7500 18420 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 18414 7488 18420 7500
rect 18472 7528 18478 7540
rect 18690 7528 18696 7540
rect 18472 7500 18696 7528
rect 18472 7488 18478 7500
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 19610 7528 19616 7540
rect 19475 7500 19616 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 20162 7488 20168 7540
rect 20220 7528 20226 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 20220 7500 20821 7528
rect 20220 7488 20226 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 18966 7469 18972 7472
rect 18509 7463 18567 7469
rect 18509 7460 18521 7463
rect 17368 7432 18521 7460
rect 17368 7420 17374 7432
rect 18509 7429 18521 7432
rect 18555 7460 18567 7463
rect 18923 7463 18972 7469
rect 18923 7460 18935 7463
rect 18555 7432 18935 7460
rect 18555 7429 18567 7432
rect 18509 7423 18567 7429
rect 18923 7429 18935 7432
rect 18969 7429 18972 7463
rect 18923 7423 18972 7429
rect 18966 7420 18972 7423
rect 19024 7420 19030 7472
rect 19061 7463 19119 7469
rect 19061 7429 19073 7463
rect 19107 7460 19119 7463
rect 19334 7460 19340 7472
rect 19107 7432 19340 7460
rect 19107 7429 19119 7432
rect 19061 7423 19119 7429
rect 19334 7420 19340 7432
rect 19392 7460 19398 7472
rect 19392 7432 20300 7460
rect 19392 7420 19398 7432
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 19153 7395 19211 7401
rect 1636 7364 1900 7392
rect 1636 7352 1642 7364
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 1872 7333 1900 7364
rect 19153 7361 19165 7395
rect 19199 7392 19211 7395
rect 19426 7392 19432 7404
rect 19199 7364 19432 7392
rect 19199 7361 19211 7364
rect 19153 7355 19211 7361
rect 19426 7352 19432 7364
rect 19484 7392 19490 7404
rect 19610 7392 19616 7404
rect 19484 7364 19616 7392
rect 19484 7352 19490 7364
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 20272 7336 20300 7432
rect 20346 7420 20352 7472
rect 20404 7460 20410 7472
rect 20487 7463 20545 7469
rect 20487 7460 20499 7463
rect 20404 7432 20499 7460
rect 20404 7420 20410 7432
rect 20487 7429 20499 7432
rect 20533 7429 20545 7463
rect 20487 7423 20545 7429
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7293 1915 7327
rect 1857 7287 1915 7293
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 19797 7327 19855 7333
rect 19797 7324 19809 7327
rect 18288 7296 19809 7324
rect 18288 7284 18294 7296
rect 19797 7293 19809 7296
rect 19843 7293 19855 7327
rect 19797 7287 19855 7293
rect 20254 7284 20260 7336
rect 20312 7324 20318 7336
rect 20714 7333 20720 7336
rect 20579 7327 20637 7333
rect 20579 7324 20591 7327
rect 20312 7296 20591 7324
rect 20312 7284 20318 7296
rect 20579 7293 20591 7296
rect 20625 7293 20637 7327
rect 20579 7287 20637 7293
rect 20688 7327 20720 7333
rect 20688 7293 20700 7327
rect 20688 7287 20720 7293
rect 20714 7284 20720 7287
rect 20772 7284 20778 7336
rect 18506 7256 18512 7268
rect 17512 7228 18512 7256
rect 17512 7200 17540 7228
rect 18506 7216 18512 7228
rect 18564 7256 18570 7268
rect 18785 7259 18843 7265
rect 18785 7256 18797 7259
rect 18564 7228 18797 7256
rect 18564 7216 18570 7228
rect 18785 7225 18797 7228
rect 18831 7256 18843 7259
rect 20349 7259 20407 7265
rect 20349 7256 20361 7259
rect 18831 7228 20361 7256
rect 18831 7225 18843 7228
rect 18785 7219 18843 7225
rect 20349 7225 20361 7228
rect 20395 7256 20407 7259
rect 21361 7259 21419 7265
rect 21361 7256 21373 7259
rect 20395 7228 21373 7256
rect 20395 7225 20407 7228
rect 20349 7219 20407 7225
rect 21361 7225 21373 7228
rect 21407 7225 21419 7259
rect 21726 7256 21732 7268
rect 21687 7228 21732 7256
rect 21361 7219 21419 7225
rect 21726 7216 21732 7228
rect 21784 7216 21790 7268
rect 106 7148 112 7200
rect 164 7188 170 7200
rect 1489 7191 1547 7197
rect 1489 7188 1501 7191
rect 164 7160 1501 7188
rect 164 7148 170 7160
rect 1489 7157 1501 7160
rect 1535 7157 1547 7191
rect 17494 7188 17500 7200
rect 17455 7160 17500 7188
rect 1489 7151 1547 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 21450 7148 21456 7200
rect 21508 7188 21514 7200
rect 22097 7191 22155 7197
rect 22097 7188 22109 7191
rect 21508 7160 22109 7188
rect 21508 7148 21514 7160
rect 22097 7157 22109 7160
rect 22143 7157 22155 7191
rect 22097 7151 22155 7157
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 1670 6984 1676 6996
rect 1631 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 18877 6987 18935 6993
rect 18877 6984 18889 6987
rect 18196 6956 18889 6984
rect 18196 6944 18202 6956
rect 18877 6953 18889 6956
rect 18923 6953 18935 6987
rect 18877 6947 18935 6953
rect 19242 6944 19248 6996
rect 19300 6984 19306 6996
rect 19610 6984 19616 6996
rect 19300 6956 19616 6984
rect 19300 6944 19306 6956
rect 19610 6944 19616 6956
rect 19668 6944 19674 6996
rect 20073 6987 20131 6993
rect 20073 6953 20085 6987
rect 20119 6984 20131 6987
rect 20346 6984 20352 6996
rect 20119 6956 20352 6984
rect 20119 6953 20131 6956
rect 20073 6947 20131 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 18233 6919 18291 6925
rect 18233 6885 18245 6919
rect 18279 6916 18291 6919
rect 18598 6916 18604 6928
rect 18279 6888 18604 6916
rect 18279 6885 18291 6888
rect 18233 6879 18291 6885
rect 18598 6876 18604 6888
rect 18656 6876 18662 6928
rect 21637 6919 21695 6925
rect 21637 6885 21649 6919
rect 21683 6916 21695 6919
rect 23566 6916 23572 6928
rect 21683 6888 23572 6916
rect 21683 6885 21695 6888
rect 21637 6879 21695 6885
rect 23566 6876 23572 6888
rect 23624 6876 23630 6928
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16540 6820 16681 6848
rect 16540 6808 16546 6820
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 16669 6811 16727 6817
rect 17008 6851 17066 6857
rect 17008 6817 17020 6851
rect 17054 6848 17066 6851
rect 17310 6848 17316 6860
rect 17054 6820 17316 6848
rect 17054 6817 17066 6820
rect 17008 6811 17066 6817
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 18966 6808 18972 6860
rect 19024 6848 19030 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 19024 6820 19257 6848
rect 19024 6808 19030 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 20530 6808 20536 6860
rect 20588 6848 20594 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20588 6820 20913 6848
rect 20588 6808 20594 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 21450 6848 21456 6860
rect 21411 6820 21456 6848
rect 20901 6811 20959 6817
rect 17126 6780 17132 6792
rect 17087 6752 17132 6780
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 17276 6752 18153 6780
rect 17276 6740 17282 6752
rect 18141 6749 18153 6752
rect 18187 6780 18199 6783
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18187 6752 18613 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 18601 6749 18613 6752
rect 18647 6780 18659 6783
rect 19426 6780 19432 6792
rect 18647 6752 19432 6780
rect 18647 6749 18659 6752
rect 18601 6743 18659 6749
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 20916 6780 20944 6811
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 22278 6780 22284 6792
rect 20916 6752 22284 6780
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 18509 6715 18567 6721
rect 18509 6712 18521 6715
rect 17696 6684 18521 6712
rect 16482 6644 16488 6656
rect 16443 6616 16488 6644
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 16807 6647 16865 6653
rect 16807 6644 16819 6647
rect 16724 6616 16819 6644
rect 16724 6604 16730 6616
rect 16807 6613 16819 6616
rect 16853 6613 16865 6647
rect 16942 6644 16948 6656
rect 16903 6616 16948 6644
rect 16807 6607 16865 6613
rect 16942 6604 16948 6616
rect 17000 6644 17006 6656
rect 17494 6644 17500 6656
rect 17000 6616 17500 6644
rect 17000 6604 17006 6616
rect 17494 6604 17500 6616
rect 17552 6644 17558 6656
rect 17696 6653 17724 6684
rect 18509 6681 18521 6684
rect 18555 6712 18567 6715
rect 19334 6712 19340 6724
rect 18555 6684 19340 6712
rect 18555 6681 18567 6684
rect 18509 6675 18567 6681
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17552 6616 17693 6644
rect 17552 6604 17558 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17681 6607 17739 6613
rect 18230 6604 18236 6656
rect 18288 6644 18294 6656
rect 18371 6647 18429 6653
rect 18371 6644 18383 6647
rect 18288 6616 18383 6644
rect 18288 6604 18294 6616
rect 18371 6613 18383 6616
rect 18417 6613 18429 6647
rect 18371 6607 18429 6613
rect 19610 6604 19616 6656
rect 19668 6644 19674 6656
rect 19705 6647 19763 6653
rect 19705 6644 19717 6647
rect 19668 6616 19717 6644
rect 19668 6604 19674 6616
rect 19705 6613 19717 6616
rect 19751 6644 19763 6647
rect 20441 6647 20499 6653
rect 20441 6644 20453 6647
rect 19751 6616 20453 6644
rect 19751 6613 19763 6616
rect 19705 6607 19763 6613
rect 20441 6613 20453 6616
rect 20487 6644 20499 6647
rect 20530 6644 20536 6656
rect 20487 6616 20536 6644
rect 20487 6613 20499 6616
rect 20441 6607 20499 6613
rect 20530 6604 20536 6616
rect 20588 6644 20594 6656
rect 20714 6644 20720 6656
rect 20588 6616 20720 6644
rect 20588 6604 20594 6616
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 1578 6400 1584 6452
rect 1636 6440 1642 6452
rect 1854 6440 1860 6452
rect 1636 6412 1860 6440
rect 1636 6400 1642 6412
rect 1854 6400 1860 6412
rect 1912 6440 1918 6452
rect 7561 6443 7619 6449
rect 7561 6440 7573 6443
rect 1912 6412 7573 6440
rect 1912 6400 1918 6412
rect 7561 6409 7573 6412
rect 7607 6409 7619 6443
rect 7561 6403 7619 6409
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10870 6440 10876 6452
rect 10643 6412 10876 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 7576 6236 7604 6403
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 15565 6443 15623 6449
rect 15565 6409 15577 6443
rect 15611 6440 15623 6443
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 15611 6412 16681 6440
rect 15611 6409 15623 6412
rect 15565 6403 15623 6409
rect 16669 6409 16681 6412
rect 16715 6440 16727 6443
rect 16758 6440 16764 6452
rect 16715 6412 16764 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 16758 6400 16764 6412
rect 16816 6440 16822 6452
rect 16942 6440 16948 6452
rect 16816 6412 16948 6440
rect 16816 6400 16822 6412
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 17126 6400 17132 6452
rect 17184 6440 17190 6452
rect 20717 6443 20775 6449
rect 20717 6440 20729 6443
rect 17184 6412 20729 6440
rect 17184 6400 17190 6412
rect 20717 6409 20729 6412
rect 20763 6440 20775 6443
rect 21266 6440 21272 6452
rect 20763 6412 21272 6440
rect 20763 6409 20775 6412
rect 20717 6403 20775 6409
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 22278 6440 22284 6452
rect 22239 6412 22284 6440
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 17310 6332 17316 6384
rect 17368 6372 17374 6384
rect 17405 6375 17463 6381
rect 17405 6372 17417 6375
rect 17368 6344 17417 6372
rect 17368 6332 17374 6344
rect 17405 6341 17417 6344
rect 17451 6341 17463 6375
rect 19334 6372 19340 6384
rect 19295 6344 19340 6372
rect 17405 6335 17463 6341
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16761 6307 16819 6313
rect 16761 6304 16773 6307
rect 15979 6276 16773 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16761 6273 16773 6276
rect 16807 6304 16819 6307
rect 17218 6304 17224 6316
rect 16807 6276 17224 6304
rect 16807 6273 16819 6276
rect 16761 6267 16819 6273
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 19426 6304 19432 6316
rect 19339 6276 19432 6304
rect 19426 6264 19432 6276
rect 19484 6304 19490 6316
rect 20346 6304 20352 6316
rect 19484 6276 20352 6304
rect 19484 6264 19490 6276
rect 20346 6264 20352 6276
rect 20404 6264 20410 6316
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 7576 6208 7757 6236
rect 7745 6205 7757 6208
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 7892 6208 8217 6236
rect 7892 6196 7898 6208
rect 8205 6205 8217 6208
rect 8251 6205 8263 6239
rect 10870 6236 10876 6248
rect 10831 6208 10876 6236
rect 8205 6199 8263 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11238 6236 11244 6248
rect 11199 6208 11244 6236
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 16390 6236 16396 6248
rect 16351 6208 16396 6236
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16540 6239 16598 6245
rect 16540 6205 16552 6239
rect 16586 6236 16598 6239
rect 16666 6236 16672 6248
rect 16586 6208 16672 6236
rect 16586 6205 16598 6208
rect 16540 6199 16598 6205
rect 8478 6168 8484 6180
rect 8439 6140 8484 6168
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 16555 6168 16583 6199
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 17954 6236 17960 6248
rect 17911 6208 17960 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 17954 6196 17960 6208
rect 18012 6236 18018 6248
rect 18598 6236 18604 6248
rect 18012 6208 18604 6236
rect 18012 6196 18018 6208
rect 18598 6196 18604 6208
rect 18656 6236 18662 6248
rect 19242 6245 19248 6248
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18656 6208 19073 6236
rect 18656 6196 18662 6208
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19208 6239 19248 6245
rect 19208 6236 19220 6239
rect 19155 6208 19220 6236
rect 19061 6199 19119 6205
rect 19208 6205 19220 6208
rect 19208 6199 19248 6205
rect 19223 6196 19248 6199
rect 19300 6196 19306 6248
rect 19797 6239 19855 6245
rect 19797 6205 19809 6239
rect 19843 6236 19855 6239
rect 20714 6236 20720 6248
rect 19843 6208 20720 6236
rect 19843 6205 19855 6208
rect 19797 6199 19855 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 18230 6168 18236 6180
rect 16555 6140 18236 6168
rect 10778 6100 10784 6112
rect 10739 6072 10784 6100
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 16298 6100 16304 6112
rect 16259 6072 16304 6100
rect 16298 6060 16304 6072
rect 16356 6100 16362 6112
rect 16555 6100 16583 6140
rect 18230 6128 18236 6140
rect 18288 6128 18294 6180
rect 19223 6168 19251 6196
rect 18800 6140 19251 6168
rect 21192 6168 21220 6199
rect 21266 6196 21272 6248
rect 21324 6236 21330 6248
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 21324 6208 21373 6236
rect 21324 6196 21330 6208
rect 21361 6205 21373 6208
rect 21407 6205 21419 6239
rect 21634 6236 21640 6248
rect 21595 6208 21640 6236
rect 21361 6199 21419 6205
rect 21634 6196 21640 6208
rect 21692 6196 21698 6248
rect 21726 6168 21732 6180
rect 21192 6140 21732 6168
rect 16356 6072 16583 6100
rect 16356 6060 16362 6072
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 17037 6103 17095 6109
rect 17037 6100 17049 6103
rect 16908 6072 17049 6100
rect 16908 6060 16914 6072
rect 17037 6069 17049 6072
rect 17083 6069 17095 6103
rect 17037 6063 17095 6069
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 18800 6109 18828 6140
rect 21726 6128 21732 6140
rect 21784 6168 21790 6180
rect 21913 6171 21971 6177
rect 21913 6168 21925 6171
rect 21784 6140 21925 6168
rect 21784 6128 21790 6140
rect 21913 6137 21925 6140
rect 21959 6137 21971 6171
rect 21913 6131 21971 6137
rect 18785 6103 18843 6109
rect 18785 6100 18797 6103
rect 18748 6072 18797 6100
rect 18748 6060 18754 6072
rect 18785 6069 18797 6072
rect 18831 6069 18843 6103
rect 18785 6063 18843 6069
rect 20165 6103 20223 6109
rect 20165 6069 20177 6103
rect 20211 6100 20223 6103
rect 20530 6100 20536 6112
rect 20211 6072 20536 6100
rect 20211 6069 20223 6072
rect 20165 6063 20223 6069
rect 20530 6060 20536 6072
rect 20588 6100 20594 6112
rect 20990 6100 20996 6112
rect 20588 6072 20996 6100
rect 20588 6060 20594 6072
rect 20990 6060 20996 6072
rect 21048 6060 21054 6112
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 2133 5899 2191 5905
rect 2133 5896 2145 5899
rect 2096 5868 2145 5896
rect 2096 5856 2102 5868
rect 2133 5865 2145 5868
rect 2179 5865 2191 5899
rect 2133 5859 2191 5865
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 11238 5896 11244 5908
rect 7984 5868 11244 5896
rect 7984 5856 7990 5868
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 15378 5896 15384 5908
rect 15339 5868 15384 5896
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 16908 5868 20637 5896
rect 16908 5856 16914 5868
rect 20625 5865 20637 5868
rect 20671 5896 20683 5899
rect 21450 5896 21456 5908
rect 20671 5868 21456 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 21450 5856 21456 5868
rect 21508 5856 21514 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 21600 5868 21645 5896
rect 21600 5856 21606 5868
rect 18138 5828 18144 5840
rect 15856 5800 18144 5828
rect 2590 5760 2596 5772
rect 2551 5732 2596 5760
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 2774 5760 2780 5772
rect 2735 5732 2780 5760
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 15856 5769 15884 5800
rect 18138 5788 18144 5800
rect 18196 5788 18202 5840
rect 18414 5788 18420 5840
rect 18472 5828 18478 5840
rect 18601 5831 18659 5837
rect 18601 5828 18613 5831
rect 18472 5800 18613 5828
rect 18472 5788 18478 5800
rect 18601 5797 18613 5800
rect 18647 5797 18659 5831
rect 19518 5828 19524 5840
rect 19479 5800 19524 5828
rect 18601 5791 18659 5797
rect 19518 5788 19524 5800
rect 19576 5828 19582 5840
rect 20070 5828 20076 5840
rect 19576 5800 20076 5828
rect 19576 5788 19582 5800
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 15528 5732 15853 5760
rect 15528 5720 15534 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 17310 5760 17316 5772
rect 17271 5732 17316 5760
rect 15841 5723 15899 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17954 5760 17960 5772
rect 17915 5732 17960 5760
rect 17954 5720 17960 5732
rect 18012 5760 18018 5772
rect 18506 5760 18512 5772
rect 18012 5732 18512 5760
rect 18012 5720 18018 5732
rect 18506 5720 18512 5732
rect 18564 5760 18570 5772
rect 18785 5763 18843 5769
rect 18785 5760 18797 5763
rect 18564 5732 18797 5760
rect 18564 5720 18570 5732
rect 18785 5729 18797 5732
rect 18831 5760 18843 5763
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 18831 5732 19809 5760
rect 18831 5729 18843 5732
rect 18785 5723 18843 5729
rect 19797 5729 19809 5732
rect 19843 5729 19855 5763
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 19797 5723 19855 5729
rect 20824 5732 20913 5760
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 19153 5695 19211 5701
rect 19153 5661 19165 5695
rect 19199 5692 19211 5695
rect 19426 5692 19432 5704
rect 19199 5664 19432 5692
rect 19199 5661 19211 5664
rect 19153 5655 19211 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 18414 5584 18420 5636
rect 18472 5624 18478 5636
rect 18782 5624 18788 5636
rect 18472 5596 18788 5624
rect 18472 5584 18478 5596
rect 18782 5584 18788 5596
rect 18840 5624 18846 5636
rect 19061 5627 19119 5633
rect 19061 5624 19073 5627
rect 18840 5596 19073 5624
rect 18840 5584 18846 5596
rect 19061 5593 19073 5596
rect 19107 5624 19119 5627
rect 20824 5624 20852 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 21048 5664 21281 5692
rect 21048 5652 21054 5664
rect 21269 5661 21281 5664
rect 21315 5692 21327 5695
rect 22278 5692 22284 5704
rect 21315 5664 22284 5692
rect 21315 5661 21327 5664
rect 21269 5655 21327 5661
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 19107 5596 20852 5624
rect 19107 5593 19119 5596
rect 19061 5587 19119 5593
rect 7834 5556 7840 5568
rect 7795 5528 7840 5556
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 10781 5559 10839 5565
rect 10781 5525 10793 5559
rect 10827 5556 10839 5559
rect 11238 5556 11244 5568
rect 10827 5528 11244 5556
rect 10827 5525 10839 5528
rect 10781 5519 10839 5525
rect 11238 5516 11244 5528
rect 11296 5556 11302 5568
rect 12526 5556 12532 5568
rect 11296 5528 12532 5556
rect 11296 5516 11302 5528
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 16390 5556 16396 5568
rect 16351 5528 16396 5556
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 16482 5516 16488 5568
rect 16540 5556 16546 5568
rect 16853 5559 16911 5565
rect 16853 5556 16865 5559
rect 16540 5528 16865 5556
rect 16540 5516 16546 5528
rect 16853 5525 16865 5528
rect 16899 5556 16911 5559
rect 17310 5556 17316 5568
rect 16899 5528 17316 5556
rect 16899 5525 16911 5528
rect 16853 5519 16911 5525
rect 17310 5516 17316 5528
rect 17368 5516 17374 5568
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 18923 5559 18981 5565
rect 18923 5556 18935 5559
rect 18748 5528 18935 5556
rect 18748 5516 18754 5528
rect 18923 5525 18935 5528
rect 18969 5525 18981 5559
rect 18923 5519 18981 5525
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 20165 5559 20223 5565
rect 20165 5556 20177 5559
rect 19392 5528 20177 5556
rect 19392 5516 19398 5528
rect 20165 5525 20177 5528
rect 20211 5525 20223 5559
rect 20165 5519 20223 5525
rect 20806 5516 20812 5568
rect 20864 5556 20870 5568
rect 21039 5559 21097 5565
rect 21039 5556 21051 5559
rect 20864 5528 21051 5556
rect 20864 5516 20870 5528
rect 21039 5525 21051 5528
rect 21085 5525 21097 5559
rect 21039 5519 21097 5525
rect 21177 5559 21235 5565
rect 21177 5525 21189 5559
rect 21223 5556 21235 5559
rect 21450 5556 21456 5568
rect 21223 5528 21456 5556
rect 21223 5525 21235 5528
rect 21177 5519 21235 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 2590 5312 2596 5364
rect 2648 5352 2654 5364
rect 2958 5352 2964 5364
rect 2648 5324 2964 5352
rect 2648 5312 2654 5324
rect 2958 5312 2964 5324
rect 3016 5352 3022 5364
rect 3513 5355 3571 5361
rect 3513 5352 3525 5355
rect 3016 5324 3525 5352
rect 3016 5312 3022 5324
rect 3513 5321 3525 5324
rect 3559 5321 3571 5355
rect 3513 5315 3571 5321
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15470 5352 15476 5364
rect 15427 5324 15476 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 16758 5352 16764 5364
rect 16719 5324 16764 5352
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18969 5355 19027 5361
rect 18969 5352 18981 5355
rect 18380 5324 18981 5352
rect 18380 5312 18386 5324
rect 18969 5321 18981 5324
rect 19015 5321 19027 5355
rect 22278 5352 22284 5364
rect 22239 5324 22284 5352
rect 18969 5315 19027 5321
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 18690 5293 18696 5296
rect 17865 5287 17923 5293
rect 17865 5253 17877 5287
rect 17911 5284 17923 5287
rect 18647 5287 18696 5293
rect 18647 5284 18659 5287
rect 17911 5256 18659 5284
rect 17911 5253 17923 5256
rect 17865 5247 17923 5253
rect 18647 5253 18659 5256
rect 18693 5253 18696 5287
rect 18647 5247 18696 5253
rect 18690 5244 18696 5247
rect 18748 5244 18754 5296
rect 18782 5244 18788 5296
rect 18840 5284 18846 5296
rect 19521 5287 19579 5293
rect 19521 5284 19533 5287
rect 18840 5256 19533 5284
rect 18840 5244 18846 5256
rect 19521 5253 19533 5256
rect 19567 5284 19579 5287
rect 20162 5284 20168 5296
rect 19567 5256 20168 5284
rect 19567 5253 19579 5256
rect 19521 5247 19579 5253
rect 20162 5244 20168 5256
rect 20220 5284 20226 5296
rect 20349 5287 20407 5293
rect 20349 5284 20361 5287
rect 20220 5256 20361 5284
rect 20220 5244 20226 5256
rect 20349 5253 20361 5256
rect 20395 5253 20407 5287
rect 20349 5247 20407 5253
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2087 5188 2728 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2130 5148 2136 5160
rect 2091 5120 2136 5148
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 2700 5157 2728 5188
rect 16298 5176 16304 5228
rect 16356 5216 16362 5228
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 16356 5188 18429 5216
rect 16356 5176 16362 5188
rect 18417 5185 18429 5188
rect 18463 5216 18475 5219
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 18463 5188 18889 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 18877 5185 18889 5188
rect 18923 5216 18935 5219
rect 18966 5216 18972 5228
rect 18923 5188 18972 5216
rect 18923 5185 18935 5188
rect 18877 5179 18935 5185
rect 18966 5176 18972 5188
rect 19024 5216 19030 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 19024 5188 20729 5216
rect 19024 5176 19030 5188
rect 20717 5185 20729 5188
rect 20763 5216 20775 5219
rect 20806 5216 20812 5228
rect 20763 5188 20812 5216
rect 20763 5185 20775 5188
rect 20717 5179 20775 5185
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 21913 5219 21971 5225
rect 21913 5216 21925 5219
rect 21376 5188 21925 5216
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 2774 5148 2780 5160
rect 2731 5120 2780 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 2774 5108 2780 5120
rect 2832 5148 2838 5160
rect 18506 5148 18512 5160
rect 2832 5120 3280 5148
rect 18467 5120 18512 5148
rect 2832 5108 2838 5120
rect 3252 5089 3280 5120
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 19610 5148 19616 5160
rect 19306 5120 19616 5148
rect 3237 5083 3295 5089
rect 3237 5049 3249 5083
rect 3283 5080 3295 5083
rect 4154 5080 4160 5092
rect 3283 5052 4160 5080
rect 3283 5049 3295 5052
rect 3237 5043 3295 5049
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 15286 5040 15292 5092
rect 15344 5080 15350 5092
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 15344 5052 15761 5080
rect 15344 5040 15350 5052
rect 15749 5049 15761 5052
rect 15795 5080 15807 5083
rect 15795 5052 18460 5080
rect 15795 5049 15807 5052
rect 15749 5043 15807 5049
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 18432 5012 18460 5052
rect 18690 5040 18696 5092
rect 18748 5080 18754 5092
rect 19306 5080 19334 5120
rect 19610 5108 19616 5120
rect 19668 5108 19674 5160
rect 20622 5108 20628 5160
rect 20680 5148 20686 5160
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 20680 5120 20913 5148
rect 20680 5108 20686 5120
rect 20901 5117 20913 5120
rect 20947 5117 20959 5151
rect 20901 5111 20959 5117
rect 21266 5108 21272 5160
rect 21324 5148 21330 5160
rect 21376 5157 21404 5188
rect 21913 5185 21925 5188
rect 21959 5185 21971 5219
rect 21913 5179 21971 5185
rect 21361 5151 21419 5157
rect 21361 5148 21373 5151
rect 21324 5120 21373 5148
rect 21324 5108 21330 5120
rect 21361 5117 21373 5120
rect 21407 5117 21419 5151
rect 21634 5148 21640 5160
rect 21595 5120 21640 5148
rect 21361 5111 21419 5117
rect 21634 5108 21640 5120
rect 21692 5108 21698 5160
rect 18748 5052 19334 5080
rect 18748 5040 18754 5052
rect 19150 5012 19156 5024
rect 18432 4984 19156 5012
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19392 4984 19993 5012
rect 19392 4972 19398 4984
rect 19981 4981 19993 4984
rect 20027 5012 20039 5015
rect 20254 5012 20260 5024
rect 20027 4984 20260 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 20254 4972 20260 4984
rect 20312 5012 20318 5024
rect 21450 5012 21456 5024
rect 20312 4984 21456 5012
rect 20312 4972 20318 4984
rect 21450 4972 21456 4984
rect 21508 4972 21514 5024
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 17957 4811 18015 4817
rect 17957 4808 17969 4811
rect 17920 4780 17969 4808
rect 17920 4768 17926 4780
rect 17957 4777 17969 4780
rect 18003 4808 18015 4811
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 18003 4780 18337 4808
rect 18003 4777 18015 4780
rect 17957 4771 18015 4777
rect 18325 4777 18337 4780
rect 18371 4808 18383 4811
rect 18506 4808 18512 4820
rect 18371 4780 18512 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 15286 4740 15292 4752
rect 11164 4712 15292 4740
rect 1578 4672 1584 4684
rect 1539 4644 1584 4672
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 11164 4681 11192 4712
rect 15286 4700 15292 4712
rect 15344 4700 15350 4752
rect 18432 4749 18460 4780
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19484 4780 19809 4808
rect 19484 4768 19490 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 20622 4808 20628 4820
rect 20583 4780 20628 4808
rect 19797 4771 19855 4777
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 18395 4712 18429 4740
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 18417 4703 18475 4709
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 11020 4644 11161 4672
rect 11020 4632 11026 4644
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 11422 4672 11428 4684
rect 11383 4644 11428 4672
rect 11149 4635 11207 4641
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 12526 4672 12532 4684
rect 12487 4644 12532 4672
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 12618 4632 12624 4684
rect 12676 4672 12682 4684
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12676 4644 13001 4672
rect 12676 4632 12682 4644
rect 12989 4641 13001 4644
rect 13035 4672 13047 4675
rect 13035 4644 13814 4672
rect 13035 4641 13047 4644
rect 12989 4635 13047 4641
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 13262 4604 13268 4616
rect 13223 4576 13268 4604
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 13786 4536 13814 4644
rect 15470 4632 15476 4684
rect 15528 4672 15534 4684
rect 15749 4675 15807 4681
rect 15749 4672 15761 4675
rect 15528 4644 15761 4672
rect 15528 4632 15534 4644
rect 15749 4641 15761 4644
rect 15795 4641 15807 4675
rect 15749 4635 15807 4641
rect 15838 4632 15844 4684
rect 15896 4672 15902 4684
rect 16301 4675 16359 4681
rect 16301 4672 16313 4675
rect 15896 4644 16313 4672
rect 15896 4632 15902 4644
rect 16301 4641 16313 4644
rect 16347 4672 16359 4675
rect 18322 4672 18328 4684
rect 16347 4644 18328 4672
rect 16347 4641 16359 4644
rect 16301 4635 16359 4641
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 20640 4672 20668 4768
rect 20806 4672 20812 4684
rect 20640 4644 20812 4672
rect 20806 4632 20812 4644
rect 20864 4672 20870 4684
rect 20901 4675 20959 4681
rect 20901 4672 20913 4675
rect 20864 4644 20913 4672
rect 20864 4632 20870 4644
rect 20901 4641 20913 4644
rect 20947 4641 20959 4675
rect 21361 4675 21419 4681
rect 21361 4672 21373 4675
rect 20901 4635 20959 4641
rect 21284 4644 21373 4672
rect 16482 4604 16488 4616
rect 16443 4576 16488 4604
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4604 18843 4607
rect 18966 4604 18972 4616
rect 18831 4576 18972 4604
rect 18831 4573 18843 4576
rect 18785 4567 18843 4573
rect 18966 4564 18972 4576
rect 19024 4604 19030 4616
rect 19426 4604 19432 4616
rect 19024 4576 19432 4604
rect 19024 4564 19030 4576
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 20622 4564 20628 4616
rect 20680 4604 20686 4616
rect 21284 4604 21312 4644
rect 21361 4641 21373 4644
rect 21407 4641 21419 4675
rect 21361 4635 21419 4641
rect 20680 4576 21312 4604
rect 21637 4607 21695 4613
rect 20680 4564 20686 4576
rect 21637 4573 21649 4607
rect 21683 4604 21695 4607
rect 23566 4604 23572 4616
rect 21683 4576 23572 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 23566 4564 23572 4576
rect 23624 4564 23630 4616
rect 18877 4539 18935 4545
rect 18877 4536 18889 4539
rect 13786 4508 18889 4536
rect 18877 4505 18889 4508
rect 18923 4505 18935 4539
rect 18877 4499 18935 4505
rect 2498 4468 2504 4480
rect 2459 4440 2504 4468
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 3326 4468 3332 4480
rect 2915 4440 3332 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3326 4428 3332 4440
rect 3384 4428 3390 4480
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 18555 4471 18613 4477
rect 18555 4468 18567 4471
rect 18472 4440 18567 4468
rect 18472 4428 18478 4440
rect 18555 4437 18567 4440
rect 18601 4437 18613 4471
rect 18555 4431 18613 4437
rect 18693 4471 18751 4477
rect 18693 4437 18705 4471
rect 18739 4468 18751 4471
rect 18782 4468 18788 4480
rect 18739 4440 18788 4468
rect 18739 4437 18751 4440
rect 18693 4431 18751 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 19334 4428 19340 4480
rect 19392 4468 19398 4480
rect 19429 4471 19487 4477
rect 19429 4468 19441 4471
rect 19392 4440 19441 4468
rect 19392 4428 19398 4440
rect 19429 4437 19441 4440
rect 19475 4437 19487 4471
rect 19429 4431 19487 4437
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 1026 4224 1032 4276
rect 1084 4264 1090 4276
rect 4433 4267 4491 4273
rect 4433 4264 4445 4267
rect 1084 4236 4445 4264
rect 1084 4224 1090 4236
rect 4433 4233 4445 4236
rect 4479 4264 4491 4267
rect 10962 4264 10968 4276
rect 4479 4236 4752 4264
rect 10923 4236 10968 4264
rect 4479 4233 4491 4236
rect 4433 4227 4491 4233
rect 1762 4156 1768 4208
rect 1820 4196 1826 4208
rect 2777 4199 2835 4205
rect 2777 4196 2789 4199
rect 1820 4168 2789 4196
rect 1820 4156 1826 4168
rect 2777 4165 2789 4168
rect 2823 4196 2835 4199
rect 2869 4199 2927 4205
rect 2869 4196 2881 4199
rect 2823 4168 2881 4196
rect 2823 4165 2835 4168
rect 2777 4159 2835 4165
rect 2869 4165 2881 4168
rect 2915 4165 2927 4199
rect 2869 4159 2927 4165
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 2222 4128 2228 4140
rect 1627 4100 2228 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 2222 4088 2228 4100
rect 2280 4128 2286 4140
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2280 4100 3065 4128
rect 2280 4088 2286 4100
rect 3053 4097 3065 4100
rect 3099 4128 3111 4131
rect 3326 4128 3332 4140
rect 3099 4100 3332 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 3476 4100 4629 4128
rect 3476 4088 3482 4100
rect 4617 4097 4629 4100
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 1486 4060 1492 4072
rect 1447 4032 1492 4060
rect 1486 4020 1492 4032
rect 1544 4020 1550 4072
rect 1765 4063 1823 4069
rect 1765 4029 1777 4063
rect 1811 4060 1823 4063
rect 2498 4060 2504 4072
rect 1811 4032 2504 4060
rect 1811 4029 1823 4032
rect 1765 4023 1823 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 4724 4069 4752 4236
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 12618 4264 12624 4276
rect 12579 4236 12624 4264
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 15838 4264 15844 4276
rect 15799 4236 15844 4264
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16298 4264 16304 4276
rect 16259 4236 16304 4264
rect 16298 4224 16304 4236
rect 16356 4224 16362 4276
rect 17862 4264 17868 4276
rect 17823 4236 17868 4264
rect 17862 4224 17868 4236
rect 17920 4224 17926 4276
rect 18509 4267 18567 4273
rect 18509 4233 18521 4267
rect 18555 4264 18567 4267
rect 18782 4264 18788 4276
rect 18555 4236 18788 4264
rect 18555 4233 18567 4236
rect 18509 4227 18567 4233
rect 18782 4224 18788 4236
rect 18840 4264 18846 4276
rect 18877 4267 18935 4273
rect 18877 4264 18889 4267
rect 18840 4236 18889 4264
rect 18840 4224 18846 4236
rect 18877 4233 18889 4236
rect 18923 4233 18935 4267
rect 18877 4227 18935 4233
rect 16316 4128 16344 4224
rect 19334 4156 19340 4208
rect 19392 4196 19398 4208
rect 19702 4196 19708 4208
rect 19392 4168 19437 4196
rect 19663 4168 19708 4196
rect 19392 4156 19398 4168
rect 19702 4156 19708 4168
rect 19760 4156 19766 4208
rect 19429 4131 19487 4137
rect 16316 4100 16528 4128
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 3145 4063 3203 4069
rect 3145 4060 3157 4063
rect 2823 4032 3157 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 3145 4029 3157 4032
rect 3191 4029 3203 4063
rect 3145 4023 3203 4029
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 5684 4032 9229 4060
rect 5684 4020 5690 4032
rect 9217 4029 9229 4032
rect 9263 4060 9275 4063
rect 9309 4063 9367 4069
rect 9309 4060 9321 4063
rect 9263 4032 9321 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9309 4029 9321 4032
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9456 4032 9781 4060
rect 9456 4020 9462 4032
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11422 4060 11428 4072
rect 11379 4032 11428 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11422 4020 11428 4032
rect 11480 4060 11486 4072
rect 16500 4069 16528 4100
rect 19429 4097 19441 4131
rect 19475 4128 19487 4131
rect 19610 4128 19616 4140
rect 19475 4100 19616 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 20824 4100 21833 4128
rect 20824 4072 20852 4100
rect 21821 4097 21833 4100
rect 21867 4128 21879 4131
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 21867 4100 22201 4128
rect 21867 4097 21879 4100
rect 21821 4091 21879 4097
rect 22189 4097 22201 4100
rect 22235 4097 22247 4131
rect 22189 4091 22247 4097
rect 16485 4063 16543 4069
rect 11480 4032 16344 4060
rect 11480 4020 11486 4032
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 10042 3992 10048 4004
rect 2271 3964 4108 3992
rect 10003 3964 10048 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 4080 3936 4108 3964
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 1486 3884 1492 3936
rect 1544 3924 1550 3936
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 1544 3896 2513 3924
rect 1544 3884 1550 3896
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 5442 3924 5448 3936
rect 4120 3896 5448 3924
rect 4120 3884 4126 3896
rect 5442 3884 5448 3896
rect 5500 3924 5506 3936
rect 10962 3924 10968 3936
rect 5500 3896 10968 3924
rect 5500 3884 5506 3896
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12584 3896 13093 3924
rect 12584 3884 12590 3896
rect 13081 3893 13093 3896
rect 13127 3924 13139 3927
rect 15470 3924 15476 3936
rect 13127 3896 15476 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 16316 3924 16344 4032
rect 16485 4029 16497 4063
rect 16531 4029 16543 4063
rect 19208 4063 19266 4069
rect 19208 4060 19220 4063
rect 16485 4023 16543 4029
rect 18984 4032 19220 4060
rect 18984 4004 19012 4032
rect 19208 4029 19220 4032
rect 19254 4029 19266 4063
rect 20806 4060 20812 4072
rect 20767 4032 20812 4060
rect 19208 4023 19266 4029
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4029 21327 4063
rect 21269 4023 21327 4029
rect 17129 3995 17187 4001
rect 17129 3961 17141 3995
rect 17175 3992 17187 3995
rect 17402 3992 17408 4004
rect 17175 3964 17408 3992
rect 17175 3961 17187 3964
rect 17129 3955 17187 3961
rect 17402 3952 17408 3964
rect 17460 3992 17466 4004
rect 18966 3992 18972 4004
rect 17460 3964 18972 3992
rect 17460 3952 17466 3964
rect 18966 3952 18972 3964
rect 19024 3952 19030 4004
rect 19061 3995 19119 4001
rect 19061 3961 19073 3995
rect 19107 3992 19119 3995
rect 20162 3992 20168 4004
rect 19107 3964 20168 3992
rect 19107 3961 19119 3964
rect 19061 3955 19119 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 21284 3992 21312 4023
rect 21542 3992 21548 4004
rect 20272 3964 21312 3992
rect 21503 3964 21548 3992
rect 20272 3936 20300 3964
rect 21542 3952 21548 3964
rect 21600 3952 21606 4004
rect 19702 3924 19708 3936
rect 16316 3896 19708 3924
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 20254 3924 20260 3936
rect 20215 3896 20260 3924
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20622 3924 20628 3936
rect 20583 3896 20628 3924
rect 20622 3884 20628 3896
rect 20680 3884 20686 3936
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 106 3680 112 3732
rect 164 3720 170 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 164 3692 4169 3720
rect 164 3680 170 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 4157 3683 4215 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 19610 3720 19616 3732
rect 19571 3692 19616 3720
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 1578 3652 1584 3664
rect 1539 3624 1584 3652
rect 1578 3612 1584 3624
rect 1636 3612 1642 3664
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 19981 3655 20039 3661
rect 19981 3652 19993 3655
rect 19484 3624 19993 3652
rect 19484 3612 19490 3624
rect 19981 3621 19993 3624
rect 20027 3621 20039 3655
rect 19981 3615 20039 3621
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 20772 3624 21404 3652
rect 20772 3612 20778 3624
rect 2130 3584 2136 3596
rect 2043 3556 2136 3584
rect 2130 3544 2136 3556
rect 2188 3544 2194 3596
rect 2222 3544 2228 3596
rect 2280 3584 2286 3596
rect 2409 3587 2467 3593
rect 2280 3556 2325 3584
rect 2280 3544 2286 3556
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 2498 3584 2504 3596
rect 2455 3556 2504 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3584 3939 3587
rect 4062 3584 4068 3596
rect 3927 3556 4068 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4304 3556 4537 3584
rect 4304 3544 4310 3556
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 16758 3544 16764 3596
rect 16816 3584 16822 3596
rect 17037 3587 17095 3593
rect 17037 3584 17049 3587
rect 16816 3556 17049 3584
rect 16816 3544 16822 3556
rect 17037 3553 17049 3556
rect 17083 3584 17095 3587
rect 17310 3584 17316 3596
rect 17083 3556 17316 3584
rect 17083 3553 17095 3556
rect 17037 3547 17095 3553
rect 17310 3544 17316 3556
rect 17368 3584 17374 3596
rect 18601 3587 18659 3593
rect 18601 3584 18613 3587
rect 17368 3556 18613 3584
rect 17368 3544 17374 3556
rect 18601 3553 18613 3556
rect 18647 3584 18659 3587
rect 19334 3584 19340 3596
rect 18647 3556 19340 3584
rect 18647 3553 18659 3556
rect 18601 3547 18659 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 21376 3593 21404 3624
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 20864 3556 20913 3584
rect 20864 3544 20870 3556
rect 20901 3553 20913 3556
rect 20947 3553 20959 3587
rect 20901 3547 20959 3553
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3584 21419 3587
rect 21450 3584 21456 3596
rect 21407 3556 21456 3584
rect 21407 3553 21419 3556
rect 21361 3547 21419 3553
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 2148 3448 2176 3544
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 2958 3516 2964 3528
rect 2915 3488 2964 3516
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 17402 3516 17408 3528
rect 17363 3488 17408 3516
rect 17402 3476 17408 3488
rect 17460 3516 17466 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 17460 3488 18061 3516
rect 17460 3476 17466 3488
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18969 3519 19027 3525
rect 18969 3485 18981 3519
rect 19015 3516 19027 3519
rect 19058 3516 19064 3528
rect 19015 3488 19064 3516
rect 19015 3485 19027 3488
rect 18969 3479 19027 3485
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3516 21695 3519
rect 22830 3516 22836 3528
rect 21683 3488 22836 3516
rect 21683 3485 21695 3488
rect 21637 3479 21695 3485
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 18414 3448 18420 3460
rect 2148 3420 3280 3448
rect 3252 3392 3280 3420
rect 17236 3420 18420 3448
rect 17236 3392 17264 3420
rect 18414 3408 18420 3420
rect 18472 3448 18478 3460
rect 18739 3451 18797 3457
rect 18739 3448 18751 3451
rect 18472 3420 18751 3448
rect 18472 3408 18478 3420
rect 18739 3417 18751 3420
rect 18785 3417 18797 3451
rect 18874 3448 18880 3460
rect 18835 3420 18880 3448
rect 18739 3411 18797 3417
rect 18874 3408 18880 3420
rect 18932 3408 18938 3460
rect 1486 3340 1492 3392
rect 1544 3380 1550 3392
rect 1949 3383 2007 3389
rect 1949 3380 1961 3383
rect 1544 3352 1961 3380
rect 1544 3340 1550 3352
rect 1949 3349 1961 3352
rect 1995 3349 2007 3383
rect 3234 3380 3240 3392
rect 3195 3352 3240 3380
rect 1949 3343 2007 3349
rect 3234 3340 3240 3352
rect 3292 3340 3298 3392
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 17218 3389 17224 3392
rect 17175 3383 17224 3389
rect 17175 3380 17187 3383
rect 16448 3352 17187 3380
rect 16448 3340 16454 3352
rect 17175 3349 17187 3352
rect 17221 3349 17224 3383
rect 17175 3343 17224 3349
rect 17218 3340 17224 3343
rect 17276 3340 17282 3392
rect 17310 3340 17316 3392
rect 17368 3380 17374 3392
rect 17494 3380 17500 3392
rect 17368 3352 17413 3380
rect 17455 3352 17500 3380
rect 17368 3340 17374 3352
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 19058 3380 19064 3392
rect 19019 3352 19064 3380
rect 19058 3340 19064 3352
rect 19116 3380 19122 3392
rect 20254 3380 20260 3392
rect 19116 3352 20260 3380
rect 19116 3340 19122 3352
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3176 2562 3188
rect 2866 3176 2872 3188
rect 2556 3148 2872 3176
rect 2556 3136 2562 3148
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3326 3176 3332 3188
rect 3287 3148 3332 3176
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 5626 3176 5632 3188
rect 5587 3148 5632 3176
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 16758 3176 16764 3188
rect 16719 3148 16764 3176
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17276 3148 17417 3176
rect 17276 3136 17282 3148
rect 17405 3145 17417 3148
rect 17451 3176 17463 3179
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17451 3148 17785 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 18325 3179 18383 3185
rect 18325 3145 18337 3179
rect 18371 3176 18383 3179
rect 18782 3176 18788 3188
rect 18371 3148 18788 3176
rect 18371 3145 18383 3148
rect 18325 3139 18383 3145
rect 1578 3108 1584 3120
rect 1539 3080 1584 3108
rect 1578 3068 1584 3080
rect 1636 3068 1642 3120
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1912 3012 1961 3040
rect 1912 3000 1918 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 5644 3040 5672 3136
rect 17129 3111 17187 3117
rect 17129 3077 17141 3111
rect 17175 3108 17187 3111
rect 17310 3108 17316 3120
rect 17175 3080 17316 3108
rect 17175 3077 17187 3080
rect 17129 3071 17187 3077
rect 17310 3068 17316 3080
rect 17368 3108 17374 3120
rect 18340 3108 18368 3139
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 21450 3136 21456 3188
rect 21508 3176 21514 3188
rect 21545 3179 21603 3185
rect 21545 3176 21557 3179
rect 21508 3148 21557 3176
rect 21508 3136 21514 3148
rect 21545 3145 21557 3148
rect 21591 3145 21603 3179
rect 21545 3139 21603 3145
rect 17368 3080 18368 3108
rect 18693 3111 18751 3117
rect 17368 3068 17374 3080
rect 18693 3077 18705 3111
rect 18739 3108 18751 3111
rect 18966 3108 18972 3120
rect 18739 3080 18972 3108
rect 18739 3077 18751 3080
rect 18693 3071 18751 3077
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 20070 3040 20076 3052
rect 4212 3012 4257 3040
rect 4816 3012 5672 3040
rect 19444 3012 20076 3040
rect 4212 3000 4218 3012
rect 1486 2972 1492 2984
rect 1447 2944 1492 2972
rect 1486 2932 1492 2944
rect 1544 2932 1550 2984
rect 1762 2972 1768 2984
rect 1675 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2972 1826 2984
rect 2498 2972 2504 2984
rect 1820 2944 2504 2972
rect 1820 2932 1826 2944
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 4816 2981 4844 3012
rect 19444 2984 19472 3012
rect 20070 3000 20076 3012
rect 20128 3040 20134 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 20128 3012 20361 3040
rect 20128 3000 20134 3012
rect 20349 3009 20361 3012
rect 20395 3040 20407 3043
rect 20395 3012 21036 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2941 4859 2975
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 4801 2935 4859 2941
rect 2038 2864 2044 2916
rect 2096 2904 2102 2916
rect 4816 2904 4844 2935
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 19242 2972 19248 2984
rect 19203 2944 19248 2972
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 19426 2972 19432 2984
rect 19387 2944 19432 2972
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 19705 2975 19763 2981
rect 19705 2941 19717 2975
rect 19751 2972 19763 2975
rect 19978 2972 19984 2984
rect 19751 2944 19984 2972
rect 19751 2941 19763 2944
rect 19705 2935 19763 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 21008 2981 21036 3012
rect 20809 2975 20867 2981
rect 20809 2941 20821 2975
rect 20855 2941 20867 2975
rect 20809 2935 20867 2941
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 2096 2876 4844 2904
rect 5261 2907 5319 2913
rect 2096 2864 2102 2876
rect 5261 2873 5273 2907
rect 5307 2904 5319 2907
rect 5350 2904 5356 2916
rect 5307 2876 5356 2904
rect 5307 2873 5319 2876
rect 5261 2867 5319 2873
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 3786 2836 3792 2848
rect 3747 2808 3792 2836
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 20622 2836 20628 2848
rect 15528 2808 20628 2836
rect 15528 2796 15534 2808
rect 20622 2796 20628 2808
rect 20680 2836 20686 2848
rect 20824 2836 20852 2935
rect 21266 2904 21272 2916
rect 21227 2876 21272 2904
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 21358 2836 21364 2848
rect 20680 2808 21364 2836
rect 20680 2796 20686 2808
rect 21358 2796 21364 2808
rect 21416 2796 21422 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2038 2632 2044 2644
rect 1995 2604 2044 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3234 2632 3240 2644
rect 3195 2604 3240 2632
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 4212 2604 4257 2632
rect 4356 2604 5181 2632
rect 4212 2592 4218 2604
rect 2501 2567 2559 2573
rect 2501 2564 2513 2567
rect 1596 2536 2513 2564
rect 1596 2508 1624 2536
rect 2501 2533 2513 2536
rect 2547 2533 2559 2567
rect 2501 2527 2559 2533
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2465 1547 2499
rect 1489 2459 1547 2465
rect 1504 2428 1532 2459
rect 1578 2456 1584 2508
rect 1636 2496 1642 2508
rect 1762 2496 1768 2508
rect 1636 2468 1681 2496
rect 1723 2468 1768 2496
rect 1636 2456 1642 2468
rect 1762 2456 1768 2468
rect 1820 2456 1826 2508
rect 4356 2505 4384 2604
rect 5169 2601 5181 2604
rect 5215 2632 5227 2635
rect 5442 2632 5448 2644
rect 5215 2604 5448 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7006 2632 7012 2644
rect 6967 2604 7012 2632
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7374 2592 7380 2644
rect 7432 2592 7438 2644
rect 17129 2635 17187 2641
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 17402 2632 17408 2644
rect 17175 2604 17408 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 18230 2592 18236 2644
rect 18288 2632 18294 2644
rect 18417 2635 18475 2641
rect 18417 2632 18429 2635
rect 18288 2604 18429 2632
rect 18288 2592 18294 2604
rect 18417 2601 18429 2604
rect 18463 2601 18475 2635
rect 18417 2595 18475 2601
rect 19242 2592 19248 2644
rect 19300 2632 19306 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 19300 2604 19717 2632
rect 19300 2592 19306 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 20622 2632 20628 2644
rect 20583 2604 20628 2632
rect 19705 2595 19763 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 5074 2564 5080 2576
rect 4632 2536 5080 2564
rect 4632 2505 4660 2536
rect 5074 2524 5080 2536
rect 5132 2564 5138 2576
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 5132 2536 6745 2564
rect 5132 2524 5138 2536
rect 6733 2533 6745 2536
rect 6779 2564 6791 2567
rect 7392 2564 7420 2592
rect 6779 2536 7420 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 7392 2505 7420 2536
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 19426 2564 19432 2576
rect 18187 2536 19432 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 18800 2505 18828 2536
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2465 4399 2499
rect 4341 2459 4399 2465
rect 4617 2499 4675 2505
rect 4617 2465 4629 2499
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2496 6423 2499
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6411 2468 7205 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17819 2468 18337 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 18785 2499 18843 2505
rect 18785 2465 18797 2499
rect 18831 2465 18843 2499
rect 18785 2459 18843 2465
rect 2130 2428 2136 2440
rect 1504 2400 2136 2428
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 3786 2388 3792 2440
rect 3844 2428 3850 2440
rect 4632 2428 4660 2459
rect 3844 2400 4660 2428
rect 3844 2388 3850 2400
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 6380 2360 6408 2459
rect 7208 2428 7236 2459
rect 7926 2428 7932 2440
rect 7208 2400 7932 2428
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 18340 2428 18368 2459
rect 20806 2428 20812 2440
rect 18340 2400 20812 2428
rect 20806 2388 20812 2400
rect 20864 2428 20870 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20864 2400 20913 2428
rect 20864 2388 20870 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 3016 2332 6408 2360
rect 3016 2320 3022 2332
rect 19426 2292 19432 2304
rect 19387 2264 19432 2292
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
<< via1 >>
rect 848 23196 900 23248
rect 1768 23196 1820 23248
rect 20720 22652 20772 22704
rect 21732 22652 21784 22704
rect 112 22040 164 22092
rect 17960 22040 18012 22092
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 17960 21131 18012 21140
rect 17960 21097 17969 21131
rect 17969 21097 18003 21131
rect 18003 21097 18012 21131
rect 17960 21088 18012 21097
rect 18328 21088 18380 21140
rect 23020 21020 23072 21072
rect 16304 20995 16356 21004
rect 16304 20961 16313 20995
rect 16313 20961 16347 20995
rect 16347 20961 16356 20995
rect 16304 20952 16356 20961
rect 16488 20952 16540 21004
rect 18420 20995 18472 21004
rect 18420 20961 18429 20995
rect 18429 20961 18463 20995
rect 18463 20961 18472 20995
rect 18420 20952 18472 20961
rect 20628 20952 20680 21004
rect 21456 20995 21508 21004
rect 21456 20961 21465 20995
rect 21465 20961 21499 20995
rect 21499 20961 21508 20995
rect 21456 20952 21508 20961
rect 19432 20748 19484 20800
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 112 20544 164 20596
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 8392 20451 8444 20460
rect 8392 20417 8401 20451
rect 8401 20417 8435 20451
rect 8435 20417 8444 20451
rect 8392 20408 8444 20417
rect 1492 20340 1544 20392
rect 4160 20383 4212 20392
rect 4160 20349 4169 20383
rect 4169 20349 4203 20383
rect 4203 20349 4212 20383
rect 4160 20340 4212 20349
rect 4068 20272 4120 20324
rect 4988 20340 5040 20392
rect 8116 20383 8168 20392
rect 8116 20349 8125 20383
rect 8125 20349 8159 20383
rect 8159 20349 8168 20383
rect 8116 20340 8168 20349
rect 8484 20340 8536 20392
rect 11612 20408 11664 20460
rect 13268 20408 13320 20460
rect 8024 20204 8076 20256
rect 10876 20340 10928 20392
rect 12808 20340 12860 20392
rect 18420 20476 18472 20528
rect 20444 20408 20496 20460
rect 21640 20451 21692 20460
rect 21640 20417 21649 20451
rect 21649 20417 21683 20451
rect 21683 20417 21692 20451
rect 21640 20408 21692 20417
rect 15200 20383 15252 20392
rect 15200 20349 15209 20383
rect 15209 20349 15243 20383
rect 15243 20349 15252 20383
rect 15200 20340 15252 20349
rect 19432 20383 19484 20392
rect 16304 20272 16356 20324
rect 19432 20349 19441 20383
rect 19441 20349 19475 20383
rect 19475 20349 19484 20383
rect 19432 20340 19484 20349
rect 20904 20383 20956 20392
rect 20904 20349 20913 20383
rect 20913 20349 20947 20383
rect 20947 20349 20956 20383
rect 20904 20340 20956 20349
rect 21456 20383 21508 20392
rect 21456 20349 21465 20383
rect 21465 20349 21499 20383
rect 21499 20349 21508 20383
rect 21456 20340 21508 20349
rect 13544 20204 13596 20256
rect 14740 20204 14792 20256
rect 16488 20204 16540 20256
rect 18420 20204 18472 20256
rect 18972 20247 19024 20256
rect 18972 20213 18981 20247
rect 18981 20213 19015 20247
rect 19015 20213 19024 20247
rect 18972 20204 19024 20213
rect 20628 20204 20680 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 4160 20000 4212 20052
rect 5632 19932 5684 19984
rect 9496 19932 9548 19984
rect 16672 19975 16724 19984
rect 16672 19941 16681 19975
rect 16681 19941 16715 19975
rect 16715 19941 16724 19975
rect 16672 19932 16724 19941
rect 19248 19975 19300 19984
rect 4804 19907 4856 19916
rect 4804 19873 4813 19907
rect 4813 19873 4847 19907
rect 4847 19873 4856 19907
rect 4804 19864 4856 19873
rect 4988 19907 5040 19916
rect 4988 19873 4997 19907
rect 4997 19873 5031 19907
rect 5031 19873 5040 19907
rect 4988 19864 5040 19873
rect 8024 19907 8076 19916
rect 8024 19873 8033 19907
rect 8033 19873 8067 19907
rect 8067 19873 8076 19907
rect 8024 19864 8076 19873
rect 8484 19907 8536 19916
rect 8484 19873 8493 19907
rect 8493 19873 8527 19907
rect 8527 19873 8536 19907
rect 8484 19864 8536 19873
rect 16212 19907 16264 19916
rect 16212 19873 16221 19907
rect 16221 19873 16255 19907
rect 16255 19873 16264 19907
rect 16212 19864 16264 19873
rect 16488 19907 16540 19916
rect 16488 19873 16497 19907
rect 16497 19873 16531 19907
rect 16531 19873 16540 19907
rect 16488 19864 16540 19873
rect 18512 19907 18564 19916
rect 18512 19873 18521 19907
rect 18521 19873 18555 19907
rect 18555 19873 18564 19907
rect 18512 19864 18564 19873
rect 18972 19907 19024 19916
rect 18972 19873 18981 19907
rect 18981 19873 19015 19907
rect 19015 19873 19024 19907
rect 18972 19864 19024 19873
rect 19248 19941 19257 19975
rect 19257 19941 19291 19975
rect 19291 19941 19300 19975
rect 19248 19932 19300 19941
rect 23572 19932 23624 19984
rect 21272 19864 21324 19916
rect 21456 19907 21508 19916
rect 21456 19873 21465 19907
rect 21465 19873 21499 19907
rect 21499 19873 21508 19907
rect 21456 19864 21508 19873
rect 18328 19796 18380 19848
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 12808 19660 12860 19712
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 8024 19499 8076 19508
rect 8024 19465 8033 19499
rect 8033 19465 8067 19499
rect 8067 19465 8076 19499
rect 8024 19456 8076 19465
rect 21272 19499 21324 19508
rect 21272 19465 21281 19499
rect 21281 19465 21315 19499
rect 21315 19465 21324 19499
rect 21272 19456 21324 19465
rect 21456 19388 21508 19440
rect 16212 19320 16264 19372
rect 19432 19320 19484 19372
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 4068 19184 4120 19236
rect 5448 19184 5500 19236
rect 13544 19184 13596 19236
rect 18512 19252 18564 19304
rect 19340 19295 19392 19304
rect 19340 19261 19349 19295
rect 19349 19261 19383 19295
rect 19383 19261 19392 19295
rect 19340 19252 19392 19261
rect 16488 19184 16540 19236
rect 18144 19184 18196 19236
rect 4804 19116 4856 19168
rect 5816 19116 5868 19168
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 9312 19116 9364 19168
rect 18328 19116 18380 19168
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 23572 18844 23624 18896
rect 1492 18819 1544 18828
rect 1492 18785 1501 18819
rect 1501 18785 1535 18819
rect 1535 18785 1544 18819
rect 1492 18776 1544 18785
rect 1676 18776 1728 18828
rect 19984 18776 20036 18828
rect 20628 18776 20680 18828
rect 21364 18819 21416 18828
rect 21364 18785 21373 18819
rect 21373 18785 21407 18819
rect 21407 18785 21416 18819
rect 21364 18776 21416 18785
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 18972 18708 19024 18760
rect 18144 18640 18196 18692
rect 19340 18640 19392 18692
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 1492 18368 1544 18420
rect 19432 18164 19484 18216
rect 20812 18164 20864 18216
rect 21364 18207 21416 18216
rect 21364 18173 21373 18207
rect 21373 18173 21407 18207
rect 21407 18173 21416 18207
rect 21364 18164 21416 18173
rect 21640 18207 21692 18216
rect 21640 18173 21649 18207
rect 21649 18173 21683 18207
rect 21683 18173 21692 18207
rect 21640 18164 21692 18173
rect 17868 18096 17920 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 14740 18028 14792 18080
rect 19984 18071 20036 18080
rect 19984 18037 19993 18071
rect 19993 18037 20027 18071
rect 20027 18037 20036 18071
rect 19984 18028 20036 18037
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 1584 17824 1636 17876
rect 8116 17824 8168 17876
rect 20812 17484 20864 17536
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 1676 17076 1728 17128
rect 112 16940 164 16992
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 19524 16736 19576 16788
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 15384 16099 15436 16108
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 15384 16065 15393 16099
rect 15393 16065 15427 16099
rect 15427 16065 15436 16099
rect 15384 16056 15436 16065
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 19248 15988 19300 16040
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 19156 15895 19208 15904
rect 19156 15861 19165 15895
rect 19165 15861 19199 15895
rect 19199 15861 19208 15895
rect 19156 15852 19208 15861
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 1400 15648 1452 15700
rect 1952 15555 2004 15564
rect 1952 15521 1961 15555
rect 1961 15521 1995 15555
rect 1995 15521 2004 15555
rect 1952 15512 2004 15521
rect 19524 15580 19576 15632
rect 23572 15580 23624 15632
rect 19340 15512 19392 15564
rect 2044 15444 2096 15496
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 18880 15104 18932 15156
rect 19248 15147 19300 15156
rect 19248 15113 19257 15147
rect 19257 15113 19291 15147
rect 19291 15113 19300 15147
rect 19248 15104 19300 15113
rect 19524 15104 19576 15156
rect 11888 14968 11940 15020
rect 13544 14968 13596 15020
rect 14188 15011 14240 15020
rect 1952 14900 2004 14952
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 12440 14764 12492 14816
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 19524 13880 19576 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 12440 13812 12492 13864
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 23572 13880 23624 13932
rect 20444 13812 20496 13864
rect 112 13676 164 13728
rect 19892 13676 19944 13728
rect 20444 13676 20496 13728
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 1952 13472 2004 13524
rect 19892 13515 19944 13524
rect 19892 13481 19901 13515
rect 19901 13481 19935 13515
rect 19935 13481 19944 13515
rect 19892 13472 19944 13481
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 5816 12928 5868 12980
rect 18972 12928 19024 12980
rect 11152 12792 11204 12844
rect 14740 12792 14792 12844
rect 10784 12767 10836 12776
rect 10784 12733 10793 12767
rect 10793 12733 10827 12767
rect 10827 12733 10836 12767
rect 10784 12724 10836 12733
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 19524 12767 19576 12776
rect 19524 12733 19533 12767
rect 19533 12733 19567 12767
rect 19567 12733 19576 12767
rect 19524 12724 19576 12733
rect 19616 12724 19668 12776
rect 10324 12631 10376 12640
rect 10324 12597 10333 12631
rect 10333 12597 10367 12631
rect 10367 12597 10376 12631
rect 10324 12588 10376 12597
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 19616 12427 19668 12436
rect 1308 12316 1360 12368
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 2044 12316 2096 12368
rect 23572 12316 23624 12368
rect 1952 12291 2004 12300
rect 1952 12257 1961 12291
rect 1961 12257 1995 12291
rect 1995 12257 2004 12291
rect 1952 12248 2004 12257
rect 20812 12248 20864 12300
rect 21272 12248 21324 12300
rect 10784 12044 10836 12096
rect 11428 12044 11480 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 20812 11840 20864 11892
rect 1952 11636 2004 11688
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 19524 10752 19576 10804
rect 1584 10591 1636 10600
rect 1584 10557 1593 10591
rect 1593 10557 1627 10591
rect 1627 10557 1636 10591
rect 1584 10548 1636 10557
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 20628 10548 20680 10600
rect 21640 10659 21692 10668
rect 21640 10625 21649 10659
rect 21649 10625 21683 10659
rect 21683 10625 21692 10659
rect 21640 10616 21692 10625
rect 112 10412 164 10464
rect 19708 10412 19760 10464
rect 21272 10480 21324 10532
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 1952 10208 2004 10260
rect 21272 10072 21324 10124
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 23572 10072 23624 10124
rect 10876 9868 10928 9920
rect 13728 9868 13780 9920
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 13728 9528 13780 9580
rect 19616 9528 19668 9580
rect 20812 9503 20864 9512
rect 20812 9469 20821 9503
rect 20821 9469 20855 9503
rect 20855 9469 20864 9503
rect 20812 9460 20864 9469
rect 19432 9392 19484 9444
rect 19524 9392 19576 9444
rect 18236 9324 18288 9376
rect 20720 9324 20772 9376
rect 21364 9324 21416 9376
rect 112 9188 164 9240
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 17868 9120 17920 9172
rect 17776 9052 17828 9104
rect 18696 9052 18748 9104
rect 1952 9027 2004 9036
rect 1952 8993 1961 9027
rect 1961 8993 1995 9027
rect 1995 8993 2004 9027
rect 1952 8984 2004 8993
rect 6552 9027 6604 9036
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 18604 8984 18656 9036
rect 1676 8916 1728 8968
rect 18512 8916 18564 8968
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 18972 8916 19024 8968
rect 20812 8848 20864 8900
rect 18236 8780 18288 8832
rect 20720 8780 20772 8832
rect 21456 8780 21508 8832
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 2596 8576 2648 8628
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 18420 8576 18472 8628
rect 18236 8304 18288 8356
rect 18512 8440 18564 8492
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 18604 8415 18656 8424
rect 18604 8381 18613 8415
rect 18613 8381 18647 8415
rect 18647 8381 18656 8415
rect 18604 8372 18656 8381
rect 19064 8372 19116 8424
rect 7104 8279 7156 8288
rect 7104 8245 7113 8279
rect 7113 8245 7147 8279
rect 7147 8245 7156 8279
rect 7104 8236 7156 8245
rect 7840 8236 7892 8288
rect 19432 8236 19484 8288
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 18604 8032 18656 8084
rect 18880 8032 18932 8084
rect 23572 7964 23624 8016
rect 20812 7896 20864 7948
rect 21456 7939 21508 7948
rect 18972 7828 19024 7880
rect 21456 7905 21465 7939
rect 21465 7905 21499 7939
rect 21499 7905 21508 7939
rect 21456 7896 21508 7905
rect 21732 7828 21784 7880
rect 18696 7803 18748 7812
rect 18696 7769 18705 7803
rect 18705 7769 18739 7803
rect 18739 7769 18748 7803
rect 18696 7760 18748 7769
rect 19064 7760 19116 7812
rect 17500 7692 17552 7744
rect 18236 7692 18288 7744
rect 19340 7692 19392 7744
rect 20352 7735 20404 7744
rect 20352 7701 20361 7735
rect 20361 7701 20395 7735
rect 20395 7701 20404 7735
rect 20352 7692 20404 7701
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 18420 7488 18472 7540
rect 18696 7488 18748 7540
rect 19616 7488 19668 7540
rect 20168 7488 20220 7540
rect 17316 7420 17368 7472
rect 18972 7420 19024 7472
rect 19340 7420 19392 7472
rect 1584 7352 1636 7404
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 19432 7352 19484 7404
rect 19616 7352 19668 7404
rect 20352 7420 20404 7472
rect 18236 7284 18288 7336
rect 20260 7284 20312 7336
rect 20720 7327 20772 7336
rect 20720 7293 20734 7327
rect 20734 7293 20772 7327
rect 20720 7284 20772 7293
rect 18512 7216 18564 7268
rect 21732 7259 21784 7268
rect 21732 7225 21741 7259
rect 21741 7225 21775 7259
rect 21775 7225 21784 7259
rect 21732 7216 21784 7225
rect 112 7148 164 7200
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 21456 7148 21508 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 18144 6944 18196 6996
rect 19248 6944 19300 6996
rect 19616 6944 19668 6996
rect 20352 6944 20404 6996
rect 18604 6876 18656 6928
rect 23572 6876 23624 6928
rect 16488 6808 16540 6860
rect 17316 6808 17368 6860
rect 18972 6808 19024 6860
rect 20536 6808 20588 6860
rect 21456 6851 21508 6860
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 17224 6740 17276 6792
rect 19432 6740 19484 6792
rect 21456 6817 21465 6851
rect 21465 6817 21499 6851
rect 21499 6817 21508 6851
rect 21456 6808 21508 6817
rect 22284 6740 22336 6792
rect 16488 6647 16540 6656
rect 16488 6613 16497 6647
rect 16497 6613 16531 6647
rect 16531 6613 16540 6647
rect 16488 6604 16540 6613
rect 16672 6604 16724 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 17500 6604 17552 6656
rect 19340 6672 19392 6724
rect 18236 6604 18288 6656
rect 19616 6604 19668 6656
rect 20536 6604 20588 6656
rect 20720 6604 20772 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 1584 6400 1636 6452
rect 1860 6400 1912 6452
rect 10876 6400 10928 6452
rect 16764 6400 16816 6452
rect 16948 6400 17000 6452
rect 17132 6400 17184 6452
rect 21272 6400 21324 6452
rect 22284 6443 22336 6452
rect 22284 6409 22293 6443
rect 22293 6409 22327 6443
rect 22327 6409 22336 6443
rect 22284 6400 22336 6409
rect 17316 6332 17368 6384
rect 19340 6375 19392 6384
rect 19340 6341 19349 6375
rect 19349 6341 19383 6375
rect 19383 6341 19392 6375
rect 19340 6332 19392 6341
rect 17224 6264 17276 6316
rect 19432 6307 19484 6316
rect 19432 6273 19441 6307
rect 19441 6273 19475 6307
rect 19475 6273 19484 6307
rect 19432 6264 19484 6273
rect 20352 6264 20404 6316
rect 7840 6196 7892 6248
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 11244 6239 11296 6248
rect 11244 6205 11253 6239
rect 11253 6205 11287 6239
rect 11287 6205 11296 6239
rect 11244 6196 11296 6205
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 8484 6171 8536 6180
rect 8484 6137 8493 6171
rect 8493 6137 8527 6171
rect 8527 6137 8536 6171
rect 8484 6128 8536 6137
rect 16672 6196 16724 6248
rect 17960 6196 18012 6248
rect 18604 6196 18656 6248
rect 19248 6239 19300 6248
rect 19248 6205 19254 6239
rect 19254 6205 19300 6239
rect 19248 6196 19300 6205
rect 20720 6196 20772 6248
rect 18236 6171 18288 6180
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 16304 6103 16356 6112
rect 16304 6069 16313 6103
rect 16313 6069 16347 6103
rect 16347 6069 16356 6103
rect 18236 6137 18245 6171
rect 18245 6137 18279 6171
rect 18279 6137 18288 6171
rect 18236 6128 18288 6137
rect 21272 6196 21324 6248
rect 21640 6239 21692 6248
rect 21640 6205 21649 6239
rect 21649 6205 21683 6239
rect 21683 6205 21692 6239
rect 21640 6196 21692 6205
rect 16304 6060 16356 6069
rect 16856 6060 16908 6112
rect 18696 6060 18748 6112
rect 21732 6128 21784 6180
rect 20536 6060 20588 6112
rect 20996 6060 21048 6112
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 2044 5856 2096 5908
rect 7932 5856 7984 5908
rect 11244 5856 11296 5908
rect 15384 5899 15436 5908
rect 15384 5865 15393 5899
rect 15393 5865 15427 5899
rect 15427 5865 15436 5899
rect 15384 5856 15436 5865
rect 16856 5856 16908 5908
rect 21456 5856 21508 5908
rect 21548 5899 21600 5908
rect 21548 5865 21557 5899
rect 21557 5865 21591 5899
rect 21591 5865 21600 5899
rect 21548 5856 21600 5865
rect 2596 5763 2648 5772
rect 2596 5729 2605 5763
rect 2605 5729 2639 5763
rect 2639 5729 2648 5763
rect 2596 5720 2648 5729
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 15476 5720 15528 5772
rect 18144 5788 18196 5840
rect 18420 5788 18472 5840
rect 19524 5831 19576 5840
rect 19524 5797 19533 5831
rect 19533 5797 19567 5831
rect 19567 5797 19576 5831
rect 19524 5788 19576 5797
rect 20076 5788 20128 5840
rect 17316 5763 17368 5772
rect 17316 5729 17325 5763
rect 17325 5729 17359 5763
rect 17359 5729 17368 5763
rect 17316 5720 17368 5729
rect 17960 5763 18012 5772
rect 17960 5729 17969 5763
rect 17969 5729 18003 5763
rect 18003 5729 18012 5763
rect 17960 5720 18012 5729
rect 18512 5720 18564 5772
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 19432 5652 19484 5704
rect 18420 5584 18472 5636
rect 18788 5584 18840 5636
rect 20996 5652 21048 5704
rect 22284 5652 22336 5704
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 11244 5516 11296 5568
rect 12532 5516 12584 5568
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 16488 5516 16540 5568
rect 17316 5516 17368 5568
rect 18696 5516 18748 5568
rect 19340 5516 19392 5568
rect 20812 5516 20864 5568
rect 21456 5516 21508 5568
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 2596 5312 2648 5364
rect 2964 5312 3016 5364
rect 15476 5312 15528 5364
rect 16764 5355 16816 5364
rect 16764 5321 16773 5355
rect 16773 5321 16807 5355
rect 16807 5321 16816 5355
rect 16764 5312 16816 5321
rect 18328 5312 18380 5364
rect 22284 5355 22336 5364
rect 22284 5321 22293 5355
rect 22293 5321 22327 5355
rect 22327 5321 22336 5355
rect 22284 5312 22336 5321
rect 18696 5244 18748 5296
rect 18788 5287 18840 5296
rect 18788 5253 18797 5287
rect 18797 5253 18831 5287
rect 18831 5253 18840 5287
rect 18788 5244 18840 5253
rect 20168 5244 20220 5296
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 16304 5176 16356 5228
rect 18972 5176 19024 5228
rect 20812 5176 20864 5228
rect 2780 5108 2832 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 4160 5040 4212 5092
rect 15292 5040 15344 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 18696 5040 18748 5092
rect 19616 5108 19668 5160
rect 20628 5108 20680 5160
rect 21272 5108 21324 5160
rect 21640 5151 21692 5160
rect 21640 5117 21649 5151
rect 21649 5117 21683 5151
rect 21683 5117 21692 5151
rect 21640 5108 21692 5117
rect 19156 4972 19208 5024
rect 19340 4972 19392 5024
rect 20260 4972 20312 5024
rect 21456 4972 21508 5024
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 17868 4768 17920 4820
rect 1584 4675 1636 4684
rect 1584 4641 1593 4675
rect 1593 4641 1627 4675
rect 1627 4641 1636 4675
rect 1584 4632 1636 4641
rect 10968 4632 11020 4684
rect 15292 4700 15344 4752
rect 18512 4768 18564 4820
rect 19432 4768 19484 4820
rect 20628 4811 20680 4820
rect 20628 4777 20637 4811
rect 20637 4777 20671 4811
rect 20671 4777 20680 4811
rect 20628 4768 20680 4777
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 12624 4632 12676 4684
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 15476 4632 15528 4684
rect 15844 4632 15896 4684
rect 18328 4632 18380 4684
rect 20812 4632 20864 4684
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 18972 4564 19024 4616
rect 19432 4564 19484 4616
rect 20628 4564 20680 4616
rect 23572 4564 23624 4616
rect 2504 4471 2556 4480
rect 2504 4437 2513 4471
rect 2513 4437 2547 4471
rect 2547 4437 2556 4471
rect 2504 4428 2556 4437
rect 3332 4428 3384 4480
rect 18420 4428 18472 4480
rect 18788 4428 18840 4480
rect 19340 4428 19392 4480
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 1032 4224 1084 4276
rect 10968 4267 11020 4276
rect 1768 4156 1820 4208
rect 2228 4088 2280 4140
rect 3332 4088 3384 4140
rect 3424 4088 3476 4140
rect 1492 4063 1544 4072
rect 1492 4029 1501 4063
rect 1501 4029 1535 4063
rect 1535 4029 1544 4063
rect 1492 4020 1544 4029
rect 2504 4020 2556 4072
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 12624 4267 12676 4276
rect 12624 4233 12633 4267
rect 12633 4233 12667 4267
rect 12667 4233 12676 4267
rect 12624 4224 12676 4233
rect 15844 4267 15896 4276
rect 15844 4233 15853 4267
rect 15853 4233 15887 4267
rect 15887 4233 15896 4267
rect 15844 4224 15896 4233
rect 16304 4267 16356 4276
rect 16304 4233 16313 4267
rect 16313 4233 16347 4267
rect 16347 4233 16356 4267
rect 16304 4224 16356 4233
rect 17868 4267 17920 4276
rect 17868 4233 17877 4267
rect 17877 4233 17911 4267
rect 17911 4233 17920 4267
rect 17868 4224 17920 4233
rect 18788 4224 18840 4276
rect 19340 4199 19392 4208
rect 19340 4165 19349 4199
rect 19349 4165 19383 4199
rect 19383 4165 19392 4199
rect 19708 4199 19760 4208
rect 19340 4156 19392 4165
rect 19708 4165 19717 4199
rect 19717 4165 19751 4199
rect 19751 4165 19760 4199
rect 19708 4156 19760 4165
rect 5632 4020 5684 4072
rect 9404 4020 9456 4072
rect 11428 4020 11480 4072
rect 19616 4088 19668 4140
rect 10048 3995 10100 4004
rect 10048 3961 10057 3995
rect 10057 3961 10091 3995
rect 10091 3961 10100 3995
rect 10048 3952 10100 3961
rect 1492 3884 1544 3936
rect 4068 3884 4120 3936
rect 5448 3884 5500 3936
rect 10968 3884 11020 3936
rect 12532 3884 12584 3936
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 15476 3884 15528 3893
rect 20812 4063 20864 4072
rect 20812 4029 20821 4063
rect 20821 4029 20855 4063
rect 20855 4029 20864 4063
rect 20812 4020 20864 4029
rect 17408 3952 17460 4004
rect 18972 3952 19024 4004
rect 20168 3952 20220 4004
rect 21548 3995 21600 4004
rect 21548 3961 21557 3995
rect 21557 3961 21591 3995
rect 21591 3961 21600 3995
rect 21548 3952 21600 3961
rect 19708 3884 19760 3936
rect 20260 3927 20312 3936
rect 20260 3893 20269 3927
rect 20269 3893 20303 3927
rect 20303 3893 20312 3927
rect 20260 3884 20312 3893
rect 20628 3927 20680 3936
rect 20628 3893 20637 3927
rect 20637 3893 20671 3927
rect 20671 3893 20680 3927
rect 20628 3884 20680 3893
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 112 3680 164 3732
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 19616 3723 19668 3732
rect 19616 3689 19625 3723
rect 19625 3689 19659 3723
rect 19659 3689 19668 3723
rect 19616 3680 19668 3689
rect 1584 3655 1636 3664
rect 1584 3621 1593 3655
rect 1593 3621 1627 3655
rect 1627 3621 1636 3655
rect 1584 3612 1636 3621
rect 19432 3612 19484 3664
rect 20720 3612 20772 3664
rect 2136 3587 2188 3596
rect 2136 3553 2145 3587
rect 2145 3553 2179 3587
rect 2179 3553 2188 3587
rect 2136 3544 2188 3553
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 2504 3544 2556 3596
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 4252 3544 4304 3596
rect 16764 3544 16816 3596
rect 17316 3544 17368 3596
rect 19340 3544 19392 3596
rect 20812 3544 20864 3596
rect 21456 3544 21508 3596
rect 2964 3476 3016 3528
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 19064 3476 19116 3528
rect 22836 3476 22888 3528
rect 18420 3451 18472 3460
rect 18420 3417 18429 3451
rect 18429 3417 18463 3451
rect 18463 3417 18472 3451
rect 18420 3408 18472 3417
rect 18880 3451 18932 3460
rect 18880 3417 18889 3451
rect 18889 3417 18923 3451
rect 18923 3417 18932 3451
rect 18880 3408 18932 3417
rect 1492 3340 1544 3392
rect 3240 3383 3292 3392
rect 3240 3349 3249 3383
rect 3249 3349 3283 3383
rect 3283 3349 3292 3383
rect 3240 3340 3292 3349
rect 16396 3340 16448 3392
rect 17224 3340 17276 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17500 3383 17552 3392
rect 17316 3340 17368 3349
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 19064 3383 19116 3392
rect 19064 3349 19073 3383
rect 19073 3349 19107 3383
rect 19107 3349 19116 3383
rect 19064 3340 19116 3349
rect 20260 3340 20312 3392
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2872 3179 2924 3188
rect 2504 3136 2556 3145
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 3332 3179 3384 3188
rect 3332 3145 3341 3179
rect 3341 3145 3375 3179
rect 3375 3145 3384 3179
rect 3332 3136 3384 3145
rect 5632 3179 5684 3188
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 17224 3136 17276 3188
rect 1584 3111 1636 3120
rect 1584 3077 1593 3111
rect 1593 3077 1627 3111
rect 1627 3077 1636 3111
rect 1584 3068 1636 3077
rect 1860 3000 1912 3052
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 17316 3068 17368 3120
rect 18788 3136 18840 3188
rect 21456 3136 21508 3188
rect 18972 3068 19024 3120
rect 20076 3043 20128 3052
rect 4160 3000 4212 3009
rect 1492 2975 1544 2984
rect 1492 2941 1501 2975
rect 1501 2941 1535 2975
rect 1535 2941 1544 2975
rect 1492 2932 1544 2941
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2504 2932 2556 2984
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 5080 2975 5132 2984
rect 2044 2864 2096 2916
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 19248 2975 19300 2984
rect 19248 2941 19257 2975
rect 19257 2941 19291 2975
rect 19291 2941 19300 2975
rect 19248 2932 19300 2941
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 19984 2932 20036 2984
rect 5356 2864 5408 2916
rect 3792 2839 3844 2848
rect 3792 2805 3801 2839
rect 3801 2805 3835 2839
rect 3835 2805 3844 2839
rect 3792 2796 3844 2805
rect 15476 2796 15528 2848
rect 20628 2796 20680 2848
rect 21272 2907 21324 2916
rect 21272 2873 21281 2907
rect 21281 2873 21315 2907
rect 21315 2873 21324 2907
rect 21272 2864 21324 2873
rect 21364 2796 21416 2848
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 2044 2592 2096 2644
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3240 2635 3292 2644
rect 3240 2601 3249 2635
rect 3249 2601 3283 2635
rect 3283 2601 3292 2635
rect 3240 2592 3292 2601
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1768 2499 1820 2508
rect 1584 2456 1636 2465
rect 1768 2465 1777 2499
rect 1777 2465 1811 2499
rect 1811 2465 1820 2499
rect 1768 2456 1820 2465
rect 5448 2592 5500 2644
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 7380 2592 7432 2644
rect 17408 2592 17460 2644
rect 18236 2592 18288 2644
rect 19248 2592 19300 2644
rect 20628 2635 20680 2644
rect 20628 2601 20637 2635
rect 20637 2601 20671 2635
rect 20671 2601 20680 2635
rect 20628 2592 20680 2601
rect 5080 2524 5132 2576
rect 19432 2524 19484 2576
rect 2136 2388 2188 2440
rect 3792 2388 3844 2440
rect 2964 2320 3016 2372
rect 7932 2388 7984 2440
rect 20812 2388 20864 2440
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
<< metal2 >>
rect 570 23610 626 24000
rect 1766 23610 1822 24000
rect 3054 23610 3110 24000
rect 570 23582 888 23610
rect 570 23520 626 23582
rect 860 23254 888 23582
rect 1412 23582 1822 23610
rect 848 23248 900 23254
rect 848 23190 900 23196
rect 110 23080 166 23089
rect 110 23015 166 23024
rect 124 22098 152 23015
rect 112 22092 164 22098
rect 112 22034 164 22040
rect 110 21312 166 21321
rect 110 21247 166 21256
rect 124 20602 152 21247
rect 112 20596 164 20602
rect 112 20538 164 20544
rect 1412 18306 1440 23582
rect 1766 23520 1822 23582
rect 2884 23582 3110 23610
rect 1768 23248 1820 23254
rect 1768 23190 1820 23196
rect 1492 20392 1544 20398
rect 1492 20334 1544 20340
rect 1504 18834 1532 20334
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1596 18970 1624 19071
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1492 18828 1544 18834
rect 1492 18770 1544 18776
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1504 18426 1532 18770
rect 1492 18420 1544 18426
rect 1492 18362 1544 18368
rect 1412 18278 1532 18306
rect 110 17912 166 17921
rect 110 17847 166 17856
rect 124 16998 152 17847
rect 112 16992 164 16998
rect 112 16934 164 16940
rect 1398 15872 1454 15881
rect 1398 15807 1454 15816
rect 1412 15706 1440 15807
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 110 14512 166 14521
rect 110 14447 166 14456
rect 124 13734 152 14447
rect 112 13728 164 13734
rect 112 13670 164 13676
rect 1306 12472 1362 12481
rect 1306 12407 1362 12416
rect 1320 12374 1348 12407
rect 1308 12368 1360 12374
rect 1308 12310 1360 12316
rect 110 11112 166 11121
rect 110 11047 166 11056
rect 124 10470 152 11047
rect 112 10464 164 10470
rect 112 10406 164 10412
rect 1504 9489 1532 18278
rect 1688 18086 1716 18770
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1596 17134 1624 17818
rect 1688 17134 1716 18022
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1676 17128 1728 17134
rect 1676 17070 1728 17076
rect 1596 14618 1624 17070
rect 1688 16454 1716 17070
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1688 16017 1716 16390
rect 1674 16008 1730 16017
rect 1674 15943 1730 15952
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1596 13870 1624 14554
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 11354 1624 13806
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1596 10606 1624 11290
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1490 9480 1546 9489
rect 1490 9415 1546 9424
rect 110 9344 166 9353
rect 110 9279 166 9288
rect 124 9246 152 9279
rect 112 9240 164 9246
rect 112 9182 164 9188
rect 1596 8090 1624 10542
rect 1674 9072 1730 9081
rect 1674 9007 1730 9016
rect 1688 8974 1716 9007
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1688 8634 1716 8910
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 110 7712 166 7721
rect 110 7647 166 7656
rect 124 7206 152 7647
rect 1596 7410 1624 8026
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 112 7200 164 7206
rect 112 7142 164 7148
rect 1596 6458 1624 7346
rect 1688 7342 1716 8570
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 7002 1716 7278
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4690 1624 4966
rect 1584 4684 1636 4690
rect 1504 4644 1584 4672
rect 1032 4276 1084 4282
rect 1032 4218 1084 4224
rect 112 3732 164 3738
rect 112 3674 164 3680
rect 124 2553 152 3674
rect 110 2544 166 2553
rect 110 2479 166 2488
rect 754 82 810 480
rect 1044 82 1072 4218
rect 1504 4078 1532 4644
rect 1584 4626 1636 4632
rect 1780 4214 1808 23190
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1964 14958 1992 15506
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 1952 14952 2004 14958
rect 2056 14929 2084 15438
rect 1952 14894 2004 14900
rect 2042 14920 2098 14929
rect 1964 13977 1992 14894
rect 2042 14855 2098 14864
rect 2056 14822 2084 14855
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1950 13968 2006 13977
rect 1950 13903 2006 13912
rect 1964 13870 1992 13903
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13530 1992 13806
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2056 12374 2084 14758
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1964 11694 1992 12242
rect 2056 11898 2084 12310
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 10713 1992 11630
rect 1950 10704 2006 10713
rect 1950 10639 2006 10648
rect 1964 10606 1992 10639
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 10266 1992 10542
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1964 8634 1992 8978
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1768 4208 1820 4214
rect 1768 4154 1820 4156
rect 1596 4150 1820 4154
rect 1596 4126 1808 4150
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3942 1532 4014
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1504 3398 1532 3878
rect 1596 3670 1624 4126
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 2990 1532 3334
rect 1596 3126 1624 3606
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1504 1465 1532 2926
rect 1596 2514 1624 3062
rect 1872 3058 1900 6394
rect 2056 5914 2084 11834
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2044 5908 2096 5914
rect 2096 5868 2176 5896
rect 2044 5850 2096 5856
rect 2148 5166 2176 5868
rect 2608 5778 2636 8570
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2608 5370 2636 5714
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2792 5166 2820 5714
rect 2884 5710 2912 23582
rect 3054 23520 3110 23582
rect 4342 23610 4398 24000
rect 5538 23610 5594 24000
rect 6826 23610 6882 24000
rect 8114 23610 8170 24000
rect 9402 23610 9458 24000
rect 10598 23610 10654 24000
rect 11886 23610 11942 24000
rect 4342 23582 4568 23610
rect 4342 23520 4398 23582
rect 4540 20466 4568 23582
rect 5538 23582 5672 23610
rect 5538 23520 5594 23582
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4080 19242 4108 20266
rect 4172 20058 4200 20334
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 5000 19922 5028 20334
rect 5644 19990 5672 23582
rect 6826 23582 6960 23610
rect 6826 23520 6882 23582
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4816 19174 4844 19858
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 5460 6905 5488 19178
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5828 12986 5856 19110
rect 6932 13814 6960 23582
rect 8114 23582 8432 23610
rect 8114 23520 8170 23582
rect 8404 20466 8432 23582
rect 9402 23582 9536 23610
rect 9402 23520 9458 23582
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 8036 19922 8064 20198
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8036 19514 8064 19858
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 8128 18873 8156 20334
rect 8496 19922 8524 20334
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 9508 19990 9536 23582
rect 10336 23582 10654 23610
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8496 19174 8524 19858
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 8114 18864 8170 18873
rect 8114 18799 8170 18808
rect 8128 17882 8156 18799
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 6840 13786 6960 13814
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 6840 9178 6868 13786
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6564 8634 6592 8978
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 7116 8294 7144 8978
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 5446 6896 5502 6905
rect 5446 6831 5502 6840
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 7852 6254 7880 8230
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 9324 7993 9352 19110
rect 10336 12646 10364 23582
rect 10598 23520 10654 23582
rect 11624 23582 11942 23610
rect 11624 20466 11652 23582
rect 11886 23520 11942 23582
rect 13174 23610 13230 24000
rect 14462 23610 14518 24000
rect 15658 23610 15714 24000
rect 16946 23610 17002 24000
rect 13174 23582 13308 23610
rect 13174 23520 13230 23582
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 13280 20466 13308 23582
rect 14200 23582 14518 23610
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 10888 19718 10916 20334
rect 12820 19718 12848 20334
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10796 12102 10824 12718
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10888 9926 10916 19654
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 13556 19242 13584 20198
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 13556 15026 13584 19178
rect 14200 15026 14228 23582
rect 14462 23520 14518 23582
rect 15396 23582 15714 23610
rect 15198 20496 15254 20505
rect 15198 20431 15254 20440
rect 15212 20398 15240 20431
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14752 18086 14780 20198
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14752 16046 14780 18022
rect 15396 16114 15424 23582
rect 15658 23520 15714 23582
rect 16684 23582 17002 23610
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16316 20330 16344 20946
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 16500 20262 16528 20946
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16500 19922 16528 20198
rect 16684 19990 16712 23582
rect 16946 23520 17002 23582
rect 18234 23610 18290 24000
rect 19522 23610 19578 24000
rect 20718 23610 20774 24000
rect 22006 23610 22062 24000
rect 23294 23610 23350 24000
rect 18234 23582 18368 23610
rect 18234 23520 18290 23582
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 17972 21146 18000 22034
rect 18340 21146 18368 23582
rect 19260 23582 19578 23610
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18432 20534 18460 20946
rect 18420 20528 18472 20534
rect 18420 20470 18472 20476
rect 18432 20262 18460 20470
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16224 19378 16252 19858
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16500 19242 16528 19858
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 18156 18698 18184 19178
rect 18340 19174 18368 19790
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18144 18692 18196 18698
rect 18144 18634 18196 18640
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 14740 16040 14792 16046
rect 17880 16017 17908 18090
rect 14740 15982 14792 15988
rect 17866 16008 17922 16017
rect 14752 15366 14780 15982
rect 17866 15943 17922 15952
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 11900 14929 11928 14962
rect 11886 14920 11942 14929
rect 11886 14855 11942 14864
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 13870 12480 14758
rect 13556 14618 13584 14962
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 12622 13968 12678 13977
rect 12622 13903 12678 13912
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 7852 5574 7880 6190
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2136 5160 2188 5166
rect 2056 5120 2136 5148
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 2514 1808 2926
rect 2056 2922 2084 5120
rect 2136 5102 2188 5108
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 4729 2268 4966
rect 2226 4720 2282 4729
rect 2226 4655 2282 4664
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2148 3602 2176 4558
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2240 3602 2268 4082
rect 2516 4078 2544 4422
rect 2504 4072 2556 4078
rect 2502 4040 2504 4049
rect 2556 4040 2558 4049
rect 2502 3975 2558 3984
rect 2516 3602 2544 3975
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2044 2916 2096 2922
rect 2044 2858 2096 2864
rect 2056 2650 2084 2858
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 2148 2446 2176 3538
rect 2516 3194 2544 3538
rect 2976 3534 3004 5306
rect 7852 5273 7880 5510
rect 7838 5264 7894 5273
rect 7838 5199 7894 5208
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4146 3372 4422
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2516 2990 2544 3130
rect 2594 3088 2650 3097
rect 2594 3023 2650 3032
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 754 54 1072 82
rect 2318 82 2374 480
rect 2608 82 2636 3023
rect 2884 2650 2912 3130
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2976 2378 3004 3470
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3252 2650 3280 3334
rect 3344 3194 3372 4082
rect 3436 4049 3464 4082
rect 3422 4040 3478 4049
rect 3422 3975 3478 3984
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3602 4108 3878
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4172 3584 4200 5034
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 4252 3596 4304 3602
rect 4172 3556 4252 3584
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 4172 3058 4200 3556
rect 4252 3538 4304 3544
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4172 2961 4200 2994
rect 5080 2984 5132 2990
rect 4158 2952 4214 2961
rect 5080 2926 5132 2932
rect 4158 2887 4214 2896
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3804 2650 3832 2790
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 3804 2446 3832 2586
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2318 54 2636 82
rect 3882 82 3938 480
rect 4172 82 4200 2586
rect 5092 2582 5120 2926
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 3882 54 4200 82
rect 5368 82 5396 2858
rect 5460 2650 5488 3878
rect 5644 3194 5672 4014
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 5538 82 5594 480
rect 5368 54 5594 82
rect 7024 82 7052 2586
rect 7392 2553 7420 2586
rect 7378 2544 7434 2553
rect 7378 2479 7434 2488
rect 7944 2446 7972 5850
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7102 82 7158 480
rect 7024 54 7158 82
rect 8496 82 8524 6122
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 9324 4154 9352 7919
rect 10888 6458 10916 9862
rect 11164 9674 11192 12786
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11164 9646 11284 9674
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10888 6254 10916 6394
rect 11256 6254 11284 9646
rect 10876 6248 10928 6254
rect 10782 6216 10838 6225
rect 10876 6190 10928 6196
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 10782 6151 10838 6160
rect 10796 6118 10824 6151
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 11256 5914 11284 6190
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11256 5574 11284 5850
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11440 4690 11468 12038
rect 12452 9081 12480 13806
rect 12438 9072 12494 9081
rect 12438 9007 12494 9016
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12544 4690 12572 5510
rect 12636 4690 12664 13903
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 14752 12850 14780 15302
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 13740 9586 13768 9862
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 17774 9480 17830 9489
rect 17774 9415 17830 9424
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 17788 9110 17816 9415
rect 17880 9178 17908 15943
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 17788 8634 17816 9046
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 17130 6896 17186 6905
rect 16488 6860 16540 6866
rect 17328 6866 17356 7414
rect 17512 7206 17540 7686
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17130 6831 17186 6840
rect 17316 6860 17368 6866
rect 16488 6802 16540 6808
rect 16500 6662 16528 6802
rect 17144 6798 17172 6831
rect 17316 6802 17368 6808
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 16396 6248 16448 6254
rect 16500 6236 16528 6598
rect 16684 6254 16712 6598
rect 16960 6458 16988 6598
rect 17144 6458 17172 6734
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 16448 6208 16528 6236
rect 16396 6190 16448 6196
rect 16304 6112 16356 6118
rect 16356 6072 16436 6100
rect 16304 6054 16356 6060
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 15304 5098 15332 5714
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15304 4758 15332 5034
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 10980 4282 11008 4626
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 9324 4126 9444 4154
rect 9416 4078 9444 4126
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 9416 3738 9444 4014
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 8758 82 8814 480
rect 8496 54 8814 82
rect 10060 82 10088 3946
rect 10980 3942 11008 4218
rect 11440 4078 11468 4626
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10322 82 10378 480
rect 10060 54 10378 82
rect 11624 82 11652 4558
rect 12544 3942 12572 4626
rect 12636 4282 12664 4626
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 11886 82 11942 480
rect 11624 54 11942 82
rect 13280 82 13308 4558
rect 13542 82 13598 480
rect 13280 54 13598 82
rect 754 0 810 54
rect 2318 0 2374 54
rect 3882 0 3938 54
rect 5538 0 5594 54
rect 7102 0 7158 54
rect 8758 0 8814 54
rect 10322 0 10378 54
rect 11886 0 11942 54
rect 13542 0 13598 54
rect 15106 82 15162 480
rect 15396 82 15424 5850
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 5370 15516 5714
rect 16408 5574 16436 6072
rect 16500 5574 16528 6208
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15488 3942 15516 4626
rect 15856 4282 15884 4626
rect 16316 4282 16344 5170
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15488 2854 15516 3878
rect 16408 3398 16436 5510
rect 16776 5370 16804 6394
rect 17236 6322 17264 6734
rect 17328 6390 17356 6802
rect 17512 6662 17540 7142
rect 18156 7002 18184 18634
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 8838 18276 9318
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8362 18276 8774
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18248 7750 18276 8298
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7342 18276 7686
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17316 6384 17368 6390
rect 17316 6326 17368 6332
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5914 16896 6054
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16868 5273 16896 5850
rect 17972 5778 18000 6190
rect 18156 5846 18184 6938
rect 18248 6662 18276 7278
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6186 18276 6598
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17328 5574 17356 5714
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 17328 5030 17356 5510
rect 18340 5370 18368 19110
rect 18432 8634 18460 20198
rect 18984 19922 19012 20198
rect 19260 19990 19288 23582
rect 19522 23520 19578 23582
rect 20456 23582 20774 23610
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 20398 19472 20742
rect 19522 20496 19578 20505
rect 20456 20466 20484 23582
rect 20718 23520 20774 23582
rect 21744 23582 22062 23610
rect 21638 22808 21694 22817
rect 21638 22743 21694 22752
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 19522 20431 19578 20440
rect 20444 20460 20496 20466
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18524 19310 18552 19858
rect 19444 19378 19472 20334
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18524 18873 18552 19246
rect 18510 18864 18566 18873
rect 18510 18799 18566 18808
rect 18524 18766 18552 18799
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18892 10713 18920 15098
rect 18984 12986 19012 18702
rect 19352 18698 19380 19246
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19444 18222 19472 19314
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19536 16794 19564 20431
rect 20444 20402 20496 20408
rect 19614 20360 19670 20369
rect 19614 20295 19670 20304
rect 19628 19378 19656 20295
rect 20640 20262 20668 20946
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 20640 18834 20668 20198
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 19996 18086 20024 18770
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 20074 16824 20130 16833
rect 19524 16788 19576 16794
rect 20074 16759 20130 16768
rect 19524 16730 19576 16736
rect 19536 16046 19564 16730
rect 20088 16114 20116 16759
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19168 13977 19196 15846
rect 19260 15552 19288 15982
rect 19536 15638 19564 15982
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19340 15564 19392 15570
rect 19260 15524 19340 15552
rect 19260 15162 19288 15524
rect 19340 15506 19392 15512
rect 19536 15162 19564 15574
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19154 13968 19210 13977
rect 19536 13938 19564 15098
rect 19154 13903 19210 13912
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 13530 19932 13670
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19536 10810 19564 12718
rect 19628 12442 19656 12718
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 18878 10704 18934 10713
rect 18878 10639 18934 10648
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18524 8498 18552 8910
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18432 5846 18460 7482
rect 18524 7274 18552 8434
rect 18616 8430 18644 8978
rect 18708 8974 18736 9046
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18616 8090 18644 8366
rect 18892 8090 18920 10639
rect 19628 9586 19656 12378
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18984 8498 19012 8910
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18616 6934 18644 8026
rect 18984 7886 19012 8434
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7546 18736 7754
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18984 7478 19012 7822
rect 19076 7818 19104 8366
rect 19444 8294 19472 9386
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7478 19380 7686
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18616 6254 18644 6870
rect 18984 6866 19012 7414
rect 19444 7410 19472 8230
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 18432 5642 18460 5782
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3097 16436 3334
rect 16394 3088 16450 3097
rect 16394 3023 16450 3032
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15106 54 15424 82
rect 16500 82 16528 4558
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 17328 3602 17356 4966
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17880 4282 17908 4762
rect 18340 4690 18368 5306
rect 18524 5166 18552 5714
rect 18708 5574 18736 6054
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18708 5302 18736 5510
rect 18800 5302 18828 5578
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18788 5296 18840 5302
rect 18788 5238 18840 5244
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4826 18552 5102
rect 18708 5098 18736 5238
rect 18696 5092 18748 5098
rect 18696 5034 18748 5040
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18800 4486 18828 5238
rect 18984 5234 19012 6802
rect 19260 6254 19288 6938
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19352 6390 19380 6666
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19352 5574 19380 6326
rect 19444 6322 19472 6734
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19444 5710 19472 6258
rect 19536 5846 19564 9386
rect 19628 7546 19656 9522
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19628 7002 19656 7346
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19628 6662 19656 6938
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18984 4706 19012 5170
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 18984 4678 19104 4706
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 16776 3194 16804 3538
rect 17420 3534 17448 3946
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17236 3194 17264 3334
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17328 3126 17356 3334
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 17420 2650 17448 3470
rect 18432 3466 18460 4422
rect 18800 4282 18828 4422
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18800 3448 18828 4218
rect 18984 4010 19012 4558
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 19076 3534 19104 4678
rect 19168 4185 19196 4966
rect 19352 4486 19380 4966
rect 19444 4826 19472 5646
rect 19616 5160 19668 5166
rect 19616 5102 19668 5108
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19444 4622 19472 4762
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 4214 19380 4422
rect 19340 4208 19392 4214
rect 19154 4176 19210 4185
rect 19340 4150 19392 4156
rect 19154 4111 19210 4120
rect 19064 3528 19116 3534
rect 18984 3488 19064 3516
rect 18880 3460 18932 3466
rect 18800 3420 18880 3448
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17512 2961 17540 3334
rect 18800 3194 18828 3420
rect 18880 3402 18932 3408
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18984 3126 19012 3488
rect 19064 3470 19116 3476
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 17498 2952 17554 2961
rect 17498 2887 17554 2896
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 16762 82 16818 480
rect 16500 54 16818 82
rect 18248 82 18276 2586
rect 19076 2553 19104 3334
rect 19168 2972 19196 4111
rect 19352 3602 19380 4150
rect 19444 3670 19472 4558
rect 19628 4146 19656 5102
rect 19720 4214 19748 10406
rect 20180 7546 20208 13806
rect 20456 13734 20484 13806
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20258 13288 20314 13297
rect 20258 13223 20314 13232
rect 20272 12850 20300 13223
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20364 7478 20392 7686
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20272 7206 20300 7278
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 19708 4208 19760 4214
rect 19708 4150 19760 4156
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19628 3738 19656 4082
rect 19720 3942 19748 4150
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19248 2984 19300 2990
rect 19168 2944 19248 2972
rect 19248 2926 19300 2932
rect 19260 2650 19288 2926
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19062 2544 19118 2553
rect 19062 2479 19118 2488
rect 19352 2292 19380 3538
rect 20088 3058 20116 5782
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 20180 4010 20208 5238
rect 20272 5030 20300 7142
rect 20364 7002 20392 7414
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20364 6322 20392 6938
rect 20456 6848 20484 13670
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20536 6860 20588 6866
rect 20456 6820 20536 6848
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20350 4176 20406 4185
rect 20456 4154 20484 6820
rect 20536 6802 20588 6808
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 6118 20576 6598
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20640 5166 20668 10542
rect 20732 9382 20760 22646
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 20902 20496 20958 20505
rect 20902 20431 20958 20440
rect 20916 20398 20944 20431
rect 21468 20398 21496 20946
rect 21652 20466 21680 22743
rect 21744 22710 21772 23582
rect 22006 23520 22062 23582
rect 23032 23582 23350 23610
rect 21732 22704 21784 22710
rect 21732 22646 21784 22652
rect 23032 21078 23060 23582
rect 23294 23520 23350 23582
rect 23570 22128 23626 22137
rect 23570 22063 23626 22072
rect 23020 21072 23072 21078
rect 23020 21014 23072 21020
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21468 19922 21496 20334
rect 23584 19990 23612 22063
rect 23572 19984 23624 19990
rect 23572 19926 23624 19932
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 21284 19514 21312 19858
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21468 19446 21496 19858
rect 23570 19680 23626 19689
rect 23570 19615 23626 19624
rect 21456 19440 21508 19446
rect 21456 19382 21508 19388
rect 23584 18902 23612 19615
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 21376 18222 21404 18770
rect 21638 18320 21694 18329
rect 21638 18255 21694 18264
rect 21652 18222 21680 18255
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 20824 17542 20852 18158
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20824 12306 20852 17478
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 23570 16144 23626 16153
rect 23570 16079 23626 16088
rect 23584 15638 23612 16079
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 23570 14920 23626 14929
rect 23570 14855 23626 14864
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 23584 13938 23612 14855
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 23570 12608 23626 12617
rect 23570 12543 23626 12552
rect 23584 12374 23612 12543
rect 23572 12368 23624 12374
rect 23572 12310 23624 12316
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 20824 11898 20852 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20824 9518 20852 11834
rect 21284 11558 21312 12242
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 21284 10538 21312 11494
rect 21638 10976 21694 10985
rect 21638 10911 21694 10920
rect 21652 10674 21680 10911
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 23662 10160 23718 10169
rect 23584 10130 23662 10146
rect 21272 10124 21324 10130
rect 21456 10124 21508 10130
rect 21324 10084 21404 10112
rect 21272 10066 21324 10072
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20824 8906 20852 9454
rect 21376 9382 21404 10084
rect 21456 10066 21508 10072
rect 23572 10124 23662 10130
rect 23624 10118 23662 10124
rect 23662 10095 23718 10104
rect 23572 10066 23624 10072
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 7993 20760 8774
rect 20718 7984 20774 7993
rect 20824 7954 20852 8842
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20718 7919 20774 7928
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20732 6662 20760 7278
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21284 6254 21312 6394
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20640 4826 20668 5102
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20406 4126 20484 4154
rect 20350 4111 20406 4120
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19444 2582 19472 2926
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19432 2304 19484 2310
rect 19352 2264 19432 2292
rect 19432 2246 19484 2252
rect 19444 2009 19472 2246
rect 19430 2000 19486 2009
rect 19430 1935 19486 1944
rect 18326 82 18382 480
rect 18248 54 18382 82
rect 15106 0 15162 54
rect 16762 0 16818 54
rect 18326 0 18382 54
rect 19890 82 19946 480
rect 19996 82 20024 2926
rect 20180 1193 20208 3946
rect 20640 3942 20668 4558
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20272 3398 20300 3878
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20640 2961 20668 3878
rect 20732 3670 20760 6190
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 21008 5710 21036 6054
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20824 5234 20852 5510
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 21284 5166 21312 6190
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 4078 20852 4626
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20824 3602 20852 4014
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20626 2952 20682 2961
rect 20626 2887 20682 2896
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 2650 20668 2790
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20824 2446 20852 3538
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20166 1184 20222 1193
rect 20166 1119 20222 1128
rect 19890 54 20024 82
rect 21284 82 21312 2858
rect 21376 2854 21404 9318
rect 21468 8838 21496 10066
rect 23570 8936 23626 8945
rect 23570 8871 23626 8880
rect 21456 8832 21508 8838
rect 21508 8792 21588 8820
rect 21456 8774 21508 8780
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21468 7206 21496 7890
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21468 6866 21496 7142
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21468 5914 21496 6802
rect 21560 5914 21588 8792
rect 23584 8022 23612 8871
rect 23572 8016 23624 8022
rect 23572 7958 23624 7964
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21744 7274 21772 7822
rect 23570 7712 23626 7721
rect 23570 7647 23626 7656
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21638 6352 21694 6361
rect 21638 6287 21694 6296
rect 21652 6254 21680 6287
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21744 6186 21772 7210
rect 23584 6934 23612 7647
rect 23572 6928 23624 6934
rect 23572 6870 23624 6876
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22296 6458 22324 6734
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 5030 21496 5510
rect 21638 5400 21694 5409
rect 22296 5370 22324 5646
rect 21638 5335 21694 5344
rect 22284 5364 22336 5370
rect 21652 5166 21680 5335
rect 22284 5306 22336 5312
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23584 4185 23612 4558
rect 23570 4176 23626 4185
rect 23570 4111 23626 4120
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21468 3194 21496 3538
rect 21560 3505 21588 3946
rect 22836 3528 22888 3534
rect 21546 3496 21602 3505
rect 22836 3470 22888 3476
rect 21546 3431 21602 3440
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21546 82 21602 480
rect 21284 54 21602 82
rect 22848 82 22876 3470
rect 23110 82 23166 480
rect 22848 54 23166 82
rect 19890 0 19946 54
rect 21546 0 21602 54
rect 23110 0 23166 54
<< via2 >>
rect 110 23024 166 23080
rect 110 21256 166 21312
rect 1582 19080 1638 19136
rect 110 17856 166 17912
rect 1398 15816 1454 15872
rect 110 14456 166 14512
rect 1306 12416 1362 12472
rect 110 11056 166 11112
rect 1674 15952 1730 16008
rect 1490 9424 1546 9480
rect 110 9288 166 9344
rect 1674 9016 1730 9072
rect 110 7656 166 7712
rect 110 2488 166 2544
rect 2042 14864 2098 14920
rect 1950 13912 2006 13968
rect 1950 10648 2006 10704
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8114 18808 8170 18864
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 5446 6840 5502 6896
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 15198 20440 15254 20496
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 17866 15952 17922 16008
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 11886 14864 11942 14920
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 12622 13912 12678 13968
rect 9310 7928 9366 7984
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 2226 4664 2282 4720
rect 2502 4020 2504 4040
rect 2504 4020 2556 4040
rect 2556 4020 2558 4040
rect 2502 3984 2558 4020
rect 7838 5208 7894 5264
rect 2594 3032 2650 3088
rect 1490 1400 1546 1456
rect 3422 3984 3478 4040
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 4158 2896 4214 2952
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 7378 2488 7434 2544
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 10782 6160 10838 6216
rect 12438 9016 12494 9072
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 17774 9424 17830 9480
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 17130 6840 17186 6896
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16854 5208 16910 5264
rect 19522 20440 19578 20496
rect 21638 22752 21694 22808
rect 18510 18808 18566 18864
rect 19614 20304 19670 20360
rect 20074 16768 20130 16824
rect 19154 13912 19210 13968
rect 18878 10648 18934 10704
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16394 3032 16450 3088
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 19154 4120 19210 4176
rect 17498 2896 17554 2952
rect 20258 13232 20314 13288
rect 19062 2488 19118 2544
rect 20350 4120 20406 4176
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 20902 20440 20958 20496
rect 23570 22072 23626 22128
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 23570 19624 23626 19680
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 21638 18264 21694 18320
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 23570 16088 23626 16144
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 23570 14864 23626 14920
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 23570 12552 23626 12608
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 21638 10920 21694 10976
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 23662 10104 23718 10160
rect 20718 7928 20774 7984
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 19430 1944 19486 2000
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20626 2896 20682 2952
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 20166 1128 20222 1184
rect 23570 8880 23626 8936
rect 23570 7656 23626 7712
rect 21638 6296 21694 6352
rect 21638 5344 21694 5400
rect 23570 4120 23626 4176
rect 21546 3440 21602 3496
<< metal3 >>
rect 23520 23264 24000 23384
rect 0 23080 480 23112
rect 0 23024 110 23080
rect 166 23024 480 23080
rect 0 22992 480 23024
rect 21633 22810 21699 22813
rect 23614 22810 23674 23264
rect 21633 22808 23674 22810
rect 21633 22752 21638 22808
rect 21694 22752 23674 22808
rect 21633 22750 23674 22752
rect 21633 22747 21699 22750
rect 23520 22130 24000 22160
rect 23484 22128 24000 22130
rect 23484 22072 23570 22128
rect 23626 22072 24000 22128
rect 23484 22070 24000 22072
rect 23520 22040 24000 22070
rect 4944 21792 5264 21793
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 0 21312 480 21344
rect 0 21256 110 21312
rect 166 21256 480 21312
rect 0 21224 480 21256
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 23520 20816 24000 20936
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 15193 20498 15259 20501
rect 19517 20498 19583 20501
rect 20897 20498 20963 20501
rect 15193 20496 20963 20498
rect 15193 20440 15198 20496
rect 15254 20440 19522 20496
rect 19578 20440 20902 20496
rect 20958 20440 20963 20496
rect 15193 20438 20963 20440
rect 15193 20435 15259 20438
rect 19517 20435 19583 20438
rect 20897 20435 20963 20438
rect 19609 20362 19675 20365
rect 23614 20362 23674 20816
rect 19609 20360 23674 20362
rect 19609 20304 19614 20360
rect 19670 20304 23674 20360
rect 19609 20302 23674 20304
rect 19609 20299 19675 20302
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 20095 17264 20096
rect 0 19592 480 19712
rect 23520 19682 24000 19712
rect 23484 19680 24000 19682
rect 23484 19624 23570 19680
rect 23626 19624 24000 19680
rect 23484 19622 24000 19624
rect 4944 19616 5264 19617
rect 62 19138 122 19592
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 23520 19592 24000 19622
rect 20944 19551 21264 19552
rect 1577 19138 1643 19141
rect 62 19136 1643 19138
rect 62 19080 1582 19136
rect 1638 19080 1643 19136
rect 62 19078 1643 19080
rect 1577 19075 1643 19078
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 8109 18866 8175 18869
rect 18505 18866 18571 18869
rect 8109 18864 18571 18866
rect 8109 18808 8114 18864
rect 8170 18808 18510 18864
rect 18566 18808 18571 18864
rect 8109 18806 18571 18808
rect 8109 18803 8175 18806
rect 18505 18803 18571 18806
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 23520 18504 24000 18624
rect 20944 18463 21264 18464
rect 21633 18322 21699 18325
rect 23614 18322 23674 18504
rect 21633 18320 23674 18322
rect 21633 18264 21638 18320
rect 21694 18264 23674 18320
rect 21633 18262 23674 18264
rect 21633 18259 21699 18262
rect 8944 17984 9264 17985
rect 0 17912 480 17944
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 0 17856 110 17912
rect 166 17856 480 17912
rect 0 17824 480 17856
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 23520 17280 24000 17400
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 16831 17264 16832
rect 20069 16826 20135 16829
rect 23614 16826 23674 17280
rect 20069 16824 23674 16826
rect 20069 16768 20074 16824
rect 20130 16768 23674 16824
rect 20069 16766 23674 16768
rect 20069 16763 20135 16766
rect 4944 16352 5264 16353
rect 0 16192 480 16312
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 62 15874 122 16192
rect 23520 16146 24000 16176
rect 23484 16144 24000 16146
rect 23484 16088 23570 16144
rect 23626 16088 24000 16144
rect 23484 16086 24000 16088
rect 23520 16056 24000 16086
rect 1669 16010 1735 16013
rect 17861 16010 17927 16013
rect 1669 16008 17927 16010
rect 1669 15952 1674 16008
rect 1730 15952 17866 16008
rect 17922 15952 17927 16008
rect 1669 15950 17927 15952
rect 1669 15947 1735 15950
rect 17861 15947 17927 15950
rect 1393 15874 1459 15877
rect 62 15872 1459 15874
rect 62 15816 1398 15872
rect 1454 15816 1459 15872
rect 62 15814 1459 15816
rect 1393 15811 1459 15814
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 2037 14922 2103 14925
rect 11881 14922 11947 14925
rect 23520 14922 24000 14952
rect 2037 14920 11947 14922
rect 2037 14864 2042 14920
rect 2098 14864 11886 14920
rect 11942 14864 11947 14920
rect 2037 14862 11947 14864
rect 23484 14920 24000 14922
rect 23484 14864 23570 14920
rect 23626 14864 24000 14920
rect 23484 14862 24000 14864
rect 2037 14859 2103 14862
rect 11881 14859 11947 14862
rect 23520 14832 24000 14862
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 0 14512 480 14544
rect 0 14456 110 14512
rect 166 14456 480 14512
rect 0 14424 480 14456
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 1945 13970 2011 13973
rect 12617 13970 12683 13973
rect 19149 13970 19215 13973
rect 1945 13968 19215 13970
rect 1945 13912 1950 13968
rect 2006 13912 12622 13968
rect 12678 13912 19154 13968
rect 19210 13912 19215 13968
rect 1945 13910 19215 13912
rect 1945 13907 2011 13910
rect 12617 13907 12683 13910
rect 19149 13907 19215 13910
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 23520 13608 24000 13728
rect 16944 13567 17264 13568
rect 20253 13290 20319 13293
rect 23614 13290 23674 13608
rect 20253 13288 23674 13290
rect 20253 13232 20258 13288
rect 20314 13232 23674 13288
rect 20253 13230 23674 13232
rect 20253 13227 20319 13230
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 0 12792 480 12912
rect 62 12474 122 12792
rect 23520 12610 24000 12640
rect 23484 12608 24000 12610
rect 23484 12552 23570 12608
rect 23626 12552 24000 12608
rect 23484 12550 24000 12552
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 23520 12520 24000 12550
rect 16944 12479 17264 12480
rect 1301 12474 1367 12477
rect 62 12472 1367 12474
rect 62 12416 1306 12472
rect 1362 12416 1367 12472
rect 62 12414 1367 12416
rect 1301 12411 1367 12414
rect 4944 12000 5264 12001
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 23520 11296 24000 11416
rect 0 11112 480 11144
rect 0 11056 110 11112
rect 166 11056 480 11112
rect 0 11024 480 11056
rect 21633 10978 21699 10981
rect 23614 10978 23674 11296
rect 21633 10976 23674 10978
rect 21633 10920 21638 10976
rect 21694 10920 23674 10976
rect 21633 10918 23674 10920
rect 21633 10915 21699 10918
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 1945 10706 2011 10709
rect 18873 10706 18939 10709
rect 1945 10704 18939 10706
rect 1945 10648 1950 10704
rect 2006 10648 18878 10704
rect 18934 10648 18939 10704
rect 1945 10646 18939 10648
rect 1945 10643 2011 10646
rect 18873 10643 18939 10646
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 23520 10160 24000 10192
rect 23520 10104 23662 10160
rect 23718 10104 24000 10160
rect 23520 10072 24000 10104
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 1485 9482 1551 9485
rect 17769 9482 17835 9485
rect 1485 9480 17835 9482
rect 1485 9424 1490 9480
rect 1546 9424 17774 9480
rect 17830 9424 17835 9480
rect 1485 9422 17835 9424
rect 1485 9419 1551 9422
rect 17769 9419 17835 9422
rect 0 9344 480 9376
rect 0 9288 110 9344
rect 166 9288 480 9344
rect 0 9256 480 9288
rect 8944 9280 9264 9281
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 9215 17264 9216
rect 1669 9074 1735 9077
rect 12433 9074 12499 9077
rect 1669 9072 12499 9074
rect 1669 9016 1674 9072
rect 1730 9016 12438 9072
rect 12494 9016 12499 9072
rect 1669 9014 12499 9016
rect 1669 9011 1735 9014
rect 12433 9011 12499 9014
rect 23520 8938 24000 8968
rect 23484 8936 24000 8938
rect 23484 8880 23570 8936
rect 23626 8880 24000 8936
rect 23484 8878 24000 8880
rect 23520 8848 24000 8878
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 8127 17264 8128
rect 9305 7986 9371 7989
rect 20713 7986 20779 7989
rect 9305 7984 20779 7986
rect 9305 7928 9310 7984
rect 9366 7928 20718 7984
rect 20774 7928 20779 7984
rect 9305 7926 20779 7928
rect 9305 7923 9371 7926
rect 20713 7923 20779 7926
rect 0 7712 480 7744
rect 23520 7714 24000 7744
rect 0 7656 110 7712
rect 166 7656 480 7712
rect 0 7624 480 7656
rect 23484 7712 24000 7714
rect 23484 7656 23570 7712
rect 23626 7656 24000 7712
rect 23484 7654 24000 7656
rect 4944 7648 5264 7649
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 23520 7624 24000 7654
rect 20944 7583 21264 7584
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 5441 6898 5507 6901
rect 17125 6898 17191 6901
rect 5441 6896 17191 6898
rect 5441 6840 5446 6896
rect 5502 6840 17130 6896
rect 17186 6840 17191 6896
rect 5441 6838 17191 6840
rect 5441 6835 5507 6838
rect 17125 6835 17191 6838
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 23520 6536 24000 6656
rect 20944 6495 21264 6496
rect 21633 6354 21699 6357
rect 23614 6354 23674 6536
rect 21633 6352 23674 6354
rect 21633 6296 21638 6352
rect 21694 6296 23674 6352
rect 21633 6294 23674 6296
rect 21633 6291 21699 6294
rect 10777 6218 10843 6221
rect 62 6216 10843 6218
rect 62 6160 10782 6216
rect 10838 6160 10843 6216
rect 62 6158 10843 6160
rect 62 5976 122 6158
rect 10777 6155 10843 6158
rect 8944 6016 9264 6017
rect 0 5856 480 5976
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 21633 5402 21699 5405
rect 23520 5402 24000 5432
rect 21633 5400 24000 5402
rect 21633 5344 21638 5400
rect 21694 5344 24000 5400
rect 21633 5342 24000 5344
rect 21633 5339 21699 5342
rect 23520 5312 24000 5342
rect 7833 5266 7899 5269
rect 16849 5266 16915 5269
rect 7833 5264 16915 5266
rect 7833 5208 7838 5264
rect 7894 5208 16854 5264
rect 16910 5208 16915 5264
rect 7833 5206 16915 5208
rect 7833 5203 7899 5206
rect 16849 5203 16915 5206
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 2221 4722 2287 4725
rect 62 4720 2287 4722
rect 62 4664 2226 4720
rect 2282 4664 2287 4720
rect 62 4662 2287 4664
rect 62 4344 122 4662
rect 2221 4659 2287 4662
rect 4944 4384 5264 4385
rect 0 4224 480 4344
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 19149 4178 19215 4181
rect 20345 4178 20411 4181
rect 23520 4178 24000 4208
rect 19149 4176 20411 4178
rect 19149 4120 19154 4176
rect 19210 4120 20350 4176
rect 20406 4120 20411 4176
rect 19149 4118 20411 4120
rect 23484 4176 24000 4178
rect 23484 4120 23570 4176
rect 23626 4120 24000 4176
rect 23484 4118 24000 4120
rect 19149 4115 19215 4118
rect 20345 4115 20411 4118
rect 23520 4088 24000 4118
rect 2497 4042 2563 4045
rect 3417 4042 3483 4045
rect 2497 4040 3483 4042
rect 2497 3984 2502 4040
rect 2558 3984 3422 4040
rect 3478 3984 3483 4040
rect 2497 3982 3483 3984
rect 2497 3979 2563 3982
rect 3417 3979 3483 3982
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 21541 3498 21607 3501
rect 21541 3496 23674 3498
rect 21541 3440 21546 3496
rect 21602 3440 23674 3496
rect 21541 3438 23674 3440
rect 21541 3435 21607 3438
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 2589 3090 2655 3093
rect 16389 3090 16455 3093
rect 2589 3088 16455 3090
rect 2589 3032 2594 3088
rect 2650 3032 16394 3088
rect 16450 3032 16455 3088
rect 2589 3030 16455 3032
rect 2589 3027 2655 3030
rect 16389 3027 16455 3030
rect 23614 2984 23674 3438
rect 4153 2954 4219 2957
rect 17493 2954 17559 2957
rect 20621 2954 20687 2957
rect 4153 2952 20687 2954
rect 4153 2896 4158 2952
rect 4214 2896 17498 2952
rect 17554 2896 20626 2952
rect 20682 2896 20687 2952
rect 4153 2894 20687 2896
rect 4153 2891 4219 2894
rect 17493 2891 17559 2894
rect 20621 2891 20687 2894
rect 23520 2864 24000 2984
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 0 2544 480 2576
rect 0 2488 110 2544
rect 166 2488 480 2544
rect 0 2456 480 2488
rect 7373 2546 7439 2549
rect 19057 2546 19123 2549
rect 7373 2544 19123 2546
rect 7373 2488 7378 2544
rect 7434 2488 19062 2544
rect 19118 2488 19123 2544
rect 7373 2486 19123 2488
rect 7373 2483 7439 2486
rect 19057 2483 19123 2486
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 19425 2002 19491 2005
rect 19425 2000 23674 2002
rect 19425 1944 19430 2000
rect 19486 1944 23674 2000
rect 19425 1942 23674 1944
rect 19425 1939 19491 1942
rect 23614 1760 23674 1942
rect 23520 1640 24000 1760
rect 1485 1458 1551 1461
rect 62 1456 1551 1458
rect 62 1400 1490 1456
rect 1546 1400 1551 1456
rect 62 1398 1551 1400
rect 62 944 122 1398
rect 1485 1395 1551 1398
rect 20161 1186 20227 1189
rect 20161 1184 23674 1186
rect 20161 1128 20166 1184
rect 20222 1128 23674 1184
rect 20161 1126 23674 1128
rect 20161 1123 20227 1126
rect 0 824 480 944
rect 23614 672 23674 1126
rect 23520 552 24000 672
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
use scs8hd_or3_4  _035_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1472 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _039_
timestamp 1586364061
transform 1 0 1472 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_17 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_17
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_13
timestamp 1586364061
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__035__B
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_21
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__035__A
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_25 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__035__C
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__B
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _074_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _075_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_45 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_46
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_50
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 774 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_53
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_62 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_92
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__067__D
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_172
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__C
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__C
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_192
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__D
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_203
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 20516 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_210
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_207
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_224
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 130 592
use scs8hd_or3_4  _042_
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__039__B
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__C
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__C
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_20
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_24
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_28
timestamp 1586364061
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_65
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 590 592
use scs8hd_or4_4  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_1  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 130 592
use scs8hd_or4_4  _072_
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__C
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_207
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 130 592
use scs8hd_or3_4  _037_
timestamp 1586364061
transform 1 0 1472 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use scs8hd_inv_8  _032_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__032__A
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__037__C
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_13
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_17
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _027_
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__027__A
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_30
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_nor2_4  _054_
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_8  _030_
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__030__A
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 314 592
use scs8hd_or4_4  _047_
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__047__D
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_inv_8  _033_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__037__A
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__037__B
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_16
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_20
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_28
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _050_
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_115
timestamp 1586364061
transform 1 0 11684 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 15732 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__D
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__D
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__B
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_201
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__033__A
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_28
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_52
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__029__A
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_or4_4  _089_
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_202
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__052__C
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__D
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_207
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_211
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_nor2_4  _068_
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_8  FILLER_6_22
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use scs8hd_nor2_4  _061_
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_74
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_7_81
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_101
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _043_
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__043__B
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_130
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use scs8hd_or4_4  _057_
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _029_
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__D
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_172
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__094__D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__C
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_188
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_or4_4  _084_
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 866 592
use scs8hd_or4_4  _077_
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__D
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_194
timestamp 1586364061
transform 1 0 18952 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_212
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _052_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_228
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__057__D
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _062_
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _094_
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__C
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_195
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_203
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _060_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__034__A
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _040_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_24
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__041__D
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _041_
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_190
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _034_
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__034__B
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__034__D
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_226
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__040__B
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 406 592
use scs8hd_or4_4  _109_
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__D
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_184
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__B
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _059_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__034__C
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_102
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _079_
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_189
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__031__A
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _031_
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_228
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_24
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_nor2_4  _058_
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 314 592
use scs8hd_or4_4  _099_
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__D
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_183
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__D
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_196
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_200
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_208
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_231
timestamp 1586364061
transform 1 0 22356 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _028_
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__028__A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _053_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_207
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_48
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_60
timestamp 1586364061
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _051_
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_211
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_224
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_12
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_24
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__048__B
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__046__B
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_198
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_nor2_4  _049_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _048_
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_108
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _046_
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__038__B
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_209
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_221
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_24
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_48
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_60
timestamp 1586364061
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _038_
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__038__A
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_225
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__036__B
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_133
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_148
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _036_
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__036__A
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_155
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_199
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_203
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_23_227
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_12
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_24
timestamp 1586364061
transform 1 0 3312 0 -1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_30
timestamp 1586364061
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_196
timestamp 1586364061
transform 1 0 19136 0 -1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_219
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_231
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_48
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_200
timestamp 1586364061
transform 1 0 19504 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_231
timestamp 1586364061
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_207
timestamp 1586364061
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_211
timestamp 1586364061
transform 1 0 20516 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 1472 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_13
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_25
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_191
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_195
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_199
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_232
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_35
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_167
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_191
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_31_202
timestamp 1586364061
transform 1 0 19688 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _063_
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_58
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _055_
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_70
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__045__B
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_107
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__044__B
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 15916 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_160
timestamp 1586364061
transform 1 0 15824 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_170
timestamp 1586364061
transform 1 0 16744 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 18492 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_6  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_198
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 1142 592
use scs8hd_nor2_4  _083_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_224
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_232
timestamp 1586364061
transform 1 0 22448 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _065_
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _056_
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_70
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_82
timestamp 1586364061
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _045_
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _044_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_162
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_162
timestamp 1586364061
transform 1 0 16008 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_167
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_174
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 17848 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_188
timestamp 1586364061
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_192
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_191
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 19136 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_205
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_195
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_198
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_211
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_210
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_224
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_228
timestamp 1586364061
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_224
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_232
timestamp 1586364061
transform 1 0 22448 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal2 s 570 23520 626 24000 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 824 480 944 6 address[1]
port 1 nsew default input
rlabel metal2 s 1766 23520 1822 24000 6 address[2]
port 2 nsew default input
rlabel metal3 s 23520 552 24000 672 6 address[3]
port 3 nsew default input
rlabel metal2 s 2318 0 2374 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 23520 1640 24000 1760 6 address[5]
port 5 nsew default input
rlabel metal3 s 23520 2864 24000 2984 6 data_out[0]
port 6 nsew default tristate
rlabel metal3 s 23520 6536 24000 6656 6 data_out[10]
port 7 nsew default tristate
rlabel metal2 s 5538 23520 5594 24000 6 data_out[11]
port 8 nsew default tristate
rlabel metal2 s 8758 0 8814 480 6 data_out[12]
port 9 nsew default tristate
rlabel metal3 s 23520 7624 24000 7744 6 data_out[13]
port 10 nsew default tristate
rlabel metal3 s 23520 8848 24000 8968 6 data_out[14]
port 11 nsew default tristate
rlabel metal2 s 6826 23520 6882 24000 6 data_out[15]
port 12 nsew default tristate
rlabel metal2 s 8114 23520 8170 24000 6 data_out[16]
port 13 nsew default tristate
rlabel metal2 s 9402 23520 9458 24000 6 data_out[17]
port 14 nsew default tristate
rlabel metal2 s 10322 0 10378 480 6 data_out[18]
port 15 nsew default tristate
rlabel metal3 s 23520 10072 24000 10192 6 data_out[19]
port 16 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 data_out[1]
port 17 nsew default tristate
rlabel metal3 s 23520 11296 24000 11416 6 data_out[20]
port 18 nsew default tristate
rlabel metal2 s 11886 0 11942 480 6 data_out[21]
port 19 nsew default tristate
rlabel metal3 s 23520 12520 24000 12640 6 data_out[22]
port 20 nsew default tristate
rlabel metal2 s 10598 23520 10654 24000 6 data_out[23]
port 21 nsew default tristate
rlabel metal3 s 23520 13608 24000 13728 6 data_out[24]
port 22 nsew default tristate
rlabel metal2 s 11886 23520 11942 24000 6 data_out[25]
port 23 nsew default tristate
rlabel metal2 s 13174 23520 13230 24000 6 data_out[26]
port 24 nsew default tristate
rlabel metal3 s 0 5856 480 5976 6 data_out[27]
port 25 nsew default tristate
rlabel metal3 s 0 7624 480 7744 6 data_out[28]
port 26 nsew default tristate
rlabel metal3 s 23520 14832 24000 14952 6 data_out[29]
port 27 nsew default tristate
rlabel metal2 s 5538 0 5594 480 6 data_out[2]
port 28 nsew default tristate
rlabel metal2 s 14462 23520 14518 24000 6 data_out[30]
port 29 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 data_out[31]
port 30 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 data_out[32]
port 31 nsew default tristate
rlabel metal3 s 23520 16056 24000 16176 6 data_out[33]
port 32 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 data_out[34]
port 33 nsew default tristate
rlabel metal2 s 15658 23520 15714 24000 6 data_out[35]
port 34 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 data_out[36]
port 35 nsew default tristate
rlabel metal3 s 23520 17280 24000 17400 6 data_out[37]
port 36 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 data_out[38]
port 37 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 data_out[39]
port 38 nsew default tristate
rlabel metal2 s 7102 0 7158 480 6 data_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 data_out[40]
port 40 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 data_out[41]
port 41 nsew default tristate
rlabel metal3 s 23520 18504 24000 18624 6 data_out[42]
port 42 nsew default tristate
rlabel metal3 s 23520 19592 24000 19712 6 data_out[43]
port 43 nsew default tristate
rlabel metal3 s 23520 20816 24000 20936 6 data_out[44]
port 44 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 data_out[45]
port 45 nsew default tristate
rlabel metal2 s 16946 23520 17002 24000 6 data_out[46]
port 46 nsew default tristate
rlabel metal2 s 18234 23520 18290 24000 6 data_out[47]
port 47 nsew default tristate
rlabel metal2 s 19522 23520 19578 24000 6 data_out[48]
port 48 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 data_out[49]
port 49 nsew default tristate
rlabel metal3 s 23520 4088 24000 4208 6 data_out[4]
port 50 nsew default tristate
rlabel metal2 s 20718 23520 20774 24000 6 data_out[50]
port 51 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 data_out[51]
port 52 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 data_out[52]
port 53 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 data_out[53]
port 54 nsew default tristate
rlabel metal2 s 22006 23520 22062 24000 6 data_out[54]
port 55 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 data_out[55]
port 56 nsew default tristate
rlabel metal3 s 23520 22040 24000 22160 6 data_out[56]
port 57 nsew default tristate
rlabel metal3 s 23520 23264 24000 23384 6 data_out[57]
port 58 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 data_out[58]
port 59 nsew default tristate
rlabel metal2 s 23294 23520 23350 24000 6 data_out[59]
port 60 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 data_out[5]
port 61 nsew default tristate
rlabel metal2 s 23110 0 23166 480 6 data_out[60]
port 62 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 data_out[6]
port 63 nsew default tristate
rlabel metal2 s 3054 23520 3110 24000 6 data_out[7]
port 64 nsew default tristate
rlabel metal3 s 23520 5312 24000 5432 6 data_out[8]
port 65 nsew default tristate
rlabel metal2 s 4342 23520 4398 24000 6 data_out[9]
port 66 nsew default tristate
rlabel metal2 s 754 0 810 480 6 enable
port 67 nsew default input
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 68 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 69 nsew default input
<< end >>
