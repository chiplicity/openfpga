magic
tech sky130A
magscale 1 2
timestamp 1605106472
<< locali >>
rect 5917 16439 5951 16745
rect 12081 6239 12115 6409
rect 3157 3383 3191 3485
<< viali >>
rect 1593 25449 1627 25483
rect 1409 25313 1443 25347
rect 1409 24701 1443 24735
rect 1593 24565 1627 24599
rect 1961 24565 1995 24599
rect 2421 24565 2455 24599
rect 1593 24361 1627 24395
rect 2697 24361 2731 24395
rect 1409 24225 1443 24259
rect 2513 24225 2547 24259
rect 1961 24021 1995 24055
rect 2421 23817 2455 23851
rect 2789 23817 2823 23851
rect 3157 23817 3191 23851
rect 7021 23817 7055 23851
rect 19993 23817 20027 23851
rect 1961 23681 1995 23715
rect 1685 23613 1719 23647
rect 2973 23613 3007 23647
rect 6837 23613 6871 23647
rect 7481 23545 7515 23579
rect 3617 23477 3651 23511
rect 4261 23273 4295 23307
rect 1961 23205 1995 23239
rect 1685 23137 1719 23171
rect 4077 23137 4111 23171
rect 3065 22729 3099 22763
rect 1869 22593 1903 22627
rect 1593 22525 1627 22559
rect 2881 22525 2915 22559
rect 3433 22525 3467 22559
rect 2421 22457 2455 22491
rect 2789 22389 2823 22423
rect 4077 22389 4111 22423
rect 1685 22049 1719 22083
rect 1961 22049 1995 22083
rect 4077 22049 4111 22083
rect 7941 22049 7975 22083
rect 8125 21981 8159 22015
rect 4261 21913 4295 21947
rect 4445 21641 4479 21675
rect 3157 21505 3191 21539
rect 1685 21437 1719 21471
rect 2973 21437 3007 21471
rect 4261 21437 4295 21471
rect 4813 21437 4847 21471
rect 1961 21369 1995 21403
rect 2513 21301 2547 21335
rect 2881 21301 2915 21335
rect 3801 21301 3835 21335
rect 4077 21301 4111 21335
rect 8033 21301 8067 21335
rect 4261 21097 4295 21131
rect 9689 21097 9723 21131
rect 11345 21097 11379 21131
rect 1869 21029 1903 21063
rect 6285 21029 6319 21063
rect 11253 21029 11287 21063
rect 11805 21029 11839 21063
rect 1593 20961 1627 20995
rect 2881 20961 2915 20995
rect 4077 20961 4111 20995
rect 6009 20961 6043 20995
rect 10057 20961 10091 20995
rect 11713 20961 11747 20995
rect 12909 20961 12943 20995
rect 10149 20893 10183 20927
rect 10241 20893 10275 20927
rect 11897 20893 11931 20927
rect 3065 20757 3099 20791
rect 7113 20757 7147 20791
rect 12449 20757 12483 20791
rect 4261 20553 4295 20587
rect 9413 20553 9447 20587
rect 11897 20553 11931 20587
rect 7021 20485 7055 20519
rect 1777 20417 1811 20451
rect 3525 20417 3559 20451
rect 7573 20417 7607 20451
rect 12449 20417 12483 20451
rect 1501 20349 1535 20383
rect 2789 20349 2823 20383
rect 3065 20349 3099 20383
rect 4077 20349 4111 20383
rect 4629 20349 4663 20383
rect 9505 20349 9539 20383
rect 11529 20349 11563 20383
rect 6653 20281 6687 20315
rect 7389 20281 7423 20315
rect 9045 20281 9079 20315
rect 9772 20281 9806 20315
rect 12265 20281 12299 20315
rect 12694 20281 12728 20315
rect 2329 20213 2363 20247
rect 2697 20213 2731 20247
rect 3985 20213 4019 20247
rect 5641 20213 5675 20247
rect 6285 20213 6319 20247
rect 7481 20213 7515 20247
rect 8677 20213 8711 20247
rect 10885 20213 10919 20247
rect 13829 20213 13863 20247
rect 5549 20009 5583 20043
rect 6009 20009 6043 20043
rect 8493 20009 8527 20043
rect 9689 20009 9723 20043
rect 10149 20009 10183 20043
rect 10701 20009 10735 20043
rect 12173 20009 12207 20043
rect 11038 19941 11072 19975
rect 1501 19873 1535 19907
rect 1777 19873 1811 19907
rect 2789 19873 2823 19907
rect 4077 19873 4111 19907
rect 4353 19873 4387 19907
rect 5365 19873 5399 19907
rect 7380 19873 7414 19907
rect 7113 19805 7147 19839
rect 10793 19805 10827 19839
rect 2329 19669 2363 19703
rect 2973 19669 3007 19703
rect 3433 19669 3467 19703
rect 4905 19669 4939 19703
rect 9413 19669 9447 19703
rect 2789 19465 2823 19499
rect 3341 19465 3375 19499
rect 8125 19465 8159 19499
rect 10793 19465 10827 19499
rect 12449 19465 12483 19499
rect 13461 19465 13495 19499
rect 9689 19397 9723 19431
rect 3801 19329 3835 19363
rect 3985 19329 4019 19363
rect 7021 19329 7055 19363
rect 11345 19329 11379 19363
rect 13001 19329 13035 19363
rect 1409 19261 1443 19295
rect 4905 19261 4939 19295
rect 5641 19261 5675 19295
rect 8309 19261 8343 19295
rect 8565 19261 8599 19295
rect 12817 19261 12851 19295
rect 1685 19193 1719 19227
rect 5181 19193 5215 19227
rect 10701 19193 10735 19227
rect 2237 19125 2271 19159
rect 3249 19125 3283 19159
rect 3709 19125 3743 19159
rect 4445 19125 4479 19159
rect 4813 19125 4847 19159
rect 6653 19125 6687 19159
rect 7573 19125 7607 19159
rect 10333 19125 10367 19159
rect 11161 19125 11195 19159
rect 11253 19125 11287 19159
rect 11805 19125 11839 19159
rect 12265 19125 12299 19159
rect 12909 19125 12943 19159
rect 2237 18921 2271 18955
rect 2973 18921 3007 18955
rect 7205 18921 7239 18955
rect 10517 18921 10551 18955
rect 12633 18921 12667 18955
rect 3433 18853 3467 18887
rect 4988 18853 5022 18887
rect 7665 18853 7699 18887
rect 1501 18785 1535 18819
rect 2789 18785 2823 18819
rect 3801 18785 3835 18819
rect 4353 18785 4387 18819
rect 4721 18785 4755 18819
rect 7573 18785 7607 18819
rect 9321 18785 9355 18819
rect 10968 18785 11002 18819
rect 1777 18717 1811 18751
rect 7757 18717 7791 18751
rect 10701 18717 10735 18751
rect 2697 18581 2731 18615
rect 6101 18581 6135 18615
rect 6745 18581 6779 18615
rect 7021 18581 7055 18615
rect 8309 18581 8343 18615
rect 9873 18581 9907 18615
rect 12081 18581 12115 18615
rect 2881 18377 2915 18411
rect 3249 18377 3283 18411
rect 6561 18377 6595 18411
rect 7573 18377 7607 18411
rect 8677 18377 8711 18411
rect 9229 18377 9263 18411
rect 12265 18377 12299 18411
rect 10793 18309 10827 18343
rect 2513 18241 2547 18275
rect 8217 18241 8251 18275
rect 9689 18241 9723 18275
rect 9873 18241 9907 18275
rect 11437 18241 11471 18275
rect 1409 18173 1443 18207
rect 2697 18173 2731 18207
rect 3801 18173 3835 18207
rect 1685 18105 1719 18139
rect 3709 18105 3743 18139
rect 4046 18105 4080 18139
rect 7941 18105 7975 18139
rect 10701 18105 10735 18139
rect 2237 18037 2271 18071
rect 5181 18037 5215 18071
rect 5825 18037 5859 18071
rect 6101 18037 6135 18071
rect 7021 18037 7055 18071
rect 7481 18037 7515 18071
rect 8033 18037 8067 18071
rect 9137 18037 9171 18071
rect 9597 18037 9631 18071
rect 10333 18037 10367 18071
rect 11161 18037 11195 18071
rect 11253 18037 11287 18071
rect 11805 18037 11839 18071
rect 3249 17833 3283 17867
rect 4077 17833 4111 17867
rect 4445 17833 4479 17867
rect 5181 17833 5215 17867
rect 7205 17833 7239 17867
rect 7757 17833 7791 17867
rect 9965 17833 9999 17867
rect 12357 17833 12391 17867
rect 6092 17765 6126 17799
rect 2237 17697 2271 17731
rect 2881 17697 2915 17731
rect 9505 17697 9539 17731
rect 11244 17697 11278 17731
rect 2329 17629 2363 17663
rect 2421 17629 2455 17663
rect 4537 17629 4571 17663
rect 4629 17629 4663 17663
rect 5825 17629 5859 17663
rect 8309 17629 8343 17663
rect 10977 17629 11011 17663
rect 1685 17493 1719 17527
rect 1869 17493 1903 17527
rect 3709 17493 3743 17527
rect 5641 17493 5675 17527
rect 8125 17493 8159 17527
rect 8769 17493 8803 17527
rect 9137 17493 9171 17527
rect 9321 17493 9355 17527
rect 10425 17493 10459 17527
rect 10793 17493 10827 17527
rect 4537 17289 4571 17323
rect 5457 17289 5491 17323
rect 6193 17289 6227 17323
rect 10885 17289 10919 17323
rect 11529 17289 11563 17323
rect 13829 17289 13863 17323
rect 2053 17153 2087 17187
rect 2145 17153 2179 17187
rect 6653 17153 6687 17187
rect 9505 17153 9539 17187
rect 11897 17153 11931 17187
rect 12449 17153 12483 17187
rect 3157 17085 3191 17119
rect 5641 17085 5675 17119
rect 7021 17085 7055 17119
rect 7288 17085 7322 17119
rect 3065 17017 3099 17051
rect 3402 17017 3436 17051
rect 9321 17017 9355 17051
rect 9750 17017 9784 17051
rect 12265 17017 12299 17051
rect 12694 17017 12728 17051
rect 1593 16949 1627 16983
rect 1961 16949 1995 16983
rect 2605 16949 2639 16983
rect 5181 16949 5215 16983
rect 5825 16949 5859 16983
rect 8401 16949 8435 16983
rect 9045 16949 9079 16983
rect 2421 16745 2455 16779
rect 4629 16745 4663 16779
rect 5917 16745 5951 16779
rect 6009 16745 6043 16779
rect 6193 16745 6227 16779
rect 8309 16745 8343 16779
rect 10057 16745 10091 16779
rect 10793 16745 10827 16779
rect 12633 16745 12667 16779
rect 1409 16677 1443 16711
rect 2881 16677 2915 16711
rect 3801 16677 3835 16711
rect 5089 16677 5123 16711
rect 1961 16609 1995 16643
rect 2237 16609 2271 16643
rect 2789 16609 2823 16643
rect 3525 16609 3559 16643
rect 4353 16609 4387 16643
rect 4997 16609 5031 16643
rect 5733 16609 5767 16643
rect 3065 16541 3099 16575
rect 5181 16541 5215 16575
rect 7849 16677 7883 16711
rect 6561 16609 6595 16643
rect 11253 16609 11287 16643
rect 11520 16609 11554 16643
rect 6653 16541 6687 16575
rect 6745 16541 6779 16575
rect 8401 16541 8435 16575
rect 8493 16541 8527 16575
rect 9045 16541 9079 16575
rect 10149 16541 10183 16575
rect 10241 16541 10275 16575
rect 5917 16405 5951 16439
rect 7297 16405 7331 16439
rect 7941 16405 7975 16439
rect 9413 16405 9447 16439
rect 9689 16405 9723 16439
rect 11069 16405 11103 16439
rect 1593 16201 1627 16235
rect 2053 16201 2087 16235
rect 3893 16201 3927 16235
rect 4997 16201 5031 16235
rect 7573 16201 7607 16235
rect 10517 16201 10551 16235
rect 11897 16201 11931 16235
rect 12633 16201 12667 16235
rect 10333 16133 10367 16167
rect 5641 16065 5675 16099
rect 6837 16065 6871 16099
rect 11069 16065 11103 16099
rect 1409 15997 1443 16031
rect 2513 15997 2547 16031
rect 2780 15997 2814 16031
rect 8033 15997 8067 16031
rect 8300 15997 8334 16031
rect 5365 15929 5399 15963
rect 6285 15929 6319 15963
rect 2421 15861 2455 15895
rect 4537 15861 4571 15895
rect 4813 15861 4847 15895
rect 5457 15861 5491 15895
rect 6561 15861 6595 15895
rect 7941 15861 7975 15895
rect 9413 15861 9447 15895
rect 9965 15861 9999 15895
rect 10885 15861 10919 15895
rect 10977 15861 11011 15895
rect 11529 15861 11563 15895
rect 1593 15657 1627 15691
rect 2053 15657 2087 15691
rect 6745 15657 6779 15691
rect 7481 15657 7515 15691
rect 7941 15657 7975 15691
rect 8585 15657 8619 15691
rect 9965 15657 9999 15691
rect 10609 15657 10643 15691
rect 12357 15657 12391 15691
rect 12909 15657 12943 15691
rect 14013 15657 14047 15691
rect 1961 15589 1995 15623
rect 7849 15589 7883 15623
rect 11222 15589 11256 15623
rect 4629 15521 4663 15555
rect 4988 15521 5022 15555
rect 7389 15521 7423 15555
rect 9505 15521 9539 15555
rect 10977 15521 11011 15555
rect 2237 15453 2271 15487
rect 2973 15453 3007 15487
rect 3893 15453 3927 15487
rect 4721 15453 4755 15487
rect 8125 15453 8159 15487
rect 2697 15385 2731 15419
rect 7205 15385 7239 15419
rect 3341 15317 3375 15351
rect 6101 15317 6135 15351
rect 7021 15317 7055 15351
rect 8861 15317 8895 15351
rect 9321 15317 9355 15351
rect 2053 15113 2087 15147
rect 3893 15113 3927 15147
rect 7665 15113 7699 15147
rect 8033 15113 8067 15147
rect 9505 15113 9539 15147
rect 10609 15113 10643 15147
rect 12449 15113 12483 15147
rect 6561 15045 6595 15079
rect 2605 14977 2639 15011
rect 4537 14977 4571 15011
rect 7113 14977 7147 15011
rect 10149 14977 10183 15011
rect 11161 14977 11195 15011
rect 13001 14977 13035 15011
rect 13829 14977 13863 15011
rect 14565 14977 14599 15011
rect 1961 14909 1995 14943
rect 2513 14909 2547 14943
rect 3801 14909 3835 14943
rect 4353 14909 4387 14943
rect 5457 14909 5491 14943
rect 6193 14909 6227 14943
rect 8125 14909 8159 14943
rect 8392 14909 8426 14943
rect 12817 14909 12851 14943
rect 14381 14909 14415 14943
rect 2421 14841 2455 14875
rect 3433 14841 3467 14875
rect 5733 14841 5767 14875
rect 10517 14841 10551 14875
rect 10977 14841 11011 14875
rect 11897 14841 11931 14875
rect 14473 14841 14507 14875
rect 4261 14773 4295 14807
rect 4997 14773 5031 14807
rect 5273 14773 5307 14807
rect 11069 14773 11103 14807
rect 12173 14773 12207 14807
rect 12909 14773 12943 14807
rect 13461 14773 13495 14807
rect 14013 14773 14047 14807
rect 1409 14569 1443 14603
rect 2053 14569 2087 14603
rect 2789 14569 2823 14603
rect 4261 14569 4295 14603
rect 4629 14569 4663 14603
rect 6653 14569 6687 14603
rect 7573 14569 7607 14603
rect 8861 14569 8895 14603
rect 10057 14569 10091 14603
rect 12449 14569 12483 14603
rect 14013 14569 14047 14603
rect 3433 14501 3467 14535
rect 9965 14501 9999 14535
rect 3893 14433 3927 14467
rect 4077 14433 4111 14467
rect 4997 14433 5031 14467
rect 5540 14433 5574 14467
rect 8125 14433 8159 14467
rect 10609 14433 10643 14467
rect 11336 14433 11370 14467
rect 23397 14433 23431 14467
rect 2881 14365 2915 14399
rect 3065 14365 3099 14399
rect 5273 14365 5307 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 11069 14365 11103 14399
rect 7757 14297 7791 14331
rect 2421 14229 2455 14263
rect 9321 14229 9355 14263
rect 23581 14229 23615 14263
rect 1685 14025 1719 14059
rect 10609 14025 10643 14059
rect 23397 14025 23431 14059
rect 2053 13957 2087 13991
rect 3525 13957 3559 13991
rect 4629 13957 4663 13991
rect 7389 13957 7423 13991
rect 11989 13957 12023 13991
rect 12633 13957 12667 13991
rect 23857 13957 23891 13991
rect 4537 13889 4571 13923
rect 5181 13889 5215 13923
rect 8125 13889 8159 13923
rect 10149 13889 10183 13923
rect 11253 13889 11287 13923
rect 2145 13821 2179 13855
rect 6009 13821 6043 13855
rect 6653 13821 6687 13855
rect 7757 13821 7791 13855
rect 8392 13821 8426 13855
rect 10517 13821 10551 13855
rect 11069 13821 11103 13855
rect 23673 13821 23707 13855
rect 24225 13821 24259 13855
rect 2412 13753 2446 13787
rect 4997 13753 5031 13787
rect 10977 13753 11011 13787
rect 4169 13685 4203 13719
rect 5089 13685 5123 13719
rect 5733 13685 5767 13719
rect 6469 13685 6503 13719
rect 6837 13685 6871 13719
rect 9505 13685 9539 13719
rect 11713 13685 11747 13719
rect 2881 13481 2915 13515
rect 6837 13481 6871 13515
rect 7849 13481 7883 13515
rect 10425 13481 10459 13515
rect 12081 13481 12115 13515
rect 1768 13413 1802 13447
rect 3433 13413 3467 13447
rect 5273 13413 5307 13447
rect 8401 13413 8435 13447
rect 1501 13345 1535 13379
rect 4077 13345 4111 13379
rect 4813 13345 4847 13379
rect 5457 13345 5491 13379
rect 5724 13345 5758 13379
rect 8309 13345 8343 13379
rect 10609 13345 10643 13379
rect 10957 13345 10991 13379
rect 22385 13345 22419 13379
rect 4353 13277 4387 13311
rect 8493 13277 8527 13311
rect 10701 13277 10735 13311
rect 8953 13209 8987 13243
rect 10241 13209 10275 13243
rect 3893 13141 3927 13175
rect 7481 13141 7515 13175
rect 7941 13141 7975 13175
rect 9413 13141 9447 13175
rect 9873 13141 9907 13175
rect 22569 13141 22603 13175
rect 1869 12937 1903 12971
rect 5917 12937 5951 12971
rect 6561 12937 6595 12971
rect 7665 12937 7699 12971
rect 8677 12937 8711 12971
rect 9413 12937 9447 12971
rect 12633 12937 12667 12971
rect 3249 12869 3283 12903
rect 7481 12869 7515 12903
rect 10793 12869 10827 12903
rect 2421 12801 2455 12835
rect 3433 12801 3467 12835
rect 7205 12801 7239 12835
rect 8217 12801 8251 12835
rect 10057 12801 10091 12835
rect 12173 12801 12207 12835
rect 3689 12733 3723 12767
rect 6101 12733 6135 12767
rect 8033 12733 8067 12767
rect 11161 12733 11195 12767
rect 22385 12733 22419 12767
rect 2237 12665 2271 12699
rect 2973 12665 3007 12699
rect 5549 12665 5583 12699
rect 9321 12665 9355 12699
rect 9781 12665 9815 12699
rect 11897 12665 11931 12699
rect 1777 12597 1811 12631
rect 2329 12597 2363 12631
rect 4813 12597 4847 12631
rect 8125 12597 8159 12631
rect 9873 12597 9907 12631
rect 10977 12597 11011 12631
rect 11437 12597 11471 12631
rect 13001 12597 13035 12631
rect 13369 12597 13403 12631
rect 1409 12393 1443 12427
rect 2973 12393 3007 12427
rect 3433 12393 3467 12427
rect 5825 12393 5859 12427
rect 7297 12393 7331 12427
rect 8033 12393 8067 12427
rect 8585 12393 8619 12427
rect 11345 12393 11379 12427
rect 6184 12325 6218 12359
rect 1777 12257 1811 12291
rect 1869 12257 1903 12291
rect 4721 12257 4755 12291
rect 4813 12257 4847 12291
rect 5917 12257 5951 12291
rect 9505 12257 9539 12291
rect 9965 12257 9999 12291
rect 10221 12257 10255 12291
rect 12716 12257 12750 12291
rect 21833 12257 21867 12291
rect 2053 12189 2087 12223
rect 3893 12189 3927 12223
rect 4997 12189 5031 12223
rect 9137 12189 9171 12223
rect 12449 12189 12483 12223
rect 4353 12121 4387 12155
rect 2605 12053 2639 12087
rect 5457 12053 5491 12087
rect 8401 12053 8435 12087
rect 11989 12053 12023 12087
rect 12357 12053 12391 12087
rect 13829 12053 13863 12087
rect 22017 12053 22051 12087
rect 1593 11849 1627 11883
rect 2053 11849 2087 11883
rect 2513 11849 2547 11883
rect 5641 11849 5675 11883
rect 6285 11849 6319 11883
rect 10609 11849 10643 11883
rect 12265 11849 12299 11883
rect 13829 11849 13863 11883
rect 14197 11849 14231 11883
rect 12449 11781 12483 11815
rect 3065 11713 3099 11747
rect 4261 11713 4295 11747
rect 8125 11713 8159 11747
rect 11161 11713 11195 11747
rect 12909 11713 12943 11747
rect 13093 11713 13127 11747
rect 1409 11645 1443 11679
rect 8392 11645 8426 11679
rect 10149 11645 10183 11679
rect 10977 11645 11011 11679
rect 21833 11645 21867 11679
rect 2421 11577 2455 11611
rect 2973 11577 3007 11611
rect 3801 11577 3835 11611
rect 4528 11577 4562 11611
rect 7665 11577 7699 11611
rect 8033 11577 8067 11611
rect 2881 11509 2915 11543
rect 4169 11509 4203 11543
rect 6561 11509 6595 11543
rect 7113 11509 7147 11543
rect 9505 11509 9539 11543
rect 10517 11509 10551 11543
rect 11069 11509 11103 11543
rect 11805 11509 11839 11543
rect 12817 11509 12851 11543
rect 13461 11509 13495 11543
rect 2881 11305 2915 11339
rect 3433 11305 3467 11339
rect 4997 11305 5031 11339
rect 6837 11305 6871 11339
rect 7757 11305 7791 11339
rect 8309 11305 8343 11339
rect 8401 11305 8435 11339
rect 9873 11305 9907 11339
rect 10333 11305 10367 11339
rect 12265 11305 12299 11339
rect 12633 11305 12667 11339
rect 13645 11305 13679 11339
rect 3801 11237 3835 11271
rect 4445 11237 4479 11271
rect 5702 11237 5736 11271
rect 7481 11237 7515 11271
rect 1501 11169 1535 11203
rect 1768 11169 1802 11203
rect 4169 11169 4203 11203
rect 5457 11169 5491 11203
rect 10425 11169 10459 11203
rect 8493 11101 8527 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 13277 11101 13311 11135
rect 7941 11033 7975 11067
rect 9413 11033 9447 11067
rect 11713 11033 11747 11067
rect 5273 10965 5307 10999
rect 9045 10965 9079 10999
rect 5457 10761 5491 10795
rect 6285 10761 6319 10795
rect 8861 10761 8895 10795
rect 11069 10761 11103 10795
rect 12265 10761 12299 10795
rect 2513 10625 2547 10659
rect 3249 10625 3283 10659
rect 3709 10625 3743 10659
rect 4721 10625 4755 10659
rect 5733 10625 5767 10659
rect 6929 10625 6963 10659
rect 8585 10625 8619 10659
rect 9505 10625 9539 10659
rect 13001 10625 13035 10659
rect 13461 10625 13495 10659
rect 4629 10557 4663 10591
rect 8493 10557 8527 10591
rect 9689 10557 9723 10591
rect 12817 10557 12851 10591
rect 14197 10557 14231 10591
rect 1593 10489 1627 10523
rect 3985 10489 4019 10523
rect 4537 10489 4571 10523
rect 8401 10489 8435 10523
rect 9321 10489 9355 10523
rect 9934 10489 9968 10523
rect 12909 10489 12943 10523
rect 13829 10489 13863 10523
rect 2053 10421 2087 10455
rect 2605 10421 2639 10455
rect 2973 10421 3007 10455
rect 3065 10421 3099 10455
rect 4169 10421 4203 10455
rect 6653 10421 6687 10455
rect 7573 10421 7607 10455
rect 7849 10421 7883 10455
rect 8033 10421 8067 10455
rect 9229 10421 9263 10455
rect 11437 10421 11471 10455
rect 12449 10421 12483 10455
rect 5089 10217 5123 10251
rect 5641 10217 5675 10251
rect 6009 10217 6043 10251
rect 8217 10217 8251 10251
rect 9413 10217 9447 10251
rect 9689 10217 9723 10251
rect 13369 10217 13403 10251
rect 3341 10149 3375 10183
rect 4537 10149 4571 10183
rect 10057 10149 10091 10183
rect 1676 10081 1710 10115
rect 3893 10081 3927 10115
rect 4445 10081 4479 10115
rect 5549 10081 5583 10115
rect 6101 10081 6135 10115
rect 7573 10081 7607 10115
rect 11693 10081 11727 10115
rect 1409 10013 1443 10047
rect 4629 10013 4663 10047
rect 6285 10013 6319 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 10149 10013 10183 10047
rect 10333 10013 10367 10047
rect 10793 10013 10827 10047
rect 11437 10013 11471 10047
rect 4077 9945 4111 9979
rect 14105 9945 14139 9979
rect 2789 9877 2823 9911
rect 6929 9877 6963 9911
rect 7205 9877 7239 9911
rect 8953 9877 8987 9911
rect 11345 9877 11379 9911
rect 12817 9877 12851 9911
rect 14381 9877 14415 9911
rect 2513 9673 2547 9707
rect 4537 9673 4571 9707
rect 12081 9673 12115 9707
rect 1501 9605 1535 9639
rect 5365 9605 5399 9639
rect 8217 9605 8251 9639
rect 12449 9605 12483 9639
rect 2053 9537 2087 9571
rect 6009 9537 6043 9571
rect 6837 9537 6871 9571
rect 9321 9537 9355 9571
rect 13093 9537 13127 9571
rect 14565 9537 14599 9571
rect 1961 9469 1995 9503
rect 3157 9469 3191 9503
rect 6561 9469 6595 9503
rect 7104 9469 7138 9503
rect 8861 9469 8895 9503
rect 12265 9469 12299 9503
rect 14473 9469 14507 9503
rect 3065 9401 3099 9435
rect 3424 9401 3458 9435
rect 9566 9401 9600 9435
rect 11989 9401 12023 9435
rect 12909 9401 12943 9435
rect 13921 9401 13955 9435
rect 14381 9401 14415 9435
rect 1869 9333 1903 9367
rect 5641 9333 5675 9367
rect 9229 9333 9263 9367
rect 10701 9333 10735 9367
rect 11621 9333 11655 9367
rect 12817 9333 12851 9367
rect 13553 9333 13587 9367
rect 14013 9333 14047 9367
rect 1685 9129 1719 9163
rect 2237 9129 2271 9163
rect 2421 9129 2455 9163
rect 3893 9129 3927 9163
rect 4997 9129 5031 9163
rect 6561 9129 6595 9163
rect 8033 9129 8067 9163
rect 9229 9129 9263 9163
rect 11345 9129 11379 9163
rect 13921 9129 13955 9163
rect 14473 9129 14507 9163
rect 16681 9129 16715 9163
rect 2789 9061 2823 9095
rect 10977 9061 11011 9095
rect 11682 9061 11716 9095
rect 5181 8993 5215 9027
rect 5448 8993 5482 9027
rect 9505 8993 9539 9027
rect 10057 8993 10091 9027
rect 11437 8993 11471 9027
rect 15301 8993 15335 9027
rect 15568 8993 15602 9027
rect 2881 8925 2915 8959
rect 2973 8925 3007 8959
rect 3525 8925 3559 8959
rect 8125 8925 8159 8959
rect 8217 8925 8251 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 7665 8857 7699 8891
rect 9321 8857 9355 8891
rect 12817 8857 12851 8891
rect 4353 8789 4387 8823
rect 4629 8789 4663 8823
rect 7205 8789 7239 8823
rect 8769 8789 8803 8823
rect 9689 8789 9723 8823
rect 13461 8789 13495 8823
rect 13737 8789 13771 8823
rect 3617 8585 3651 8619
rect 6285 8585 6319 8619
rect 8309 8585 8343 8619
rect 9689 8585 9723 8619
rect 10149 8585 10183 8619
rect 11805 8585 11839 8619
rect 4905 8517 4939 8551
rect 6837 8517 6871 8551
rect 8585 8517 8619 8551
rect 12633 8517 12667 8551
rect 15577 8517 15611 8551
rect 16129 8517 16163 8551
rect 2237 8449 2271 8483
rect 4445 8449 4479 8483
rect 5733 8449 5767 8483
rect 7389 8449 7423 8483
rect 9137 8449 9171 8483
rect 10793 8449 10827 8483
rect 11161 8449 11195 8483
rect 13277 8449 13311 8483
rect 5089 8381 5123 8415
rect 7297 8381 7331 8415
rect 9045 8381 9079 8415
rect 10517 8381 10551 8415
rect 13001 8381 13035 8415
rect 14197 8381 14231 8415
rect 20269 8381 20303 8415
rect 21005 8381 21039 8415
rect 2053 8313 2087 8347
rect 2482 8313 2516 8347
rect 4813 8313 4847 8347
rect 5641 8313 5675 8347
rect 6561 8313 6595 8347
rect 7849 8313 7883 8347
rect 8953 8313 8987 8347
rect 12173 8313 12207 8347
rect 13093 8313 13127 8347
rect 14105 8313 14139 8347
rect 14464 8313 14498 8347
rect 16681 8313 16715 8347
rect 20545 8313 20579 8347
rect 1685 8245 1719 8279
rect 5181 8245 5215 8279
rect 5549 8245 5583 8279
rect 7205 8245 7239 8279
rect 10057 8245 10091 8279
rect 10609 8245 10643 8279
rect 13645 8245 13679 8279
rect 2789 8041 2823 8075
rect 3433 8041 3467 8075
rect 4537 8041 4571 8075
rect 8861 8041 8895 8075
rect 9689 8041 9723 8075
rect 10609 8041 10643 8075
rect 13093 8041 13127 8075
rect 14105 8041 14139 8075
rect 14657 8041 14691 8075
rect 15761 8041 15795 8075
rect 18153 8041 18187 8075
rect 3801 7973 3835 8007
rect 6009 7973 6043 8007
rect 9137 7973 9171 8007
rect 10241 7973 10275 8007
rect 11314 7973 11348 8007
rect 1409 7905 1443 7939
rect 1676 7905 1710 7939
rect 5917 7905 5951 7939
rect 7665 7905 7699 7939
rect 8125 7905 8159 7939
rect 10977 7905 11011 7939
rect 14013 7905 14047 7939
rect 15301 7905 15335 7939
rect 16773 7905 16807 7939
rect 17040 7905 17074 7939
rect 6101 7837 6135 7871
rect 8217 7837 8251 7871
rect 8309 7837 8343 7871
rect 11069 7837 11103 7871
rect 14197 7837 14231 7871
rect 5181 7769 5215 7803
rect 7389 7769 7423 7803
rect 4905 7701 4939 7735
rect 5549 7701 5583 7735
rect 6929 7701 6963 7735
rect 7481 7701 7515 7735
rect 7757 7701 7791 7735
rect 10793 7701 10827 7735
rect 12449 7701 12483 7735
rect 13461 7701 13495 7735
rect 13645 7701 13679 7735
rect 16497 7701 16531 7735
rect 4169 7497 4203 7531
rect 4813 7497 4847 7531
rect 9321 7497 9355 7531
rect 12909 7497 12943 7531
rect 13277 7497 13311 7531
rect 15853 7497 15887 7531
rect 6193 7429 6227 7463
rect 8769 7429 8803 7463
rect 1409 7361 1443 7395
rect 5181 7361 5215 7395
rect 6653 7361 6687 7395
rect 9781 7361 9815 7395
rect 16957 7361 16991 7395
rect 2789 7293 2823 7327
rect 3056 7293 3090 7327
rect 7389 7293 7423 7327
rect 7656 7293 7690 7327
rect 9873 7293 9907 7327
rect 10140 7293 10174 7327
rect 13369 7293 13403 7327
rect 13625 7293 13659 7327
rect 19717 7293 19751 7327
rect 20453 7293 20487 7327
rect 2145 7225 2179 7259
rect 2513 7225 2547 7259
rect 16221 7225 16255 7259
rect 16865 7225 16899 7259
rect 19993 7225 20027 7259
rect 5273 7157 5307 7191
rect 5733 7157 5767 7191
rect 7205 7157 7239 7191
rect 11253 7157 11287 7191
rect 11805 7157 11839 7191
rect 12265 7157 12299 7191
rect 14749 7157 14783 7191
rect 16405 7157 16439 7191
rect 16773 7157 16807 7191
rect 17417 7157 17451 7191
rect 1685 6953 1719 6987
rect 3801 6953 3835 6987
rect 6101 6953 6135 6987
rect 8217 6953 8251 6987
rect 11621 6953 11655 6987
rect 13461 6953 13495 6987
rect 14013 6953 14047 6987
rect 5365 6885 5399 6919
rect 10885 6885 10919 6919
rect 12348 6885 12382 6919
rect 2789 6817 2823 6851
rect 2881 6817 2915 6851
rect 6745 6817 6779 6851
rect 7104 6817 7138 6851
rect 8861 6817 8895 6851
rect 9321 6817 9355 6851
rect 9873 6817 9907 6851
rect 11989 6817 12023 6851
rect 12081 6817 12115 6851
rect 14749 6817 14783 6851
rect 15393 6817 15427 6851
rect 16497 6817 16531 6851
rect 17121 6817 17155 6851
rect 20913 6817 20947 6851
rect 2973 6749 3007 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 6837 6749 6871 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 15669 6749 15703 6783
rect 16865 6749 16899 6783
rect 2421 6681 2455 6715
rect 4997 6681 5031 6715
rect 6377 6681 6411 6715
rect 10333 6681 10367 6715
rect 14473 6681 14507 6715
rect 14565 6681 14599 6715
rect 2053 6613 2087 6647
rect 3433 6613 3467 6647
rect 4353 6613 4387 6647
rect 4905 6613 4939 6647
rect 6561 6613 6595 6647
rect 10517 6613 10551 6647
rect 18245 6613 18279 6647
rect 21097 6613 21131 6647
rect 3341 6409 3375 6443
rect 5365 6409 5399 6443
rect 5641 6409 5675 6443
rect 9781 6409 9815 6443
rect 10885 6409 10919 6443
rect 12081 6409 12115 6443
rect 12173 6409 12207 6443
rect 12449 6409 12483 6443
rect 16037 6409 16071 6443
rect 17325 6409 17359 6443
rect 20913 6409 20947 6443
rect 11897 6341 11931 6375
rect 2513 6273 2547 6307
rect 4169 6273 4203 6307
rect 4813 6273 4847 6307
rect 6285 6273 6319 6307
rect 6653 6273 6687 6307
rect 7389 6273 7423 6307
rect 8401 6273 8435 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 14105 6273 14139 6307
rect 18061 6273 18095 6307
rect 2329 6205 2363 6239
rect 4629 6205 4663 6239
rect 7205 6205 7239 6239
rect 12081 6205 12115 6239
rect 12817 6205 12851 6239
rect 13461 6205 13495 6239
rect 14372 6205 14406 6239
rect 16589 6205 16623 6239
rect 19165 6205 19199 6239
rect 19901 6205 19935 6239
rect 3709 6137 3743 6171
rect 7297 6137 7331 6171
rect 7849 6137 7883 6171
rect 8309 6137 8343 6171
rect 8646 6137 8680 6171
rect 11345 6137 11379 6171
rect 14013 6137 14047 6171
rect 16865 6137 16899 6171
rect 19441 6137 19475 6171
rect 1593 6069 1627 6103
rect 1961 6069 1995 6103
rect 2421 6069 2455 6103
rect 3065 6069 3099 6103
rect 4261 6069 4295 6103
rect 4721 6069 4755 6103
rect 6837 6069 6871 6103
rect 10517 6069 10551 6103
rect 15485 6069 15519 6103
rect 16405 6069 16439 6103
rect 17785 6069 17819 6103
rect 18521 6069 18555 6103
rect 1409 5865 1443 5899
rect 1869 5865 1903 5899
rect 3801 5865 3835 5899
rect 4261 5865 4295 5899
rect 6837 5865 6871 5899
rect 7941 5865 7975 5899
rect 9689 5865 9723 5899
rect 10609 5865 10643 5899
rect 12909 5865 12943 5899
rect 13277 5865 13311 5899
rect 13645 5865 13679 5899
rect 14013 5865 14047 5899
rect 14657 5865 14691 5899
rect 16589 5865 16623 5899
rect 17141 5865 17175 5899
rect 17233 5865 17267 5899
rect 18337 5865 18371 5899
rect 2421 5797 2455 5831
rect 8953 5797 8987 5831
rect 9321 5797 9355 5831
rect 11152 5797 11186 5831
rect 18797 5797 18831 5831
rect 1777 5729 1811 5763
rect 4905 5729 4939 5763
rect 5724 5729 5758 5763
rect 8309 5729 8343 5763
rect 15301 5729 15335 5763
rect 18705 5729 18739 5763
rect 2053 5661 2087 5695
rect 5457 5661 5491 5695
rect 8401 5661 8435 5695
rect 8585 5661 8619 5695
rect 10241 5661 10275 5695
rect 10885 5661 10919 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 15485 5661 15519 5695
rect 17325 5661 17359 5695
rect 18889 5661 18923 5695
rect 7849 5593 7883 5627
rect 16773 5593 16807 5627
rect 2881 5525 2915 5559
rect 3157 5525 3191 5559
rect 5273 5525 5307 5559
rect 7481 5525 7515 5559
rect 12265 5525 12299 5559
rect 18061 5525 18095 5559
rect 1685 5321 1719 5355
rect 3249 5321 3283 5355
rect 5181 5321 5215 5355
rect 6653 5321 6687 5355
rect 7389 5321 7423 5355
rect 9413 5321 9447 5355
rect 10885 5321 10919 5355
rect 11437 5321 11471 5355
rect 13645 5321 13679 5355
rect 14105 5321 14139 5355
rect 14933 5321 14967 5355
rect 16957 5321 16991 5355
rect 17417 5321 17451 5355
rect 19441 5321 19475 5355
rect 12449 5253 12483 5287
rect 4721 5185 4755 5219
rect 5733 5185 5767 5219
rect 8585 5185 8619 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 16129 5185 16163 5219
rect 1869 5117 1903 5151
rect 5641 5117 5675 5151
rect 9505 5117 9539 5151
rect 9761 5117 9795 5151
rect 14197 5117 14231 5151
rect 15853 5117 15887 5151
rect 16589 5117 16623 5151
rect 17785 5117 17819 5151
rect 18061 5117 18095 5151
rect 20545 5117 20579 5151
rect 21097 5117 21131 5151
rect 2114 5049 2148 5083
rect 7757 5049 7791 5083
rect 12265 5049 12299 5083
rect 14473 5049 14507 5083
rect 15945 5049 15979 5083
rect 18306 5049 18340 5083
rect 3801 4981 3835 5015
rect 4261 4981 4295 5015
rect 4997 4981 5031 5015
rect 5549 4981 5583 5015
rect 6285 4981 6319 5015
rect 6929 4981 6963 5015
rect 7941 4981 7975 5015
rect 8309 4981 8343 5015
rect 8401 4981 8435 5015
rect 8953 4981 8987 5015
rect 11805 4981 11839 5015
rect 12817 4981 12851 5015
rect 15301 4981 15335 5015
rect 15485 4981 15519 5015
rect 20729 4981 20763 5015
rect 6653 4777 6687 4811
rect 7573 4777 7607 4811
rect 9689 4777 9723 4811
rect 13737 4777 13771 4811
rect 16037 4777 16071 4811
rect 16681 4777 16715 4811
rect 19073 4777 19107 4811
rect 7849 4709 7883 4743
rect 8401 4709 8435 4743
rect 9045 4709 9079 4743
rect 15117 4709 15151 4743
rect 1501 4641 1535 4675
rect 1768 4641 1802 4675
rect 5273 4641 5307 4675
rect 5540 4641 5574 4675
rect 8493 4641 8527 4675
rect 9505 4641 9539 4675
rect 10057 4641 10091 4675
rect 10885 4641 10919 4675
rect 11888 4641 11922 4675
rect 14105 4641 14139 4675
rect 15301 4641 15335 4675
rect 16773 4641 16807 4675
rect 17029 4641 17063 4675
rect 19257 4641 19291 4675
rect 20913 4641 20947 4675
rect 8677 4573 8711 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 11621 4573 11655 4607
rect 15577 4573 15611 4607
rect 13001 4505 13035 4539
rect 14657 4505 14691 4539
rect 2881 4437 2915 4471
rect 3433 4437 3467 4471
rect 3801 4437 3835 4471
rect 4261 4437 4295 4471
rect 4629 4437 4663 4471
rect 5089 4437 5123 4471
rect 8033 4437 8067 4471
rect 14289 4437 14323 4471
rect 18153 4437 18187 4471
rect 18797 4437 18831 4471
rect 19441 4437 19475 4471
rect 19901 4437 19935 4471
rect 21097 4437 21131 4471
rect 3065 4233 3099 4267
rect 8769 4233 8803 4267
rect 9781 4233 9815 4267
rect 10885 4233 10919 4267
rect 14473 4233 14507 4267
rect 5365 4165 5399 4199
rect 9689 4165 9723 4199
rect 2237 4097 2271 4131
rect 2697 4097 2731 4131
rect 10425 4097 10459 4131
rect 12265 4097 12299 4131
rect 15025 4097 15059 4131
rect 15485 4097 15519 4131
rect 17509 4097 17543 4131
rect 18613 4097 18647 4131
rect 19533 4097 19567 4131
rect 20085 4097 20119 4131
rect 20177 4097 20211 4131
rect 2145 4029 2179 4063
rect 3249 4029 3283 4063
rect 3505 4029 3539 4063
rect 6193 4029 6227 4063
rect 6837 4029 6871 4063
rect 10241 4029 10275 4063
rect 12449 4029 12483 4063
rect 12716 4029 12750 4063
rect 18521 4029 18555 4063
rect 19073 4029 19107 4063
rect 19993 4029 20027 4063
rect 21189 4029 21223 4063
rect 21741 4029 21775 4063
rect 7082 3961 7116 3995
rect 9321 3961 9355 3995
rect 15393 3961 15427 3995
rect 15730 3961 15764 3995
rect 17877 3961 17911 3995
rect 18429 3961 18463 3995
rect 22293 3961 22327 3995
rect 1685 3893 1719 3927
rect 2053 3893 2087 3927
rect 4629 3893 4663 3927
rect 5641 3893 5675 3927
rect 6653 3893 6687 3927
rect 8217 3893 8251 3927
rect 10149 3893 10183 3927
rect 11161 3893 11195 3927
rect 11345 3893 11379 3927
rect 11897 3893 11931 3927
rect 13829 3893 13863 3927
rect 16865 3893 16899 3927
rect 18061 3893 18095 3927
rect 19625 3893 19659 3927
rect 21005 3893 21039 3927
rect 21373 3893 21407 3927
rect 2789 3689 2823 3723
rect 7849 3689 7883 3723
rect 8953 3689 8987 3723
rect 9505 3689 9539 3723
rect 12173 3689 12207 3723
rect 16681 3689 16715 3723
rect 17233 3689 17267 3723
rect 18889 3689 18923 3723
rect 1777 3621 1811 3655
rect 2697 3621 2731 3655
rect 8401 3621 8435 3655
rect 9934 3621 9968 3655
rect 17601 3621 17635 3655
rect 20085 3621 20119 3655
rect 2145 3553 2179 3587
rect 5457 3553 5491 3587
rect 5724 3553 5758 3587
rect 7481 3553 7515 3587
rect 8309 3553 8343 3587
rect 9689 3553 9723 3587
rect 12541 3553 12575 3587
rect 13921 3553 13955 3587
rect 14657 3553 14691 3587
rect 15117 3553 15151 3587
rect 15568 3553 15602 3587
rect 18153 3553 18187 3587
rect 19349 3553 19383 3587
rect 20913 3553 20947 3587
rect 22017 3553 22051 3587
rect 24041 3553 24075 3587
rect 2973 3485 3007 3519
rect 3157 3485 3191 3519
rect 4445 3485 4479 3519
rect 8493 3485 8527 3519
rect 12633 3485 12667 3519
rect 12725 3485 12759 3519
rect 14105 3485 14139 3519
rect 15301 3485 15335 3519
rect 18245 3485 18279 3519
rect 18429 3485 18463 3519
rect 19625 3485 19659 3519
rect 2329 3417 2363 3451
rect 3709 3417 3743 3451
rect 7941 3417 7975 3451
rect 11713 3417 11747 3451
rect 12081 3417 12115 3451
rect 13277 3417 13311 3451
rect 13645 3417 13679 3451
rect 17785 3417 17819 3451
rect 3157 3349 3191 3383
rect 3433 3349 3467 3383
rect 4261 3349 4295 3383
rect 5273 3349 5307 3383
rect 6837 3349 6871 3383
rect 11069 3349 11103 3383
rect 21097 3349 21131 3383
rect 22201 3349 22235 3383
rect 24225 3349 24259 3383
rect 3985 3145 4019 3179
rect 6561 3145 6595 3179
rect 8033 3145 8067 3179
rect 10609 3145 10643 3179
rect 11161 3145 11195 3179
rect 11805 3145 11839 3179
rect 12265 3145 12299 3179
rect 12725 3145 12759 3179
rect 14657 3145 14691 3179
rect 15577 3145 15611 3179
rect 17417 3145 17451 3179
rect 17877 3145 17911 3179
rect 19441 3145 19475 3179
rect 20821 3145 20855 3179
rect 21649 3145 21683 3179
rect 22017 3145 22051 3179
rect 23489 3145 23523 3179
rect 24225 3145 24259 3179
rect 5181 3077 5215 3111
rect 6837 3077 6871 3111
rect 10057 3077 10091 3111
rect 11437 3077 11471 3111
rect 15301 3077 15335 3111
rect 18061 3077 18095 3111
rect 23857 3077 23891 3111
rect 1409 3009 1443 3043
rect 5733 3009 5767 3043
rect 7481 3009 7515 3043
rect 8585 3009 8619 3043
rect 13185 3009 13219 3043
rect 16221 3009 16255 3043
rect 16405 3009 16439 3043
rect 16773 3009 16807 3043
rect 18521 3009 18555 3043
rect 18705 3009 18739 3043
rect 19073 3009 19107 3043
rect 21189 3009 21223 3043
rect 2605 2941 2639 2975
rect 5549 2941 5583 2975
rect 5641 2941 5675 2975
rect 7205 2941 7239 2975
rect 8677 2941 8711 2975
rect 8944 2941 8978 2975
rect 11253 2941 11287 2975
rect 13277 2941 13311 2975
rect 13544 2941 13578 2975
rect 16129 2941 16163 2975
rect 18429 2941 18463 2975
rect 19625 2941 19659 2975
rect 20361 2941 20395 2975
rect 20913 2941 20947 2975
rect 22201 2941 22235 2975
rect 22753 2941 22787 2975
rect 23673 2941 23707 2975
rect 2053 2873 2087 2907
rect 2872 2873 2906 2907
rect 5089 2873 5123 2907
rect 6285 2873 6319 2907
rect 19901 2873 19935 2907
rect 2329 2805 2363 2839
rect 4721 2805 4755 2839
rect 7297 2805 7331 2839
rect 15761 2805 15795 2839
rect 22385 2805 22419 2839
rect 1961 2601 1995 2635
rect 2513 2601 2547 2635
rect 3065 2601 3099 2635
rect 5733 2601 5767 2635
rect 9229 2601 9263 2635
rect 9781 2601 9815 2635
rect 10241 2601 10275 2635
rect 11345 2601 11379 2635
rect 12633 2601 12667 2635
rect 13737 2601 13771 2635
rect 15945 2601 15979 2635
rect 16497 2601 16531 2635
rect 18061 2601 18095 2635
rect 19441 2601 19475 2635
rect 24777 2601 24811 2635
rect 2421 2533 2455 2567
rect 3893 2533 3927 2567
rect 4620 2533 4654 2567
rect 10149 2533 10183 2567
rect 16865 2533 16899 2567
rect 19901 2533 19935 2567
rect 21465 2533 21499 2567
rect 4353 2465 4387 2499
rect 6745 2465 6779 2499
rect 7297 2465 7331 2499
rect 8033 2465 8067 2499
rect 11437 2465 11471 2499
rect 13001 2465 13035 2499
rect 14105 2465 14139 2499
rect 14197 2465 14231 2499
rect 15209 2465 15243 2499
rect 15853 2465 15887 2499
rect 17049 2465 17083 2499
rect 17601 2465 17635 2499
rect 18337 2465 18371 2499
rect 19073 2465 19107 2499
rect 19625 2465 19659 2499
rect 20361 2465 20395 2499
rect 21189 2465 21223 2499
rect 21925 2465 21959 2499
rect 22477 2465 22511 2499
rect 23029 2465 23063 2499
rect 2697 2397 2731 2431
rect 3433 2397 3467 2431
rect 6377 2397 6411 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 8677 2397 8711 2431
rect 10425 2397 10459 2431
rect 10793 2397 10827 2431
rect 12081 2397 12115 2431
rect 13093 2397 13127 2431
rect 13277 2397 13311 2431
rect 14933 2397 14967 2431
rect 16037 2397 16071 2431
rect 18521 2397 18555 2431
rect 2053 2329 2087 2363
rect 6929 2329 6963 2363
rect 8309 2329 8343 2363
rect 12449 2329 12483 2363
rect 15485 2329 15519 2363
rect 17233 2329 17267 2363
rect 9505 2261 9539 2295
rect 11621 2261 11655 2295
rect 14381 2261 14415 2295
rect 22661 2261 22695 2295
<< metal1 >>
rect 3234 26324 3240 26376
rect 3292 26364 3298 26376
rect 10042 26364 10048 26376
rect 3292 26336 10048 26364
rect 3292 26324 3298 26336
rect 10042 26324 10048 26336
rect 10100 26324 10106 26376
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1578 25480 1584 25492
rect 1539 25452 1584 25480
rect 1578 25440 1584 25452
rect 1636 25440 1642 25492
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2590 25344 2596 25356
rect 1443 25316 2596 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2590 25304 2596 25316
rect 2648 25304 2654 25356
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1443 24704 1992 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1964 24608 1992 24704
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 1946 24596 1952 24608
rect 1907 24568 1952 24596
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 2409 24599 2467 24605
rect 2409 24565 2421 24599
rect 2455 24596 2467 24599
rect 2590 24596 2596 24608
rect 2455 24568 2596 24596
rect 2455 24565 2467 24568
rect 2409 24559 2467 24565
rect 2590 24556 2596 24568
rect 2648 24556 2654 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 2682 24392 2688 24404
rect 2643 24364 2688 24392
rect 2682 24352 2688 24364
rect 2740 24352 2746 24404
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 2498 24256 2504 24268
rect 2459 24228 2504 24256
rect 2498 24216 2504 24228
rect 2556 24216 2562 24268
rect 1670 24012 1676 24064
rect 1728 24052 1734 24064
rect 1949 24055 2007 24061
rect 1949 24052 1961 24055
rect 1728 24024 1961 24052
rect 1728 24012 1734 24024
rect 1949 24021 1961 24024
rect 1995 24021 2007 24055
rect 1949 24015 2007 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1394 23808 1400 23860
rect 1452 23848 1458 23860
rect 1854 23848 1860 23860
rect 1452 23820 1860 23848
rect 1452 23808 1458 23820
rect 1854 23808 1860 23820
rect 1912 23848 1918 23860
rect 2409 23851 2467 23857
rect 2409 23848 2421 23851
rect 1912 23820 2421 23848
rect 1912 23808 1918 23820
rect 2409 23817 2421 23820
rect 2455 23817 2467 23851
rect 2409 23811 2467 23817
rect 2498 23808 2504 23860
rect 2556 23848 2562 23860
rect 2777 23851 2835 23857
rect 2777 23848 2789 23851
rect 2556 23820 2789 23848
rect 2556 23808 2562 23820
rect 2777 23817 2789 23820
rect 2823 23817 2835 23851
rect 3142 23848 3148 23860
rect 3103 23820 3148 23848
rect 2777 23811 2835 23817
rect 3142 23808 3148 23820
rect 3200 23808 3206 23860
rect 7006 23848 7012 23860
rect 6967 23820 7012 23848
rect 7006 23808 7012 23820
rect 7064 23808 7070 23860
rect 19981 23851 20039 23857
rect 19981 23817 19993 23851
rect 20027 23848 20039 23851
rect 20990 23848 20996 23860
rect 20027 23820 20996 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 20990 23808 20996 23820
rect 21048 23808 21054 23860
rect 1949 23715 2007 23721
rect 1949 23681 1961 23715
rect 1995 23712 2007 23715
rect 2516 23712 2544 23808
rect 1995 23684 2544 23712
rect 1995 23681 2007 23684
rect 1949 23675 2007 23681
rect 1670 23644 1676 23656
rect 1631 23616 1676 23644
rect 1670 23604 1676 23616
rect 1728 23604 1734 23656
rect 2961 23647 3019 23653
rect 2961 23613 2973 23647
rect 3007 23644 3019 23647
rect 6825 23647 6883 23653
rect 3007 23616 3648 23644
rect 3007 23613 3019 23616
rect 2961 23607 3019 23613
rect 3620 23520 3648 23616
rect 6825 23613 6837 23647
rect 6871 23613 6883 23647
rect 6825 23607 6883 23613
rect 6840 23576 6868 23607
rect 7466 23576 7472 23588
rect 6840 23548 7472 23576
rect 7466 23536 7472 23548
rect 7524 23536 7530 23588
rect 3602 23508 3608 23520
rect 3563 23480 3608 23508
rect 3602 23468 3608 23480
rect 3660 23468 3666 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 4249 23307 4307 23313
rect 4249 23304 4261 23307
rect 4212 23276 4261 23304
rect 4212 23264 4218 23276
rect 4249 23273 4261 23276
rect 4295 23273 4307 23307
rect 4249 23267 4307 23273
rect 1946 23236 1952 23248
rect 1907 23208 1952 23236
rect 1946 23196 1952 23208
rect 2004 23196 2010 23248
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23168 1731 23171
rect 2774 23168 2780 23180
rect 1719 23140 2780 23168
rect 1719 23137 1731 23140
rect 1673 23131 1731 23137
rect 2774 23128 2780 23140
rect 2832 23128 2838 23180
rect 3970 23128 3976 23180
rect 4028 23168 4034 23180
rect 4065 23171 4123 23177
rect 4065 23168 4077 23171
rect 4028 23140 4077 23168
rect 4028 23128 4034 23140
rect 4065 23137 4077 23140
rect 4111 23137 4123 23171
rect 4065 23131 4123 23137
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 3050 22760 3056 22772
rect 3011 22732 3056 22760
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 1581 22559 1639 22565
rect 1581 22525 1593 22559
rect 1627 22556 1639 22559
rect 2869 22559 2927 22565
rect 1627 22528 2452 22556
rect 1627 22525 1639 22528
rect 1581 22519 1639 22525
rect 2424 22500 2452 22528
rect 2869 22525 2881 22559
rect 2915 22556 2927 22559
rect 3142 22556 3148 22568
rect 2915 22528 3148 22556
rect 2915 22525 2927 22528
rect 2869 22519 2927 22525
rect 3142 22516 3148 22528
rect 3200 22556 3206 22568
rect 3421 22559 3479 22565
rect 3421 22556 3433 22559
rect 3200 22528 3433 22556
rect 3200 22516 3206 22528
rect 3421 22525 3433 22528
rect 3467 22525 3479 22559
rect 3421 22519 3479 22525
rect 2406 22488 2412 22500
rect 2367 22460 2412 22488
rect 2406 22448 2412 22460
rect 2464 22448 2470 22500
rect 2774 22420 2780 22432
rect 2735 22392 2780 22420
rect 2774 22380 2780 22392
rect 2832 22380 2838 22432
rect 3970 22380 3976 22432
rect 4028 22420 4034 22432
rect 4065 22423 4123 22429
rect 4065 22420 4077 22423
rect 4028 22392 4077 22420
rect 4028 22380 4034 22392
rect 4065 22389 4077 22392
rect 4111 22389 4123 22423
rect 4065 22383 4123 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 3970 22148 3976 22160
rect 2792 22120 3976 22148
rect 1673 22083 1731 22089
rect 1673 22049 1685 22083
rect 1719 22049 1731 22083
rect 1673 22043 1731 22049
rect 1949 22083 2007 22089
rect 1949 22049 1961 22083
rect 1995 22080 2007 22083
rect 2792 22080 2820 22120
rect 3970 22108 3976 22120
rect 4028 22108 4034 22160
rect 4065 22083 4123 22089
rect 4065 22080 4077 22083
rect 1995 22052 2820 22080
rect 3988 22052 4077 22080
rect 1995 22049 2007 22052
rect 1949 22043 2007 22049
rect 1688 22012 1716 22043
rect 3988 22024 4016 22052
rect 4065 22049 4077 22052
rect 4111 22049 4123 22083
rect 4065 22043 4123 22049
rect 7929 22083 7987 22089
rect 7929 22049 7941 22083
rect 7975 22080 7987 22083
rect 8018 22080 8024 22092
rect 7975 22052 8024 22080
rect 7975 22049 7987 22052
rect 7929 22043 7987 22049
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 2958 22012 2964 22024
rect 1688 21984 2964 22012
rect 2958 21972 2964 21984
rect 3016 21972 3022 22024
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 8110 22012 8116 22024
rect 8071 21984 8116 22012
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 4246 21944 4252 21956
rect 4207 21916 4252 21944
rect 4246 21904 4252 21916
rect 4304 21904 4310 21956
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 4430 21672 4436 21684
rect 4391 21644 4436 21672
rect 4430 21632 4436 21644
rect 4488 21632 4494 21684
rect 3142 21536 3148 21548
rect 3103 21508 3148 21536
rect 3142 21496 3148 21508
rect 3200 21496 3206 21548
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21468 1731 21471
rect 2961 21471 3019 21477
rect 1719 21440 2544 21468
rect 1719 21437 1731 21440
rect 1673 21431 1731 21437
rect 1946 21400 1952 21412
rect 1907 21372 1952 21400
rect 1946 21360 1952 21372
rect 2004 21360 2010 21412
rect 2516 21344 2544 21440
rect 2961 21437 2973 21471
rect 3007 21468 3019 21471
rect 4246 21468 4252 21480
rect 3007 21440 3832 21468
rect 4207 21440 4252 21468
rect 3007 21437 3019 21440
rect 2961 21431 3019 21437
rect 3804 21344 3832 21440
rect 4246 21428 4252 21440
rect 4304 21468 4310 21480
rect 4801 21471 4859 21477
rect 4801 21468 4813 21471
rect 4304 21440 4813 21468
rect 4304 21428 4310 21440
rect 4801 21437 4813 21440
rect 4847 21437 4859 21471
rect 4801 21431 4859 21437
rect 2498 21332 2504 21344
rect 2459 21304 2504 21332
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 2869 21335 2927 21341
rect 2869 21301 2881 21335
rect 2915 21332 2927 21335
rect 2958 21332 2964 21344
rect 2915 21304 2964 21332
rect 2915 21301 2927 21304
rect 2869 21295 2927 21301
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 3786 21332 3792 21344
rect 3747 21304 3792 21332
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 3970 21292 3976 21344
rect 4028 21332 4034 21344
rect 4065 21335 4123 21341
rect 4065 21332 4077 21335
rect 4028 21304 4077 21332
rect 4028 21292 4034 21304
rect 4065 21301 4077 21304
rect 4111 21301 4123 21335
rect 8018 21332 8024 21344
rect 7979 21304 8024 21332
rect 4065 21295 4123 21301
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 3510 21088 3516 21140
rect 3568 21128 3574 21140
rect 4249 21131 4307 21137
rect 4249 21128 4261 21131
rect 3568 21100 4261 21128
rect 3568 21088 3574 21100
rect 4249 21097 4261 21100
rect 4295 21097 4307 21131
rect 9674 21128 9680 21140
rect 9635 21100 9680 21128
rect 4249 21091 4307 21097
rect 9674 21088 9680 21100
rect 9732 21088 9738 21140
rect 11330 21128 11336 21140
rect 11291 21100 11336 21128
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 1857 21063 1915 21069
rect 1857 21029 1869 21063
rect 1903 21060 1915 21063
rect 3970 21060 3976 21072
rect 1903 21032 3976 21060
rect 1903 21029 1915 21032
rect 1857 21023 1915 21029
rect 3970 21020 3976 21032
rect 4028 21020 4034 21072
rect 6270 21060 6276 21072
rect 6231 21032 6276 21060
rect 6270 21020 6276 21032
rect 6328 21020 6334 21072
rect 11241 21063 11299 21069
rect 11241 21029 11253 21063
rect 11287 21060 11299 21063
rect 11793 21063 11851 21069
rect 11793 21060 11805 21063
rect 11287 21032 11805 21060
rect 11287 21029 11299 21032
rect 11241 21023 11299 21029
rect 11793 21029 11805 21032
rect 11839 21060 11851 21063
rect 12342 21060 12348 21072
rect 11839 21032 12348 21060
rect 11839 21029 11851 21032
rect 11793 21023 11851 21029
rect 12342 21020 12348 21032
rect 12400 21020 12406 21072
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20992 1639 20995
rect 2314 20992 2320 21004
rect 1627 20964 2320 20992
rect 1627 20961 1639 20964
rect 1581 20955 1639 20961
rect 2314 20952 2320 20964
rect 2372 20952 2378 21004
rect 2866 20992 2872 21004
rect 2827 20964 2872 20992
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 4062 20992 4068 21004
rect 4023 20964 4068 20992
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 5994 20992 6000 21004
rect 5955 20964 6000 20992
rect 5994 20952 6000 20964
rect 6052 20952 6058 21004
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 10045 20995 10103 21001
rect 10045 20992 10057 20995
rect 9732 20964 10057 20992
rect 9732 20952 9738 20964
rect 10045 20961 10057 20964
rect 10091 20961 10103 20995
rect 10045 20955 10103 20961
rect 11701 20995 11759 21001
rect 11701 20961 11713 20995
rect 11747 20992 11759 20995
rect 11974 20992 11980 21004
rect 11747 20964 11980 20992
rect 11747 20961 11759 20964
rect 11701 20955 11759 20961
rect 11974 20952 11980 20964
rect 12032 20992 12038 21004
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12032 20964 12909 20992
rect 12032 20952 12038 20964
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 10134 20924 10140 20936
rect 10095 20896 10140 20924
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 10226 20884 10232 20936
rect 10284 20924 10290 20936
rect 11885 20927 11943 20933
rect 10284 20896 10329 20924
rect 10284 20884 10290 20896
rect 11885 20893 11897 20927
rect 11931 20893 11943 20927
rect 11885 20887 11943 20893
rect 11514 20816 11520 20868
rect 11572 20856 11578 20868
rect 11900 20856 11928 20887
rect 11572 20828 11928 20856
rect 11572 20816 11578 20828
rect 3050 20788 3056 20800
rect 3011 20760 3056 20788
rect 3050 20748 3056 20760
rect 3108 20748 3114 20800
rect 7101 20791 7159 20797
rect 7101 20757 7113 20791
rect 7147 20788 7159 20791
rect 7558 20788 7564 20800
rect 7147 20760 7564 20788
rect 7147 20757 7159 20760
rect 7101 20751 7159 20757
rect 7558 20748 7564 20760
rect 7616 20748 7622 20800
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 12492 20760 12537 20788
rect 12492 20748 12498 20760
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 4246 20584 4252 20596
rect 4207 20556 4252 20584
rect 4246 20544 4252 20556
rect 4304 20544 4310 20596
rect 9401 20587 9459 20593
rect 9401 20553 9413 20587
rect 9447 20584 9459 20587
rect 9674 20584 9680 20596
rect 9447 20556 9680 20584
rect 9447 20553 9459 20556
rect 9401 20547 9459 20553
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 11885 20587 11943 20593
rect 11885 20553 11897 20587
rect 11931 20584 11943 20587
rect 11974 20584 11980 20596
rect 11931 20556 11980 20584
rect 11931 20553 11943 20556
rect 11885 20547 11943 20553
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 5994 20476 6000 20528
rect 6052 20516 6058 20528
rect 7009 20519 7067 20525
rect 7009 20516 7021 20519
rect 6052 20488 7021 20516
rect 6052 20476 6058 20488
rect 7009 20485 7021 20488
rect 7055 20485 7067 20519
rect 7009 20479 7067 20485
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 2866 20448 2872 20460
rect 1811 20420 2872 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 2866 20408 2872 20420
rect 2924 20448 2930 20460
rect 3513 20451 3571 20457
rect 3513 20448 3525 20451
rect 2924 20420 3525 20448
rect 2924 20408 2930 20420
rect 3513 20417 3525 20420
rect 3559 20417 3571 20451
rect 7558 20448 7564 20460
rect 7519 20420 7564 20448
rect 3513 20411 3571 20417
rect 7558 20408 7564 20420
rect 7616 20408 7622 20460
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 12492 20420 12537 20448
rect 12492 20408 12498 20420
rect 1489 20383 1547 20389
rect 1489 20349 1501 20383
rect 1535 20380 1547 20383
rect 2777 20383 2835 20389
rect 1535 20352 2360 20380
rect 1535 20349 1547 20352
rect 1489 20343 1547 20349
rect 2332 20253 2360 20352
rect 2777 20349 2789 20383
rect 2823 20349 2835 20383
rect 2777 20343 2835 20349
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20380 3111 20383
rect 4065 20383 4123 20389
rect 4065 20380 4077 20383
rect 3099 20352 4077 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 4065 20349 4077 20352
rect 4111 20380 4123 20383
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 4111 20352 4629 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 9490 20380 9496 20392
rect 9451 20352 9496 20380
rect 4617 20343 4675 20349
rect 2317 20247 2375 20253
rect 2317 20213 2329 20247
rect 2363 20244 2375 20247
rect 2406 20244 2412 20256
rect 2363 20216 2412 20244
rect 2363 20213 2375 20216
rect 2317 20207 2375 20213
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 2685 20247 2743 20253
rect 2685 20213 2697 20247
rect 2731 20244 2743 20247
rect 2792 20244 2820 20343
rect 9490 20340 9496 20352
rect 9548 20340 9554 20392
rect 10226 20380 10232 20392
rect 9692 20352 10232 20380
rect 6641 20315 6699 20321
rect 6641 20281 6653 20315
rect 6687 20312 6699 20315
rect 6914 20312 6920 20324
rect 6687 20284 6920 20312
rect 6687 20281 6699 20284
rect 6641 20275 6699 20281
rect 6914 20272 6920 20284
rect 6972 20312 6978 20324
rect 7377 20315 7435 20321
rect 7377 20312 7389 20315
rect 6972 20284 7389 20312
rect 6972 20272 6978 20284
rect 7377 20281 7389 20284
rect 7423 20281 7435 20315
rect 7377 20275 7435 20281
rect 9033 20315 9091 20321
rect 9033 20281 9045 20315
rect 9079 20312 9091 20315
rect 9692 20312 9720 20352
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 11514 20380 11520 20392
rect 11475 20352 11520 20380
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 9766 20321 9772 20324
rect 9079 20284 9720 20312
rect 9079 20281 9091 20284
rect 9033 20275 9091 20281
rect 9760 20275 9772 20321
rect 9824 20312 9830 20324
rect 9824 20284 9908 20312
rect 9766 20272 9772 20275
rect 9824 20272 9830 20284
rect 3326 20244 3332 20256
rect 2731 20216 3332 20244
rect 2731 20213 2743 20216
rect 2685 20207 2743 20213
rect 3326 20204 3332 20216
rect 3384 20204 3390 20256
rect 3973 20247 4031 20253
rect 3973 20213 3985 20247
rect 4019 20244 4031 20247
rect 4062 20244 4068 20256
rect 4019 20216 4068 20244
rect 4019 20213 4031 20216
rect 3973 20207 4031 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5629 20247 5687 20253
rect 5629 20213 5641 20247
rect 5675 20244 5687 20247
rect 6178 20244 6184 20256
rect 5675 20216 6184 20244
rect 5675 20213 5687 20216
rect 5629 20207 5687 20213
rect 6178 20204 6184 20216
rect 6236 20204 6242 20256
rect 6273 20247 6331 20253
rect 6273 20213 6285 20247
rect 6319 20244 6331 20247
rect 7466 20244 7472 20256
rect 6319 20216 7472 20244
rect 6319 20213 6331 20216
rect 6273 20207 6331 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 8665 20247 8723 20253
rect 8665 20213 8677 20247
rect 8711 20244 8723 20247
rect 9775 20244 9803 20272
rect 8711 20216 9803 20244
rect 10244 20244 10272 20340
rect 12158 20272 12164 20324
rect 12216 20312 12222 20324
rect 12253 20315 12311 20321
rect 12253 20312 12265 20315
rect 12216 20284 12265 20312
rect 12216 20272 12222 20284
rect 12253 20281 12265 20284
rect 12299 20312 12311 20315
rect 12682 20315 12740 20321
rect 12682 20312 12694 20315
rect 12299 20284 12694 20312
rect 12299 20281 12311 20284
rect 12253 20275 12311 20281
rect 12682 20281 12694 20284
rect 12728 20281 12740 20315
rect 12682 20275 12740 20281
rect 10686 20244 10692 20256
rect 10244 20216 10692 20244
rect 8711 20213 8723 20216
rect 8665 20207 8723 20213
rect 10686 20204 10692 20216
rect 10744 20244 10750 20256
rect 10873 20247 10931 20253
rect 10873 20244 10885 20247
rect 10744 20216 10885 20244
rect 10744 20204 10750 20216
rect 10873 20213 10885 20216
rect 10919 20213 10931 20247
rect 13814 20244 13820 20256
rect 13775 20216 13820 20244
rect 10873 20207 10931 20213
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 5534 20040 5540 20052
rect 5495 20012 5540 20040
rect 5534 20000 5540 20012
rect 5592 20000 5598 20052
rect 5994 20040 6000 20052
rect 5955 20012 6000 20040
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 7558 20000 7564 20052
rect 7616 20040 7622 20052
rect 8110 20040 8116 20052
rect 7616 20012 8116 20040
rect 7616 20000 7622 20012
rect 8110 20000 8116 20012
rect 8168 20040 8174 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 8168 20012 8493 20040
rect 8168 20000 8174 20012
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 9674 20040 9680 20052
rect 9635 20012 9680 20040
rect 8481 20003 8539 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10134 20040 10140 20052
rect 10095 20012 10140 20040
rect 10134 20000 10140 20012
rect 10192 20000 10198 20052
rect 10686 20040 10692 20052
rect 10647 20012 10692 20040
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 12158 20040 12164 20052
rect 12119 20012 12164 20040
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 10704 19972 10732 20000
rect 11026 19975 11084 19981
rect 11026 19972 11038 19975
rect 10704 19944 11038 19972
rect 11026 19941 11038 19944
rect 11072 19941 11084 19975
rect 11026 19935 11084 19941
rect 1486 19904 1492 19916
rect 1447 19876 1492 19904
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 2774 19904 2780 19916
rect 1811 19876 2780 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2774 19864 2780 19876
rect 2832 19904 2838 19916
rect 4062 19904 4068 19916
rect 2832 19876 2877 19904
rect 4023 19876 4068 19904
rect 2832 19864 2838 19876
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4341 19907 4399 19913
rect 4341 19873 4353 19907
rect 4387 19904 4399 19907
rect 5353 19907 5411 19913
rect 5353 19904 5365 19907
rect 4387 19876 5365 19904
rect 4387 19873 4399 19876
rect 4341 19867 4399 19873
rect 5353 19873 5365 19876
rect 5399 19904 5411 19907
rect 5442 19904 5448 19916
rect 5399 19876 5448 19904
rect 5399 19873 5411 19876
rect 5353 19867 5411 19873
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 7374 19913 7380 19916
rect 7368 19904 7380 19913
rect 7335 19876 7380 19904
rect 7368 19867 7380 19876
rect 7374 19864 7380 19867
rect 7432 19864 7438 19916
rect 7098 19836 7104 19848
rect 7059 19808 7104 19836
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 10686 19796 10692 19848
rect 10744 19836 10750 19848
rect 10781 19839 10839 19845
rect 10781 19836 10793 19839
rect 10744 19808 10793 19836
rect 10744 19796 10750 19808
rect 10781 19805 10793 19808
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 2314 19700 2320 19712
rect 2275 19672 2320 19700
rect 2314 19660 2320 19672
rect 2372 19660 2378 19712
rect 2958 19700 2964 19712
rect 2919 19672 2964 19700
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 3418 19700 3424 19712
rect 3379 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 4890 19700 4896 19712
rect 4851 19672 4896 19700
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 9401 19703 9459 19709
rect 9401 19700 9413 19703
rect 8352 19672 9413 19700
rect 8352 19660 8358 19672
rect 9401 19669 9413 19672
rect 9447 19700 9459 19703
rect 9490 19700 9496 19712
rect 9447 19672 9496 19700
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3326 19496 3332 19508
rect 2832 19468 2877 19496
rect 3287 19468 3332 19496
rect 2832 19456 2838 19468
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 8110 19496 8116 19508
rect 8071 19468 8116 19496
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10781 19499 10839 19505
rect 10781 19496 10793 19499
rect 10192 19468 10793 19496
rect 10192 19456 10198 19468
rect 10781 19465 10793 19468
rect 10827 19465 10839 19499
rect 10781 19459 10839 19465
rect 12342 19456 12348 19508
rect 12400 19496 12406 19508
rect 12437 19499 12495 19505
rect 12437 19496 12449 19499
rect 12400 19468 12449 19496
rect 12400 19456 12406 19468
rect 12437 19465 12449 19468
rect 12483 19465 12495 19499
rect 12437 19459 12495 19465
rect 12526 19456 12532 19508
rect 12584 19496 12590 19508
rect 13449 19499 13507 19505
rect 13449 19496 13461 19499
rect 12584 19468 13461 19496
rect 12584 19456 12590 19468
rect 13449 19465 13461 19468
rect 13495 19465 13507 19499
rect 13449 19459 13507 19465
rect 3418 19320 3424 19372
rect 3476 19360 3482 19372
rect 3786 19360 3792 19372
rect 3476 19332 3792 19360
rect 3476 19320 3482 19332
rect 3786 19320 3792 19332
rect 3844 19320 3850 19372
rect 3970 19360 3976 19372
rect 3931 19332 3976 19360
rect 3970 19320 3976 19332
rect 4028 19320 4034 19372
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6972 19332 7021 19360
rect 6972 19320 6978 19332
rect 7009 19329 7021 19332
rect 7055 19329 7067 19363
rect 8128 19360 8156 19456
rect 9677 19431 9735 19437
rect 9677 19397 9689 19431
rect 9723 19397 9735 19431
rect 9677 19391 9735 19397
rect 9692 19360 9720 19391
rect 9766 19360 9772 19372
rect 8128 19332 8432 19360
rect 9679 19332 9772 19360
rect 7009 19323 7067 19329
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19261 1455 19295
rect 1397 19255 1455 19261
rect 1412 19156 1440 19255
rect 4798 19252 4804 19304
rect 4856 19292 4862 19304
rect 4893 19295 4951 19301
rect 4893 19292 4905 19295
rect 4856 19264 4905 19292
rect 4856 19252 4862 19264
rect 4893 19261 4905 19264
rect 4939 19261 4951 19295
rect 4893 19255 4951 19261
rect 5534 19252 5540 19304
rect 5592 19292 5598 19304
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5592 19264 5641 19292
rect 5592 19252 5598 19264
rect 5629 19261 5641 19264
rect 5675 19261 5687 19295
rect 8294 19292 8300 19304
rect 8255 19264 8300 19292
rect 5629 19255 5687 19261
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8404 19292 8432 19332
rect 9766 19320 9772 19332
rect 9824 19360 9830 19372
rect 11333 19363 11391 19369
rect 11333 19360 11345 19363
rect 9824 19332 11345 19360
rect 9824 19320 9830 19332
rect 11333 19329 11345 19332
rect 11379 19329 11391 19363
rect 11333 19323 11391 19329
rect 12158 19320 12164 19372
rect 12216 19360 12222 19372
rect 12618 19360 12624 19372
rect 12216 19332 12624 19360
rect 12216 19320 12222 19332
rect 12618 19320 12624 19332
rect 12676 19360 12682 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12676 19332 13001 19360
rect 12676 19320 12682 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 8553 19295 8611 19301
rect 8553 19292 8565 19295
rect 8404 19264 8565 19292
rect 8553 19261 8565 19264
rect 8599 19261 8611 19295
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 8553 19255 8611 19261
rect 11808 19264 12817 19292
rect 1673 19227 1731 19233
rect 1673 19193 1685 19227
rect 1719 19224 1731 19227
rect 2774 19224 2780 19236
rect 1719 19196 2780 19224
rect 1719 19193 1731 19196
rect 1673 19187 1731 19193
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 4154 19184 4160 19236
rect 4212 19224 4218 19236
rect 5169 19227 5227 19233
rect 5169 19224 5181 19227
rect 4212 19196 5181 19224
rect 4212 19184 4218 19196
rect 5169 19193 5181 19196
rect 5215 19193 5227 19227
rect 5169 19187 5227 19193
rect 10689 19227 10747 19233
rect 10689 19193 10701 19227
rect 10735 19224 10747 19227
rect 10735 19196 11284 19224
rect 10735 19193 10747 19196
rect 10689 19187 10747 19193
rect 2225 19159 2283 19165
rect 2225 19156 2237 19159
rect 1412 19128 2237 19156
rect 2225 19125 2237 19128
rect 2271 19156 2283 19159
rect 2498 19156 2504 19168
rect 2271 19128 2504 19156
rect 2271 19125 2283 19128
rect 2225 19119 2283 19125
rect 2498 19116 2504 19128
rect 2556 19116 2562 19168
rect 2590 19116 2596 19168
rect 2648 19156 2654 19168
rect 3237 19159 3295 19165
rect 3237 19156 3249 19159
rect 2648 19128 3249 19156
rect 2648 19116 2654 19128
rect 3237 19125 3249 19128
rect 3283 19156 3295 19159
rect 3697 19159 3755 19165
rect 3697 19156 3709 19159
rect 3283 19128 3709 19156
rect 3283 19125 3295 19128
rect 3237 19119 3295 19125
rect 3697 19125 3709 19128
rect 3743 19125 3755 19159
rect 3697 19119 3755 19125
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4430 19156 4436 19168
rect 4120 19128 4436 19156
rect 4120 19116 4126 19128
rect 4430 19116 4436 19128
rect 4488 19116 4494 19168
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 4890 19116 4896 19168
rect 4948 19156 4954 19168
rect 6641 19159 6699 19165
rect 6641 19156 6653 19159
rect 4948 19128 6653 19156
rect 4948 19116 4954 19128
rect 6641 19125 6653 19128
rect 6687 19156 6699 19159
rect 6730 19156 6736 19168
rect 6687 19128 6736 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6730 19116 6736 19128
rect 6788 19156 6794 19168
rect 7098 19156 7104 19168
rect 6788 19128 7104 19156
rect 6788 19116 6794 19128
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7374 19116 7380 19168
rect 7432 19156 7438 19168
rect 7561 19159 7619 19165
rect 7561 19156 7573 19159
rect 7432 19128 7573 19156
rect 7432 19116 7438 19128
rect 7561 19125 7573 19128
rect 7607 19156 7619 19159
rect 8662 19156 8668 19168
rect 7607 19128 8668 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 9122 19116 9128 19168
rect 9180 19156 9186 19168
rect 11256 19165 11284 19196
rect 11808 19168 11836 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 10321 19159 10379 19165
rect 10321 19156 10333 19159
rect 9180 19128 10333 19156
rect 9180 19116 9186 19128
rect 10321 19125 10333 19128
rect 10367 19156 10379 19159
rect 11149 19159 11207 19165
rect 11149 19156 11161 19159
rect 10367 19128 11161 19156
rect 10367 19125 10379 19128
rect 10321 19119 10379 19125
rect 11149 19125 11161 19128
rect 11195 19125 11207 19159
rect 11149 19119 11207 19125
rect 11241 19159 11299 19165
rect 11241 19125 11253 19159
rect 11287 19156 11299 19159
rect 11330 19156 11336 19168
rect 11287 19128 11336 19156
rect 11287 19125 11299 19128
rect 11241 19119 11299 19125
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 11790 19156 11796 19168
rect 11751 19128 11796 19156
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 12897 19159 12955 19165
rect 12897 19156 12909 19159
rect 12299 19128 12909 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 12897 19125 12909 19128
rect 12943 19156 12955 19159
rect 14366 19156 14372 19168
rect 12943 19128 14372 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 2222 18952 2228 18964
rect 1544 18924 2228 18952
rect 1544 18912 1550 18924
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 2958 18952 2964 18964
rect 2919 18924 2964 18952
rect 2958 18912 2964 18924
rect 3016 18912 3022 18964
rect 7190 18952 7196 18964
rect 7151 18924 7196 18952
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 10505 18955 10563 18961
rect 10505 18952 10517 18955
rect 9824 18924 10517 18952
rect 9824 18912 9830 18924
rect 10505 18921 10517 18924
rect 10551 18921 10563 18955
rect 12618 18952 12624 18964
rect 12579 18924 12624 18952
rect 10505 18915 10563 18921
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 3421 18887 3479 18893
rect 3421 18853 3433 18887
rect 3467 18884 3479 18887
rect 3970 18884 3976 18896
rect 3467 18856 3976 18884
rect 3467 18853 3479 18856
rect 3421 18847 3479 18853
rect 3970 18844 3976 18856
rect 4028 18884 4034 18896
rect 4976 18887 5034 18893
rect 4976 18884 4988 18887
rect 4028 18856 4988 18884
rect 4028 18844 4034 18856
rect 4976 18853 4988 18856
rect 5022 18884 5034 18887
rect 5166 18884 5172 18896
rect 5022 18856 5172 18884
rect 5022 18853 5034 18856
rect 4976 18847 5034 18853
rect 5166 18844 5172 18856
rect 5224 18844 5230 18896
rect 6914 18844 6920 18896
rect 6972 18884 6978 18896
rect 7653 18887 7711 18893
rect 7653 18884 7665 18887
rect 6972 18856 7665 18884
rect 6972 18844 6978 18856
rect 7653 18853 7665 18856
rect 7699 18853 7711 18887
rect 7653 18847 7711 18853
rect 1489 18819 1547 18825
rect 1489 18785 1501 18819
rect 1535 18785 1547 18819
rect 1489 18779 1547 18785
rect 1504 18680 1532 18779
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 3234 18816 3240 18828
rect 2832 18788 3240 18816
rect 2832 18776 2838 18788
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 3789 18819 3847 18825
rect 3789 18785 3801 18819
rect 3835 18816 3847 18819
rect 3878 18816 3884 18828
rect 3835 18788 3884 18816
rect 3835 18785 3847 18788
rect 3789 18779 3847 18785
rect 3878 18776 3884 18788
rect 3936 18816 3942 18828
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 3936 18788 4353 18816
rect 3936 18776 3942 18788
rect 4341 18785 4353 18788
rect 4387 18816 4399 18819
rect 4706 18816 4712 18828
rect 4387 18788 4712 18816
rect 4387 18785 4399 18788
rect 4341 18779 4399 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 6178 18776 6184 18828
rect 6236 18816 6242 18828
rect 10962 18825 10968 18828
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 6236 18788 7573 18816
rect 6236 18776 6242 18788
rect 7561 18785 7573 18788
rect 7607 18785 7619 18819
rect 7561 18779 7619 18785
rect 9309 18819 9367 18825
rect 9309 18785 9321 18819
rect 9355 18816 9367 18819
rect 10956 18816 10968 18825
rect 9355 18788 10968 18816
rect 9355 18785 9367 18788
rect 9309 18779 9367 18785
rect 10956 18779 10968 18788
rect 10962 18776 10968 18779
rect 11020 18776 11026 18828
rect 1762 18748 1768 18760
rect 1723 18720 1768 18748
rect 1762 18708 1768 18720
rect 1820 18708 1826 18760
rect 7742 18748 7748 18760
rect 7703 18720 7748 18748
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 10686 18748 10692 18760
rect 10647 18720 10692 18748
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 1504 18652 2728 18680
rect 2700 18624 2728 18652
rect 2682 18612 2688 18624
rect 2643 18584 2688 18612
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 6086 18612 6092 18624
rect 6047 18584 6092 18612
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 6730 18612 6736 18624
rect 6691 18584 6736 18612
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 6914 18572 6920 18624
rect 6972 18612 6978 18624
rect 7009 18615 7067 18621
rect 7009 18612 7021 18615
rect 6972 18584 7021 18612
rect 6972 18572 6978 18584
rect 7009 18581 7021 18584
rect 7055 18581 7067 18615
rect 8294 18612 8300 18624
rect 8255 18584 8300 18612
rect 7009 18575 7067 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 9861 18615 9919 18621
rect 9861 18612 9873 18615
rect 9732 18584 9873 18612
rect 9732 18572 9738 18584
rect 9861 18581 9873 18584
rect 9907 18581 9919 18615
rect 12066 18612 12072 18624
rect 12027 18584 12072 18612
rect 9861 18575 9919 18581
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2866 18408 2872 18420
rect 2827 18380 2872 18408
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3234 18408 3240 18420
rect 3195 18380 3240 18408
rect 3234 18368 3240 18380
rect 3292 18368 3298 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6236 18380 6561 18408
rect 6236 18368 6242 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 6549 18371 6607 18377
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7561 18411 7619 18417
rect 7561 18408 7573 18411
rect 7524 18380 7573 18408
rect 7524 18368 7530 18380
rect 7561 18377 7573 18380
rect 7607 18377 7619 18411
rect 8662 18408 8668 18420
rect 8623 18380 8668 18408
rect 7561 18371 7619 18377
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9214 18408 9220 18420
rect 9175 18380 9220 18408
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 12253 18411 12311 18417
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 12434 18408 12440 18420
rect 12299 18380 12440 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 2501 18275 2559 18281
rect 2501 18272 2513 18275
rect 1412 18244 2513 18272
rect 1412 18216 1440 18244
rect 2501 18241 2513 18244
rect 2547 18241 2559 18275
rect 2501 18235 2559 18241
rect 8205 18275 8263 18281
rect 8205 18241 8217 18275
rect 8251 18272 8263 18275
rect 8680 18272 8708 18368
rect 10781 18343 10839 18349
rect 10781 18340 10793 18343
rect 9692 18312 10793 18340
rect 9692 18284 9720 18312
rect 10781 18309 10793 18312
rect 10827 18309 10839 18343
rect 10781 18303 10839 18309
rect 9674 18272 9680 18284
rect 8251 18244 8708 18272
rect 9635 18244 9680 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 11425 18275 11483 18281
rect 9907 18244 10364 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 1394 18204 1400 18216
rect 1355 18176 1400 18204
rect 1394 18164 1400 18176
rect 1452 18164 1458 18216
rect 1762 18164 1768 18216
rect 1820 18204 1826 18216
rect 2685 18207 2743 18213
rect 2685 18204 2697 18207
rect 1820 18176 2697 18204
rect 1820 18164 1826 18176
rect 2685 18173 2697 18176
rect 2731 18204 2743 18207
rect 2774 18204 2780 18216
rect 2731 18176 2780 18204
rect 2731 18173 2743 18176
rect 2685 18167 2743 18173
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18204 3847 18207
rect 3878 18204 3884 18216
rect 3835 18176 3884 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 4062 18145 4068 18148
rect 1673 18139 1731 18145
rect 1673 18105 1685 18139
rect 1719 18105 1731 18139
rect 1673 18099 1731 18105
rect 3697 18139 3755 18145
rect 3697 18105 3709 18139
rect 3743 18136 3755 18139
rect 4034 18139 4068 18145
rect 4034 18136 4046 18139
rect 3743 18108 4046 18136
rect 3743 18105 3755 18108
rect 3697 18099 3755 18105
rect 4034 18105 4046 18108
rect 4120 18136 4126 18148
rect 7929 18139 7987 18145
rect 7929 18136 7941 18139
rect 4120 18108 4182 18136
rect 7024 18108 7941 18136
rect 4034 18099 4068 18105
rect 1688 18068 1716 18099
rect 4062 18096 4068 18099
rect 4120 18096 4126 18108
rect 1762 18068 1768 18080
rect 1688 18040 1768 18068
rect 1762 18028 1768 18040
rect 1820 18028 1826 18080
rect 2225 18071 2283 18077
rect 2225 18037 2237 18071
rect 2271 18068 2283 18071
rect 2314 18068 2320 18080
rect 2271 18040 2320 18068
rect 2271 18037 2283 18040
rect 2225 18031 2283 18037
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 5166 18068 5172 18080
rect 5127 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 5810 18068 5816 18080
rect 5771 18040 5816 18068
rect 5810 18028 5816 18040
rect 5868 18068 5874 18080
rect 6089 18071 6147 18077
rect 6089 18068 6101 18071
rect 5868 18040 6101 18068
rect 5868 18028 5874 18040
rect 6089 18037 6101 18040
rect 6135 18037 6147 18071
rect 6089 18031 6147 18037
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 7024 18077 7052 18108
rect 7929 18105 7941 18108
rect 7975 18105 7987 18139
rect 7929 18099 7987 18105
rect 7009 18071 7067 18077
rect 7009 18068 7021 18071
rect 6972 18040 7021 18068
rect 6972 18028 6978 18040
rect 7009 18037 7021 18040
rect 7055 18037 7067 18071
rect 7009 18031 7067 18037
rect 7469 18071 7527 18077
rect 7469 18037 7481 18071
rect 7515 18068 7527 18071
rect 8018 18068 8024 18080
rect 7515 18040 8024 18068
rect 7515 18037 7527 18040
rect 7469 18031 7527 18037
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9582 18068 9588 18080
rect 9171 18040 9588 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10336 18077 10364 18244
rect 11425 18241 11437 18275
rect 11471 18272 11483 18275
rect 11514 18272 11520 18284
rect 11471 18244 11520 18272
rect 11471 18241 11483 18244
rect 11425 18235 11483 18241
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 10735 18108 11284 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 11256 18080 11284 18108
rect 10321 18071 10379 18077
rect 10321 18037 10333 18071
rect 10367 18068 10379 18071
rect 10962 18068 10968 18080
rect 10367 18040 10968 18068
rect 10367 18037 10379 18040
rect 10321 18031 10379 18037
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11146 18068 11152 18080
rect 11107 18040 11152 18068
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 11296 18040 11341 18068
rect 11296 18028 11302 18040
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11572 18040 11805 18068
rect 11572 18028 11578 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3237 17867 3295 17873
rect 3237 17864 3249 17867
rect 2832 17836 3249 17864
rect 2832 17824 2838 17836
rect 3237 17833 3249 17836
rect 3283 17833 3295 17867
rect 3237 17827 3295 17833
rect 3786 17824 3792 17876
rect 3844 17864 3850 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3844 17836 4077 17864
rect 3844 17824 3850 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 5166 17864 5172 17876
rect 4479 17836 4752 17864
rect 5127 17836 5172 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 4212 17768 4660 17796
rect 4212 17756 4218 17768
rect 2038 17688 2044 17740
rect 2096 17728 2102 17740
rect 2225 17731 2283 17737
rect 2225 17728 2237 17731
rect 2096 17700 2237 17728
rect 2096 17688 2102 17700
rect 2225 17697 2237 17700
rect 2271 17728 2283 17731
rect 2869 17731 2927 17737
rect 2869 17728 2881 17731
rect 2271 17700 2881 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 2869 17697 2881 17700
rect 2915 17697 2927 17731
rect 2869 17691 2927 17697
rect 4632 17672 4660 17768
rect 4724 17728 4752 17836
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 7193 17867 7251 17873
rect 7193 17833 7205 17867
rect 7239 17864 7251 17867
rect 7282 17864 7288 17876
rect 7239 17836 7288 17864
rect 7239 17833 7251 17836
rect 7193 17827 7251 17833
rect 7282 17824 7288 17836
rect 7340 17864 7346 17876
rect 7742 17864 7748 17876
rect 7340 17836 7748 17864
rect 7340 17824 7346 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 9953 17867 10011 17873
rect 9953 17864 9965 17867
rect 9732 17836 9965 17864
rect 9732 17824 9738 17836
rect 9953 17833 9965 17836
rect 9999 17833 10011 17867
rect 9953 17827 10011 17833
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 12345 17867 12403 17873
rect 12345 17864 12357 17867
rect 11112 17836 12357 17864
rect 11112 17824 11118 17836
rect 12345 17833 12357 17836
rect 12391 17833 12403 17867
rect 12345 17827 12403 17833
rect 6086 17805 6092 17808
rect 6080 17796 6092 17805
rect 6047 17768 6092 17796
rect 6080 17759 6092 17768
rect 6086 17756 6092 17759
rect 6144 17756 6150 17808
rect 12434 17796 12440 17808
rect 10980 17768 12440 17796
rect 5166 17728 5172 17740
rect 4724 17700 5172 17728
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 9030 17688 9036 17740
rect 9088 17728 9094 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 9088 17700 9505 17728
rect 9088 17688 9094 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 2314 17660 2320 17672
rect 2275 17632 2320 17660
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17629 2467 17663
rect 2409 17623 2467 17629
rect 2130 17552 2136 17604
rect 2188 17592 2194 17604
rect 2424 17592 2452 17623
rect 4338 17620 4344 17672
rect 4396 17660 4402 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4396 17632 4537 17660
rect 4396 17620 4402 17632
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 4525 17623 4583 17629
rect 4614 17620 4620 17672
rect 4672 17660 4678 17672
rect 5810 17660 5816 17672
rect 4672 17632 4765 17660
rect 5723 17632 5816 17660
rect 4672 17620 4678 17632
rect 5810 17620 5816 17632
rect 5868 17620 5874 17672
rect 8294 17660 8300 17672
rect 8255 17632 8300 17660
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 10686 17660 10692 17672
rect 10428 17632 10692 17660
rect 2188 17564 2452 17592
rect 2188 17552 2194 17564
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 1854 17524 1860 17536
rect 1815 17496 1860 17524
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 3697 17527 3755 17533
rect 3697 17493 3709 17527
rect 3743 17524 3755 17527
rect 5442 17524 5448 17536
rect 3743 17496 5448 17524
rect 3743 17493 3755 17496
rect 3697 17487 3755 17493
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5629 17527 5687 17533
rect 5629 17524 5641 17527
rect 5592 17496 5641 17524
rect 5592 17484 5598 17496
rect 5629 17493 5641 17496
rect 5675 17493 5687 17527
rect 5828 17524 5856 17620
rect 6730 17524 6736 17536
rect 5828 17496 6736 17524
rect 5629 17487 5687 17493
rect 6730 17484 6736 17496
rect 6788 17524 6794 17536
rect 7374 17524 7380 17536
rect 6788 17496 7380 17524
rect 6788 17484 6794 17496
rect 7374 17484 7380 17496
rect 7432 17524 7438 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7432 17496 8125 17524
rect 7432 17484 7438 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 8202 17484 8208 17536
rect 8260 17524 8266 17536
rect 8757 17527 8815 17533
rect 8757 17524 8769 17527
rect 8260 17496 8769 17524
rect 8260 17484 8266 17496
rect 8757 17493 8769 17496
rect 8803 17524 8815 17527
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 8803 17496 9137 17524
rect 8803 17493 8815 17496
rect 8757 17487 8815 17493
rect 9125 17493 9137 17496
rect 9171 17524 9183 17527
rect 9309 17527 9367 17533
rect 9309 17524 9321 17527
rect 9171 17496 9321 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9309 17493 9321 17496
rect 9355 17524 9367 17527
rect 9490 17524 9496 17536
rect 9355 17496 9496 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9490 17484 9496 17496
rect 9548 17524 9554 17536
rect 10428 17533 10456 17632
rect 10686 17620 10692 17632
rect 10744 17660 10750 17672
rect 10980 17669 11008 17768
rect 12434 17756 12440 17768
rect 12492 17756 12498 17808
rect 11232 17731 11290 17737
rect 11232 17697 11244 17731
rect 11278 17728 11290 17731
rect 11514 17728 11520 17740
rect 11278 17700 11520 17728
rect 11278 17697 11290 17700
rect 11232 17691 11290 17697
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 10965 17663 11023 17669
rect 10965 17660 10977 17663
rect 10744 17632 10977 17660
rect 10744 17620 10750 17632
rect 10965 17629 10977 17632
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 10413 17527 10471 17533
rect 10413 17524 10425 17527
rect 9548 17496 10425 17524
rect 9548 17484 9554 17496
rect 10413 17493 10425 17496
rect 10459 17493 10471 17527
rect 10778 17524 10784 17536
rect 10739 17496 10784 17524
rect 10413 17487 10471 17493
rect 10778 17484 10784 17496
rect 10836 17524 10842 17536
rect 11146 17524 11152 17536
rect 10836 17496 11152 17524
rect 10836 17484 10842 17496
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17320 4583 17323
rect 4614 17320 4620 17332
rect 4571 17292 4620 17320
rect 4571 17289 4583 17292
rect 4525 17283 4583 17289
rect 4614 17280 4620 17292
rect 4672 17320 4678 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 4672 17292 5457 17320
rect 4672 17280 4678 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 6086 17280 6092 17332
rect 6144 17320 6150 17332
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 6144 17292 6193 17320
rect 6144 17280 6150 17292
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6181 17283 6239 17289
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 10873 17323 10931 17329
rect 10873 17320 10885 17323
rect 9732 17292 10885 17320
rect 9732 17280 9738 17292
rect 10873 17289 10885 17292
rect 10919 17289 10931 17323
rect 11514 17320 11520 17332
rect 11427 17292 11520 17320
rect 10873 17283 10931 17289
rect 11514 17280 11520 17292
rect 11572 17320 11578 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 11572 17292 13829 17320
rect 11572 17280 11578 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 13817 17283 13875 17289
rect 1670 17144 1676 17196
rect 1728 17184 1734 17196
rect 2041 17187 2099 17193
rect 2041 17184 2053 17187
rect 1728 17156 2053 17184
rect 1728 17144 1734 17156
rect 2041 17153 2053 17156
rect 2087 17153 2099 17187
rect 2041 17147 2099 17153
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 6641 17187 6699 17193
rect 2188 17156 2233 17184
rect 2188 17144 2194 17156
rect 6641 17153 6653 17187
rect 6687 17184 6699 17187
rect 9490 17184 9496 17196
rect 6687 17156 7144 17184
rect 9451 17156 9496 17184
rect 6687 17153 6699 17156
rect 6641 17147 6699 17153
rect 2590 17076 2596 17128
rect 2648 17116 2654 17128
rect 3145 17119 3203 17125
rect 3145 17116 3157 17119
rect 2648 17088 3157 17116
rect 2648 17076 2654 17088
rect 3145 17085 3157 17088
rect 3191 17116 3203 17119
rect 3878 17116 3884 17128
rect 3191 17088 3884 17116
rect 3191 17085 3203 17088
rect 3145 17079 3203 17085
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5592 17088 5641 17116
rect 5592 17076 5598 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17085 7067 17119
rect 7116 17116 7144 17156
rect 9490 17144 9496 17156
rect 9548 17144 9554 17196
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17184 11943 17187
rect 12434 17184 12440 17196
rect 11931 17156 12440 17184
rect 11931 17153 11943 17156
rect 11885 17147 11943 17153
rect 12434 17144 12440 17156
rect 12492 17184 12498 17196
rect 12492 17156 12585 17184
rect 12492 17144 12498 17156
rect 7282 17125 7288 17128
rect 7276 17116 7288 17125
rect 7116 17088 7288 17116
rect 7009 17079 7067 17085
rect 7276 17079 7288 17088
rect 3050 17048 3056 17060
rect 2963 17020 3056 17048
rect 3050 17008 3056 17020
rect 3108 17048 3114 17060
rect 3390 17051 3448 17057
rect 3390 17048 3402 17051
rect 3108 17020 3402 17048
rect 3108 17008 3114 17020
rect 3390 17017 3402 17020
rect 3436 17017 3448 17051
rect 3390 17011 3448 17017
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 1670 16980 1676 16992
rect 1627 16952 1676 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 2593 16983 2651 16989
rect 2593 16980 2605 16983
rect 2188 16952 2605 16980
rect 2188 16940 2194 16952
rect 2593 16949 2605 16952
rect 2639 16949 2651 16983
rect 5166 16980 5172 16992
rect 5127 16952 5172 16980
rect 2593 16943 2651 16949
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 5810 16980 5816 16992
rect 5771 16952 5816 16980
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 7024 16980 7052 17079
rect 7282 17076 7288 17079
rect 7340 17076 7346 17128
rect 9309 17051 9367 17057
rect 9309 17048 9321 17051
rect 8404 17020 9321 17048
rect 8404 16992 8432 17020
rect 9309 17017 9321 17020
rect 9355 17048 9367 17051
rect 9738 17051 9796 17057
rect 9738 17048 9750 17051
rect 9355 17020 9750 17048
rect 9355 17017 9367 17020
rect 9309 17011 9367 17017
rect 9738 17017 9750 17020
rect 9784 17017 9796 17051
rect 9738 17011 9796 17017
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 10836 17020 12265 17048
rect 10836 17008 10842 17020
rect 12253 17017 12265 17020
rect 12299 17048 12311 17051
rect 12618 17048 12624 17060
rect 12299 17020 12624 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12618 17008 12624 17020
rect 12676 17057 12682 17060
rect 12676 17051 12740 17057
rect 12676 17017 12694 17051
rect 12728 17017 12740 17051
rect 12676 17011 12740 17017
rect 12676 17008 12682 17011
rect 7282 16980 7288 16992
rect 7024 16952 7288 16980
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 8386 16980 8392 16992
rect 8347 16952 8392 16980
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2406 16776 2412 16788
rect 2367 16748 2412 16776
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 4617 16779 4675 16785
rect 4617 16776 4629 16779
rect 4304 16748 4629 16776
rect 4304 16736 4310 16748
rect 4617 16745 4629 16748
rect 4663 16745 4675 16779
rect 4617 16739 4675 16745
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 5905 16779 5963 16785
rect 5905 16776 5917 16779
rect 5500 16748 5917 16776
rect 5500 16736 5506 16748
rect 5905 16745 5917 16748
rect 5951 16776 5963 16779
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5951 16748 6009 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 5997 16745 6009 16748
rect 6043 16745 6055 16779
rect 5997 16739 6055 16745
rect 6181 16779 6239 16785
rect 6181 16745 6193 16779
rect 6227 16776 6239 16779
rect 6822 16776 6828 16788
rect 6227 16748 6828 16776
rect 6227 16745 6239 16748
rect 6181 16739 6239 16745
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 8297 16779 8355 16785
rect 8297 16776 8309 16779
rect 7616 16748 8309 16776
rect 7616 16736 7622 16748
rect 8297 16745 8309 16748
rect 8343 16776 8355 16779
rect 9122 16776 9128 16788
rect 8343 16748 9128 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 10045 16779 10103 16785
rect 10045 16745 10057 16779
rect 10091 16776 10103 16779
rect 10134 16776 10140 16788
rect 10091 16748 10140 16776
rect 10091 16745 10103 16748
rect 10045 16739 10103 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 1397 16711 1455 16717
rect 1397 16677 1409 16711
rect 1443 16708 1455 16711
rect 2682 16708 2688 16720
rect 1443 16680 2688 16708
rect 1443 16677 1455 16680
rect 1397 16671 1455 16677
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 2869 16711 2927 16717
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 3786 16708 3792 16720
rect 2915 16680 3556 16708
rect 3747 16680 3792 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 3528 16652 3556 16680
rect 3786 16668 3792 16680
rect 3844 16668 3850 16720
rect 4890 16668 4896 16720
rect 4948 16708 4954 16720
rect 5077 16711 5135 16717
rect 5077 16708 5089 16711
rect 4948 16680 5089 16708
rect 4948 16668 4954 16680
rect 5077 16677 5089 16680
rect 5123 16677 5135 16711
rect 5077 16671 5135 16677
rect 6086 16668 6092 16720
rect 6144 16708 6150 16720
rect 7837 16711 7895 16717
rect 6144 16680 6776 16708
rect 6144 16668 6150 16680
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2130 16600 2136 16652
rect 2188 16640 2194 16652
rect 2225 16643 2283 16649
rect 2225 16640 2237 16643
rect 2188 16612 2237 16640
rect 2188 16600 2194 16612
rect 2225 16609 2237 16612
rect 2271 16609 2283 16643
rect 2225 16603 2283 16609
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 3510 16640 3516 16652
rect 2832 16612 2877 16640
rect 3471 16612 3516 16640
rect 2832 16600 2838 16612
rect 3510 16600 3516 16612
rect 3568 16600 3574 16652
rect 4338 16640 4344 16652
rect 4299 16612 4344 16640
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 4522 16600 4528 16652
rect 4580 16640 4586 16652
rect 4985 16643 5043 16649
rect 4985 16640 4997 16643
rect 4580 16612 4997 16640
rect 4580 16600 4586 16612
rect 4985 16609 4997 16612
rect 5031 16609 5043 16643
rect 4985 16603 5043 16609
rect 5721 16643 5779 16649
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 5994 16640 6000 16652
rect 5767 16612 6000 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 6546 16640 6552 16652
rect 6507 16612 6552 16640
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6748 16584 6776 16680
rect 7837 16677 7849 16711
rect 7883 16708 7895 16711
rect 8386 16708 8392 16720
rect 7883 16680 8392 16708
rect 7883 16677 7895 16680
rect 7837 16671 7895 16677
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 12434 16708 12440 16720
rect 11256 16680 12440 16708
rect 8404 16640 8432 16668
rect 11256 16649 11284 16680
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 11241 16643 11299 16649
rect 8404 16612 8524 16640
rect 2682 16532 2688 16584
rect 2740 16572 2746 16584
rect 3050 16572 3056 16584
rect 2740 16544 3056 16572
rect 2740 16532 2746 16544
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 5166 16572 5172 16584
rect 5127 16544 5172 16572
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 6638 16572 6644 16584
rect 6599 16544 6644 16572
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 6730 16532 6736 16584
rect 6788 16572 6794 16584
rect 6788 16544 6881 16572
rect 6788 16532 6794 16544
rect 8018 16532 8024 16584
rect 8076 16572 8082 16584
rect 8496 16581 8524 16612
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11508 16643 11566 16649
rect 11508 16609 11520 16643
rect 11554 16640 11566 16643
rect 11882 16640 11888 16652
rect 11554 16612 11888 16640
rect 11554 16609 11566 16612
rect 11508 16603 11566 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 8389 16575 8447 16581
rect 8389 16572 8401 16575
rect 8076 16544 8401 16572
rect 8076 16532 8082 16544
rect 8389 16541 8401 16544
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 9033 16575 9091 16581
rect 9033 16541 9045 16575
rect 9079 16572 9091 16575
rect 9490 16572 9496 16584
rect 9079 16544 9496 16572
rect 9079 16541 9091 16544
rect 9033 16535 9091 16541
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 9950 16532 9956 16584
rect 10008 16572 10014 16584
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 10008 16544 10149 16572
rect 10008 16532 10014 16544
rect 10137 16541 10149 16544
rect 10183 16541 10195 16575
rect 10137 16535 10195 16541
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 10244 16504 10272 16535
rect 9416 16476 10272 16504
rect 9416 16448 9444 16476
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16436 5963 16439
rect 6086 16436 6092 16448
rect 5951 16408 6092 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 7282 16436 7288 16448
rect 7243 16408 7288 16436
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 7926 16436 7932 16448
rect 7887 16408 7932 16436
rect 7926 16396 7932 16408
rect 7984 16396 7990 16448
rect 9398 16436 9404 16448
rect 9359 16408 9404 16436
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 9674 16436 9680 16448
rect 9635 16408 9680 16436
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11057 16439 11115 16445
rect 11057 16436 11069 16439
rect 11020 16408 11069 16436
rect 11020 16396 11026 16408
rect 11057 16405 11069 16408
rect 11103 16405 11115 16439
rect 11057 16399 11115 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2041 16235 2099 16241
rect 2041 16201 2053 16235
rect 2087 16232 2099 16235
rect 2682 16232 2688 16244
rect 2087 16204 2688 16232
rect 2087 16201 2099 16204
rect 2041 16195 2099 16201
rect 2682 16192 2688 16204
rect 2740 16232 2746 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 2740 16204 3893 16232
rect 2740 16192 2746 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 4982 16232 4988 16244
rect 4943 16204 4988 16232
rect 3881 16195 3939 16201
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 7558 16232 7564 16244
rect 7519 16204 7564 16232
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16232 10563 16235
rect 10686 16232 10692 16244
rect 10551 16204 10692 16232
rect 10551 16201 10563 16204
rect 10505 16195 10563 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12621 16235 12679 16241
rect 12621 16232 12633 16235
rect 12492 16204 12633 16232
rect 12492 16192 12498 16204
rect 12621 16201 12633 16204
rect 12667 16201 12679 16235
rect 12621 16195 12679 16201
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 10321 16167 10379 16173
rect 10321 16164 10333 16167
rect 10284 16136 10333 16164
rect 10284 16124 10290 16136
rect 10321 16133 10333 16136
rect 10367 16133 10379 16167
rect 10321 16127 10379 16133
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16096 5687 16099
rect 5994 16096 6000 16108
rect 5675 16068 6000 16096
rect 5675 16065 5687 16068
rect 5629 16059 5687 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 6822 16096 6828 16108
rect 6783 16068 6828 16096
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10836 16068 11069 16096
rect 10836 16056 10842 16068
rect 11057 16065 11069 16068
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1762 16028 1768 16040
rect 1443 16000 1768 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 2590 16028 2596 16040
rect 2547 16000 2596 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 2590 15988 2596 16000
rect 2648 15988 2654 16040
rect 2768 16031 2826 16037
rect 2768 15997 2780 16031
rect 2814 15997 2826 16031
rect 2768 15991 2826 15997
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 16028 8079 16031
rect 8110 16028 8116 16040
rect 8067 16000 8116 16028
rect 8067 15997 8079 16000
rect 8021 15991 8079 15997
rect 2682 15920 2688 15972
rect 2740 15960 2746 15972
rect 2792 15960 2820 15991
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 8288 16031 8346 16037
rect 8288 15997 8300 16031
rect 8334 16028 8346 16031
rect 8570 16028 8576 16040
rect 8334 16000 8576 16028
rect 8334 15997 8346 16000
rect 8288 15991 8346 15997
rect 8570 15988 8576 16000
rect 8628 16028 8634 16040
rect 9582 16028 9588 16040
rect 8628 16000 9588 16028
rect 8628 15988 8634 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 5353 15963 5411 15969
rect 5353 15960 5365 15963
rect 2740 15932 2820 15960
rect 4816 15932 5365 15960
rect 2740 15920 2746 15932
rect 4816 15904 4844 15932
rect 5353 15929 5365 15932
rect 5399 15929 5411 15963
rect 5353 15923 5411 15929
rect 6273 15963 6331 15969
rect 6273 15929 6285 15963
rect 6319 15960 6331 15963
rect 6638 15960 6644 15972
rect 6319 15932 6644 15960
rect 6319 15929 6331 15932
rect 6273 15923 6331 15929
rect 6638 15920 6644 15932
rect 6696 15960 6702 15972
rect 7190 15960 7196 15972
rect 6696 15932 7196 15960
rect 6696 15920 6702 15932
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 2406 15892 2412 15904
rect 2367 15864 2412 15892
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5258 15852 5264 15904
rect 5316 15892 5322 15904
rect 5445 15895 5503 15901
rect 5445 15892 5457 15895
rect 5316 15864 5457 15892
rect 5316 15852 5322 15864
rect 5445 15861 5457 15864
rect 5491 15861 5503 15895
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 5445 15855 5503 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15892 7987 15895
rect 8018 15892 8024 15904
rect 7975 15864 8024 15892
rect 7975 15861 7987 15864
rect 7929 15855 7987 15861
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 9398 15892 9404 15904
rect 8904 15864 9404 15892
rect 8904 15852 8910 15864
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 9950 15892 9956 15904
rect 9911 15864 9956 15892
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10870 15892 10876 15904
rect 10831 15864 10876 15892
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 10962 15852 10968 15904
rect 11020 15892 11026 15904
rect 11020 15864 11065 15892
rect 11020 15852 11026 15864
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11204 15864 11529 15892
rect 11204 15852 11210 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 2041 15691 2099 15697
rect 2041 15688 2053 15691
rect 1912 15660 2053 15688
rect 1912 15648 1918 15660
rect 2041 15657 2053 15660
rect 2087 15657 2099 15691
rect 6730 15688 6736 15700
rect 6691 15660 6736 15688
rect 2041 15651 2099 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7466 15688 7472 15700
rect 7427 15660 7472 15688
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 7926 15688 7932 15700
rect 7887 15660 7932 15688
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 8570 15688 8576 15700
rect 8531 15660 8576 15688
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 9953 15691 10011 15697
rect 9953 15657 9965 15691
rect 9999 15688 10011 15691
rect 10597 15691 10655 15697
rect 10597 15688 10609 15691
rect 9999 15660 10609 15688
rect 9999 15657 10011 15660
rect 9953 15651 10011 15657
rect 10597 15657 10609 15660
rect 10643 15688 10655 15691
rect 10870 15688 10876 15700
rect 10643 15660 10876 15688
rect 10643 15657 10655 15660
rect 10597 15651 10655 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11940 15660 12357 15688
rect 11940 15648 11946 15660
rect 12345 15657 12357 15660
rect 12391 15688 12403 15691
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12391 15660 12909 15688
rect 12391 15657 12403 15660
rect 12345 15651 12403 15657
rect 12897 15657 12909 15660
rect 12943 15688 12955 15691
rect 12986 15688 12992 15700
rect 12943 15660 12992 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 13998 15688 14004 15700
rect 13959 15660 14004 15688
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 1670 15580 1676 15632
rect 1728 15620 1734 15632
rect 1949 15623 2007 15629
rect 1949 15620 1961 15623
rect 1728 15592 1961 15620
rect 1728 15580 1734 15592
rect 1949 15589 1961 15592
rect 1995 15589 2007 15623
rect 1949 15583 2007 15589
rect 7650 15580 7656 15632
rect 7708 15620 7714 15632
rect 7837 15623 7895 15629
rect 7837 15620 7849 15623
rect 7708 15592 7849 15620
rect 7708 15580 7714 15592
rect 7837 15589 7849 15592
rect 7883 15620 7895 15623
rect 8202 15620 8208 15632
rect 7883 15592 8208 15620
rect 7883 15589 7895 15592
rect 7837 15583 7895 15589
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 11146 15580 11152 15632
rect 11204 15629 11210 15632
rect 11204 15623 11268 15629
rect 11204 15589 11222 15623
rect 11256 15589 11268 15623
rect 11204 15583 11268 15589
rect 11204 15580 11210 15583
rect 4982 15561 4988 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4976 15552 4988 15561
rect 4663 15524 4988 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4976 15515 4988 15524
rect 4982 15512 4988 15515
rect 5040 15512 5046 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 7024 15524 7389 15552
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15484 2283 15487
rect 2961 15487 3019 15493
rect 2961 15484 2973 15487
rect 2271 15456 2973 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2961 15453 2973 15456
rect 3007 15484 3019 15487
rect 3418 15484 3424 15496
rect 3007 15456 3424 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 3878 15484 3884 15496
rect 3839 15456 3884 15484
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 4706 15484 4712 15496
rect 4667 15456 4712 15484
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 2682 15416 2688 15428
rect 2595 15388 2688 15416
rect 2682 15376 2688 15388
rect 2740 15416 2746 15428
rect 4246 15416 4252 15428
rect 2740 15388 4252 15416
rect 2740 15376 2746 15388
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3329 15351 3387 15357
rect 3329 15348 3341 15351
rect 2832 15320 3341 15348
rect 2832 15308 2838 15320
rect 3329 15317 3341 15320
rect 3375 15317 3387 15351
rect 3329 15311 3387 15317
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 5408 15320 6101 15348
rect 5408 15308 5414 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7024 15357 7052 15524
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 7377 15515 7435 15521
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 9364 15524 9505 15552
rect 9364 15512 9370 15524
rect 9493 15521 9505 15524
rect 9539 15521 9551 15555
rect 9493 15515 9551 15521
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 10870 15552 10876 15564
rect 9732 15524 10876 15552
rect 9732 15512 9738 15524
rect 10870 15512 10876 15524
rect 10928 15552 10934 15564
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 10928 15524 10977 15552
rect 10928 15512 10934 15524
rect 10965 15521 10977 15524
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 8110 15484 8116 15496
rect 8023 15456 8116 15484
rect 8110 15444 8116 15456
rect 8168 15484 8174 15496
rect 8570 15484 8576 15496
rect 8168 15456 8576 15484
rect 8168 15444 8174 15456
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 7193 15419 7251 15425
rect 7193 15385 7205 15419
rect 7239 15416 7251 15419
rect 7282 15416 7288 15428
rect 7239 15388 7288 15416
rect 7239 15385 7251 15388
rect 7193 15379 7251 15385
rect 7282 15376 7288 15388
rect 7340 15416 7346 15428
rect 8202 15416 8208 15428
rect 7340 15388 8208 15416
rect 7340 15376 7346 15388
rect 8202 15376 8208 15388
rect 8260 15376 8266 15428
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 6972 15320 7021 15348
rect 6972 15308 6978 15320
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 8846 15348 8852 15360
rect 8807 15320 8852 15348
rect 7009 15311 7067 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 9088 15320 9321 15348
rect 9088 15308 9094 15320
rect 9309 15317 9321 15320
rect 9355 15348 9367 15351
rect 9398 15348 9404 15360
rect 9355 15320 9404 15348
rect 9355 15317 9367 15320
rect 9309 15311 9367 15317
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 3568 15116 3893 15144
rect 3568 15104 3574 15116
rect 3881 15113 3893 15116
rect 3927 15113 3939 15147
rect 7650 15144 7656 15156
rect 7611 15116 7656 15144
rect 3881 15107 3939 15113
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 8021 15147 8079 15153
rect 8021 15113 8033 15147
rect 8067 15144 8079 15147
rect 8110 15144 8116 15156
rect 8067 15116 8116 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 9490 15144 9496 15156
rect 9451 15116 9496 15144
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 10192 15116 10609 15144
rect 10192 15104 10198 15116
rect 10597 15113 10609 15116
rect 10643 15113 10655 15147
rect 10597 15107 10655 15113
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12492 15116 12537 15144
rect 12492 15104 12498 15116
rect 6546 15076 6552 15088
rect 6507 15048 6552 15076
rect 6546 15036 6552 15048
rect 6604 15036 6610 15088
rect 13998 15036 14004 15088
rect 14056 15076 14062 15088
rect 14056 15048 14596 15076
rect 14056 15036 14062 15048
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 4525 15011 4583 15017
rect 4525 15008 4537 15011
rect 4304 14980 4537 15008
rect 4304 14968 4310 14980
rect 4525 14977 4537 14980
rect 4571 15008 4583 15011
rect 4614 15008 4620 15020
rect 4571 14980 4620 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4614 14968 4620 14980
rect 4672 15008 4678 15020
rect 5350 15008 5356 15020
rect 4672 14980 5356 15008
rect 4672 14968 4678 14980
rect 5350 14968 5356 14980
rect 5408 14968 5414 15020
rect 7098 15008 7104 15020
rect 7059 14980 7104 15008
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 15008 10195 15011
rect 11146 15008 11152 15020
rect 10183 14980 11152 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 11146 14968 11152 14980
rect 11204 15008 11210 15020
rect 12434 15008 12440 15020
rect 11204 14980 12440 15008
rect 11204 14968 11210 14980
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 12986 15008 12992 15020
rect 12544 14980 12848 15008
rect 12947 14980 12992 15008
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 1949 14943 2007 14949
rect 1949 14940 1961 14943
rect 1820 14912 1961 14940
rect 1820 14900 1826 14912
rect 1949 14909 1961 14912
rect 1995 14940 2007 14943
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 1995 14912 2513 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2501 14909 2513 14912
rect 2547 14940 2559 14943
rect 3789 14943 3847 14949
rect 2547 14912 3464 14940
rect 2547 14909 2559 14912
rect 2501 14903 2559 14909
rect 2406 14872 2412 14884
rect 2367 14844 2412 14872
rect 2406 14832 2412 14844
rect 2464 14832 2470 14884
rect 3436 14881 3464 14912
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 4341 14943 4399 14949
rect 4341 14940 4353 14943
rect 3835 14912 4353 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4341 14909 4353 14912
rect 4387 14940 4399 14943
rect 4890 14940 4896 14952
rect 4387 14912 4896 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5442 14940 5448 14952
rect 5403 14912 5448 14940
rect 5442 14900 5448 14912
rect 5500 14940 5506 14952
rect 6181 14943 6239 14949
rect 6181 14940 6193 14943
rect 5500 14912 6193 14940
rect 5500 14900 5506 14912
rect 6181 14909 6193 14912
rect 6227 14909 6239 14943
rect 8110 14940 8116 14952
rect 8071 14912 8116 14940
rect 6181 14903 6239 14909
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 8380 14943 8438 14949
rect 8380 14909 8392 14943
rect 8426 14940 8438 14943
rect 8846 14940 8852 14952
rect 8426 14912 8852 14940
rect 8426 14909 8438 14912
rect 8380 14903 8438 14909
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 3421 14875 3479 14881
rect 3421 14841 3433 14875
rect 3467 14872 3479 14875
rect 4798 14872 4804 14884
rect 3467 14844 4804 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 4264 14813 4292 14844
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 5718 14872 5724 14884
rect 5679 14844 5724 14872
rect 5718 14832 5724 14844
rect 5776 14832 5782 14884
rect 8128 14872 8156 14900
rect 9582 14872 9588 14884
rect 8128 14844 9588 14872
rect 9582 14832 9588 14844
rect 9640 14832 9646 14884
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 10505 14875 10563 14881
rect 10505 14872 10517 14875
rect 10192 14844 10517 14872
rect 10192 14832 10198 14844
rect 10505 14841 10517 14844
rect 10551 14872 10563 14875
rect 10965 14875 11023 14881
rect 10965 14872 10977 14875
rect 10551 14844 10977 14872
rect 10551 14841 10563 14844
rect 10505 14835 10563 14841
rect 10965 14841 10977 14844
rect 11011 14841 11023 14875
rect 11882 14872 11888 14884
rect 11795 14844 11888 14872
rect 10965 14835 11023 14841
rect 11882 14832 11888 14844
rect 11940 14872 11946 14884
rect 12544 14872 12572 14980
rect 12820 14949 12848 14980
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 13814 15008 13820 15020
rect 13775 14980 13820 15008
rect 13814 14968 13820 14980
rect 13872 15008 13878 15020
rect 14568 15017 14596 15048
rect 14553 15011 14611 15017
rect 13872 14980 14412 15008
rect 13872 14968 13878 14980
rect 14384 14949 14412 14980
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 11940 14844 12572 14872
rect 11940 14832 11946 14844
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 14461 14875 14519 14881
rect 14461 14872 14473 14875
rect 14148 14844 14473 14872
rect 14148 14832 14154 14844
rect 14461 14841 14473 14844
rect 14507 14841 14519 14875
rect 14461 14835 14519 14841
rect 4249 14807 4307 14813
rect 4249 14773 4261 14807
rect 4295 14773 4307 14807
rect 4982 14804 4988 14816
rect 4943 14776 4988 14804
rect 4249 14767 4307 14773
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5258 14804 5264 14816
rect 5219 14776 5264 14804
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 11054 14804 11060 14816
rect 11015 14776 11060 14804
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 12158 14804 12164 14816
rect 12119 14776 12164 14804
rect 12158 14764 12164 14776
rect 12216 14804 12222 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12216 14776 12909 14804
rect 12216 14764 12222 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 13446 14804 13452 14816
rect 13407 14776 13452 14804
rect 12897 14767 12955 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 14001 14807 14059 14813
rect 14001 14804 14013 14807
rect 13964 14776 14013 14804
rect 13964 14764 13970 14776
rect 14001 14773 14013 14776
rect 14047 14773 14059 14807
rect 14001 14767 14059 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1394 14600 1400 14612
rect 1355 14572 1400 14600
rect 1394 14560 1400 14572
rect 1452 14560 1458 14612
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 1728 14572 2053 14600
rect 1728 14560 1734 14572
rect 2041 14569 2053 14572
rect 2087 14600 2099 14603
rect 2406 14600 2412 14612
rect 2087 14572 2412 14600
rect 2087 14569 2099 14572
rect 2041 14563 2099 14569
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 2866 14600 2872 14612
rect 2823 14572 2872 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 4120 14572 4261 14600
rect 4120 14560 4126 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4614 14600 4620 14612
rect 4575 14572 4620 14600
rect 4249 14563 4307 14569
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 5040 14572 6653 14600
rect 5040 14560 5046 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 6641 14563 6699 14569
rect 7561 14603 7619 14609
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 7926 14600 7932 14612
rect 7607 14572 7932 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8846 14600 8852 14612
rect 8759 14572 8852 14600
rect 8846 14560 8852 14572
rect 8904 14600 8910 14612
rect 9490 14600 9496 14612
rect 8904 14572 9496 14600
rect 8904 14560 8910 14572
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10134 14600 10140 14612
rect 10091 14572 10140 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 13998 14600 14004 14612
rect 12492 14572 12537 14600
rect 13959 14572 14004 14600
rect 12492 14560 12498 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 2682 14532 2688 14544
rect 2188 14504 2688 14532
rect 2188 14492 2194 14504
rect 2682 14492 2688 14504
rect 2740 14532 2746 14544
rect 3421 14535 3479 14541
rect 3421 14532 3433 14535
rect 2740 14504 3433 14532
rect 2740 14492 2746 14504
rect 3421 14501 3433 14504
rect 3467 14501 3479 14535
rect 3421 14495 3479 14501
rect 9953 14535 10011 14541
rect 9953 14501 9965 14535
rect 9999 14532 10011 14535
rect 11054 14532 11060 14544
rect 9999 14504 11060 14532
rect 9999 14501 10011 14504
rect 9953 14495 10011 14501
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 3881 14467 3939 14473
rect 3881 14433 3893 14467
rect 3927 14464 3939 14467
rect 4062 14464 4068 14476
rect 3927 14436 4068 14464
rect 3927 14433 3939 14436
rect 3881 14427 3939 14433
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 5534 14473 5540 14476
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 4212 14436 4997 14464
rect 4212 14424 4218 14436
rect 4985 14433 4997 14436
rect 5031 14433 5043 14467
rect 5528 14464 5540 14473
rect 5495 14436 5540 14464
rect 4985 14427 5043 14433
rect 5528 14427 5540 14436
rect 5534 14424 5540 14427
rect 5592 14424 5598 14476
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 8113 14467 8171 14473
rect 8113 14464 8125 14467
rect 7340 14436 8125 14464
rect 7340 14424 7346 14436
rect 8113 14433 8125 14436
rect 8159 14464 8171 14467
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 8159 14436 10609 14464
rect 8159 14433 8171 14436
rect 8113 14427 8171 14433
rect 10597 14433 10609 14436
rect 10643 14464 10655 14467
rect 10962 14464 10968 14476
rect 10643 14436 10968 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 11324 14467 11382 14473
rect 11324 14433 11336 14467
rect 11370 14464 11382 14467
rect 11698 14464 11704 14476
rect 11370 14436 11704 14464
rect 11370 14433 11382 14436
rect 11324 14427 11382 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 23382 14464 23388 14476
rect 23343 14436 23388 14464
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 2038 14356 2044 14408
rect 2096 14396 2102 14408
rect 2869 14399 2927 14405
rect 2869 14396 2881 14399
rect 2096 14368 2881 14396
rect 2096 14356 2102 14368
rect 2869 14365 2881 14368
rect 2915 14365 2927 14399
rect 3050 14396 3056 14408
rect 3011 14368 3056 14396
rect 2869 14359 2927 14365
rect 2884 14328 2912 14359
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 5166 14396 5172 14408
rect 4764 14368 5172 14396
rect 4764 14356 4770 14368
rect 5166 14356 5172 14368
rect 5224 14396 5230 14408
rect 5261 14399 5319 14405
rect 5261 14396 5273 14399
rect 5224 14368 5273 14396
rect 5224 14356 5230 14368
rect 5261 14365 5273 14368
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 8205 14399 8263 14405
rect 8205 14396 8217 14399
rect 7432 14368 8217 14396
rect 7432 14356 7438 14368
rect 8205 14365 8217 14368
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 5074 14328 5080 14340
rect 2884 14300 5080 14328
rect 5074 14288 5080 14300
rect 5132 14288 5138 14340
rect 7742 14328 7748 14340
rect 7703 14300 7748 14328
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 8312 14328 8340 14359
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 10928 14368 11069 14396
rect 10928 14356 10934 14368
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 7892 14300 8340 14328
rect 7892 14288 7898 14300
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 9306 14260 9312 14272
rect 9267 14232 9312 14260
rect 9306 14220 9312 14232
rect 9364 14260 9370 14272
rect 9674 14260 9680 14272
rect 9364 14232 9680 14260
rect 9364 14220 9370 14232
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 23569 14263 23627 14269
rect 23569 14229 23581 14263
rect 23615 14260 23627 14263
rect 24946 14260 24952 14272
rect 23615 14232 24952 14260
rect 23615 14229 23627 14232
rect 23569 14223 23627 14229
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14056 1731 14059
rect 2866 14056 2872 14068
rect 1719 14028 2872 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 11054 14056 11060 14068
rect 10643 14028 11060 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 23382 14056 23388 14068
rect 23343 14028 23388 14056
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 2038 13988 2044 14000
rect 1999 13960 2044 13988
rect 2038 13948 2044 13960
rect 2096 13948 2102 14000
rect 3418 13948 3424 14000
rect 3476 13988 3482 14000
rect 3513 13991 3571 13997
rect 3513 13988 3525 13991
rect 3476 13960 3525 13988
rect 3476 13948 3482 13960
rect 3513 13957 3525 13960
rect 3559 13957 3571 13991
rect 3513 13951 3571 13957
rect 4430 13948 4436 14000
rect 4488 13988 4494 14000
rect 4617 13991 4675 13997
rect 4617 13988 4629 13991
rect 4488 13960 4629 13988
rect 4488 13948 4494 13960
rect 4617 13957 4629 13960
rect 4663 13957 4675 13991
rect 4617 13951 4675 13957
rect 7282 13948 7288 14000
rect 7340 13988 7346 14000
rect 7377 13991 7435 13997
rect 7377 13988 7389 13991
rect 7340 13960 7389 13988
rect 7340 13948 7346 13960
rect 7377 13957 7389 13960
rect 7423 13957 7435 13991
rect 7377 13951 7435 13957
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 11977 13991 12035 13997
rect 11977 13988 11989 13991
rect 10744 13960 11989 13988
rect 10744 13948 10750 13960
rect 11977 13957 11989 13960
rect 12023 13988 12035 13991
rect 12621 13991 12679 13997
rect 12621 13988 12633 13991
rect 12023 13960 12633 13988
rect 12023 13957 12035 13960
rect 11977 13951 12035 13957
rect 12621 13957 12633 13960
rect 12667 13988 12679 13991
rect 13446 13988 13452 14000
rect 12667 13960 13452 13988
rect 12667 13957 12679 13960
rect 12621 13951 12679 13957
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 23845 13991 23903 13997
rect 23845 13957 23857 13991
rect 23891 13988 23903 13991
rect 24854 13988 24860 14000
rect 23891 13960 24860 13988
rect 23891 13957 23903 13960
rect 23845 13951 23903 13957
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 4571 13892 5181 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 8110 13920 8116 13932
rect 8071 13892 8116 13920
rect 5169 13883 5227 13889
rect 2130 13852 2136 13864
rect 2091 13824 2136 13852
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 2866 13852 2872 13864
rect 2740 13824 2872 13852
rect 2740 13812 2746 13824
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 5184 13852 5212 13883
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 11241 13923 11299 13929
rect 11241 13920 11253 13923
rect 10183 13892 11253 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 11241 13889 11253 13892
rect 11287 13920 11299 13923
rect 11698 13920 11704 13932
rect 11287 13892 11704 13920
rect 11287 13889 11299 13892
rect 11241 13883 11299 13889
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 5442 13852 5448 13864
rect 5184 13824 5448 13852
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5552 13824 6009 13852
rect 2400 13787 2458 13793
rect 2400 13753 2412 13787
rect 2446 13753 2458 13787
rect 4982 13784 4988 13796
rect 4943 13756 4988 13784
rect 2400 13747 2458 13753
rect 2424 13716 2452 13747
rect 4982 13744 4988 13756
rect 5040 13784 5046 13796
rect 5552 13784 5580 13824
rect 5997 13821 6009 13824
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 6641 13855 6699 13861
rect 6641 13852 6653 13855
rect 6604 13824 6653 13852
rect 6604 13812 6610 13824
rect 6641 13821 6653 13824
rect 6687 13821 6699 13855
rect 6914 13852 6920 13864
rect 6641 13815 6699 13821
rect 6840 13824 6920 13852
rect 6840 13784 6868 13824
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 7374 13812 7380 13864
rect 7432 13852 7438 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7432 13824 7757 13852
rect 7432 13812 7438 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 8380 13855 8438 13861
rect 8380 13821 8392 13855
rect 8426 13852 8438 13855
rect 8846 13852 8852 13864
rect 8426 13824 8852 13852
rect 8426 13821 8438 13824
rect 8380 13815 8438 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10870 13852 10876 13864
rect 10551 13824 10876 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10870 13812 10876 13824
rect 10928 13852 10934 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 10928 13824 11069 13852
rect 10928 13812 10934 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 11057 13815 11115 13821
rect 23658 13812 23664 13824
rect 23716 13852 23722 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23716 13824 24225 13852
rect 23716 13812 23722 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 10962 13784 10968 13796
rect 5040 13756 5580 13784
rect 6472 13756 6868 13784
rect 10923 13756 10968 13784
rect 5040 13744 5046 13756
rect 6472 13728 6500 13756
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 2682 13716 2688 13728
rect 2424 13688 2688 13716
rect 2682 13676 2688 13688
rect 2740 13676 2746 13728
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 3108 13688 4169 13716
rect 3108 13676 3114 13688
rect 4157 13685 4169 13688
rect 4203 13716 4215 13719
rect 4430 13716 4436 13728
rect 4203 13688 4436 13716
rect 4203 13685 4215 13688
rect 4157 13679 4215 13685
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 5077 13719 5135 13725
rect 5077 13685 5089 13719
rect 5123 13716 5135 13719
rect 5258 13716 5264 13728
rect 5123 13688 5264 13716
rect 5123 13685 5135 13688
rect 5077 13679 5135 13685
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 6454 13716 6460 13728
rect 6415 13688 6460 13716
rect 6454 13676 6460 13688
rect 6512 13676 6518 13728
rect 6822 13716 6828 13728
rect 6783 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 9490 13716 9496 13728
rect 9451 13688 9496 13716
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 11698 13716 11704 13728
rect 11659 13688 11704 13716
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2866 13512 2872 13524
rect 2827 13484 2872 13512
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 6825 13515 6883 13521
rect 6825 13512 6837 13515
rect 5776 13484 6837 13512
rect 5776 13472 5782 13484
rect 6825 13481 6837 13484
rect 6871 13512 6883 13515
rect 7834 13512 7840 13524
rect 6871 13484 7840 13512
rect 6871 13481 6883 13484
rect 6825 13475 6883 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 10413 13515 10471 13521
rect 10413 13512 10425 13515
rect 9732 13484 10425 13512
rect 9732 13472 9738 13484
rect 10413 13481 10425 13484
rect 10459 13481 10471 13515
rect 10413 13475 10471 13481
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11756 13484 12081 13512
rect 11756 13472 11762 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 1756 13447 1814 13453
rect 1756 13413 1768 13447
rect 1802 13444 1814 13447
rect 2590 13444 2596 13456
rect 1802 13416 2596 13444
rect 1802 13413 1814 13416
rect 1756 13407 1814 13413
rect 2590 13404 2596 13416
rect 2648 13444 2654 13456
rect 3050 13444 3056 13456
rect 2648 13416 3056 13444
rect 2648 13404 2654 13416
rect 3050 13404 3056 13416
rect 3108 13444 3114 13456
rect 3421 13447 3479 13453
rect 3421 13444 3433 13447
rect 3108 13416 3433 13444
rect 3108 13404 3114 13416
rect 3421 13413 3433 13416
rect 3467 13413 3479 13447
rect 5258 13444 5264 13456
rect 5219 13416 5264 13444
rect 3421 13407 3479 13413
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 6362 13404 6368 13456
rect 6420 13444 6426 13456
rect 7650 13444 7656 13456
rect 6420 13416 7656 13444
rect 6420 13404 6426 13416
rect 7650 13404 7656 13416
rect 7708 13444 7714 13456
rect 8389 13447 8447 13453
rect 8389 13444 8401 13447
rect 7708 13416 8401 13444
rect 7708 13404 7714 13416
rect 8389 13413 8401 13416
rect 8435 13444 8447 13447
rect 8570 13444 8576 13456
rect 8435 13416 8576 13444
rect 8435 13413 8447 13416
rect 8389 13407 8447 13413
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 11422 13444 11428 13456
rect 10612 13416 11428 13444
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13376 1547 13379
rect 1578 13376 1584 13388
rect 1535 13348 1584 13376
rect 1535 13345 1547 13348
rect 1489 13339 1547 13345
rect 1578 13336 1584 13348
rect 1636 13376 1642 13388
rect 2130 13376 2136 13388
rect 1636 13348 2136 13376
rect 1636 13336 1642 13348
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 4065 13379 4123 13385
rect 4065 13376 4077 13379
rect 2832 13348 4077 13376
rect 2832 13336 2838 13348
rect 4065 13345 4077 13348
rect 4111 13376 4123 13379
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4111 13348 4813 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 5166 13336 5172 13388
rect 5224 13376 5230 13388
rect 5445 13379 5503 13385
rect 5445 13376 5457 13379
rect 5224 13348 5457 13376
rect 5224 13336 5230 13348
rect 5445 13345 5457 13348
rect 5491 13345 5503 13379
rect 5445 13339 5503 13345
rect 5712 13379 5770 13385
rect 5712 13345 5724 13379
rect 5758 13376 5770 13379
rect 5994 13376 6000 13388
rect 5758 13348 6000 13376
rect 5758 13345 5770 13348
rect 5712 13339 5770 13345
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 10612 13385 10640 13416
rect 11422 13404 11428 13416
rect 11480 13404 11486 13456
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 10778 13336 10784 13388
rect 10836 13376 10842 13388
rect 10945 13379 11003 13385
rect 10945 13376 10957 13379
rect 10836 13348 10957 13376
rect 10836 13336 10842 13348
rect 10945 13345 10957 13348
rect 10991 13345 11003 13379
rect 22370 13376 22376 13388
rect 22331 13348 22376 13376
rect 10945 13339 11003 13345
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13308 4399 13311
rect 5350 13308 5356 13320
rect 4387 13280 5356 13308
rect 4387 13277 4399 13280
rect 4341 13271 4399 13277
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 8478 13308 8484 13320
rect 8439 13280 8484 13308
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 10686 13308 10692 13320
rect 10647 13280 10692 13308
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 7834 13200 7840 13252
rect 7892 13240 7898 13252
rect 8941 13243 8999 13249
rect 8941 13240 8953 13243
rect 7892 13212 8953 13240
rect 7892 13200 7898 13212
rect 8941 13209 8953 13212
rect 8987 13240 8999 13243
rect 10229 13243 10287 13249
rect 10229 13240 10241 13243
rect 8987 13212 10241 13240
rect 8987 13209 8999 13212
rect 8941 13203 8999 13209
rect 10229 13209 10241 13212
rect 10275 13209 10287 13243
rect 10229 13203 10287 13209
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 2590 13172 2596 13184
rect 1820 13144 2596 13172
rect 1820 13132 1826 13144
rect 2590 13132 2596 13144
rect 2648 13132 2654 13184
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 3970 13172 3976 13184
rect 3927 13144 3976 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7926 13172 7932 13184
rect 7887 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9398 13172 9404 13184
rect 9359 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 9861 13175 9919 13181
rect 9861 13172 9873 13175
rect 9824 13144 9873 13172
rect 9824 13132 9830 13144
rect 9861 13141 9873 13144
rect 9907 13141 9919 13175
rect 10244 13172 10272 13203
rect 11882 13172 11888 13184
rect 10244 13144 11888 13172
rect 9861 13135 9919 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 22557 13175 22615 13181
rect 22557 13141 22569 13175
rect 22603 13172 22615 13175
rect 23474 13172 23480 13184
rect 22603 13144 23480 13172
rect 22603 13141 22615 13144
rect 22557 13135 22615 13141
rect 23474 13132 23480 13144
rect 23532 13132 23538 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1854 12968 1860 12980
rect 1815 12940 1860 12968
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 2130 12928 2136 12980
rect 2188 12968 2194 12980
rect 4062 12968 4068 12980
rect 2188 12940 4068 12968
rect 2188 12928 2194 12940
rect 2866 12900 2872 12912
rect 2424 12872 2872 12900
rect 2424 12841 2452 12872
rect 2866 12860 2872 12872
rect 2924 12900 2930 12912
rect 3237 12903 3295 12909
rect 3237 12900 3249 12903
rect 2924 12872 3249 12900
rect 2924 12860 2930 12872
rect 3237 12869 3249 12872
rect 3283 12869 3295 12903
rect 3237 12863 3295 12869
rect 3427 12841 3455 12940
rect 4062 12928 4068 12940
rect 4120 12968 4126 12980
rect 5534 12968 5540 12980
rect 4120 12940 5540 12968
rect 4120 12928 4126 12940
rect 5534 12928 5540 12940
rect 5592 12968 5598 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5592 12940 5917 12968
rect 5592 12928 5598 12940
rect 5905 12937 5917 12940
rect 5951 12968 5963 12971
rect 6086 12968 6092 12980
rect 5951 12940 6092 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6546 12968 6552 12980
rect 6507 12940 6552 12968
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7064 12940 7665 12968
rect 7064 12928 7070 12940
rect 7653 12937 7665 12940
rect 7699 12937 7711 12971
rect 7653 12931 7711 12937
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 8628 12940 8677 12968
rect 8628 12928 8634 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 8665 12931 8723 12937
rect 8846 12928 8852 12980
rect 8904 12968 8910 12980
rect 9401 12971 9459 12977
rect 9401 12968 9413 12971
rect 8904 12940 9413 12968
rect 8904 12928 8910 12940
rect 9401 12937 9413 12940
rect 9447 12937 9459 12971
rect 12618 12968 12624 12980
rect 12579 12940 12624 12968
rect 9401 12931 9459 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 7469 12903 7527 12909
rect 7469 12900 7481 12903
rect 5132 12872 7481 12900
rect 5132 12860 5138 12872
rect 7469 12869 7481 12872
rect 7515 12900 7527 12903
rect 8294 12900 8300 12912
rect 7515 12872 8300 12900
rect 7515 12869 7527 12872
rect 7469 12863 7527 12869
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 10778 12900 10784 12912
rect 10060 12872 10784 12900
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12832 7251 12835
rect 8110 12832 8116 12844
rect 7239 12804 8116 12832
rect 7239 12801 7251 12804
rect 7193 12795 7251 12801
rect 8110 12792 8116 12804
rect 8168 12832 8174 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 8168 12804 8217 12832
rect 8168 12792 8174 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 10060 12841 10088 12872
rect 10778 12860 10784 12872
rect 10836 12900 10842 12912
rect 10962 12900 10968 12912
rect 10836 12872 10968 12900
rect 10836 12860 10842 12872
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 9732 12804 10057 12832
rect 9732 12792 9738 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 11940 12804 12173 12832
rect 11940 12792 11946 12804
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 3677 12767 3735 12773
rect 3677 12764 3689 12767
rect 3568 12736 3689 12764
rect 3568 12724 3574 12736
rect 3677 12733 3689 12736
rect 3723 12733 3735 12767
rect 3677 12727 3735 12733
rect 5810 12724 5816 12776
rect 5868 12764 5874 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5868 12736 6101 12764
rect 5868 12724 5874 12736
rect 6089 12733 6101 12736
rect 6135 12764 6147 12767
rect 6454 12764 6460 12776
rect 6135 12736 6460 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 8021 12767 8079 12773
rect 8021 12764 8033 12767
rect 7524 12736 8033 12764
rect 7524 12724 7530 12736
rect 8021 12733 8033 12736
rect 8067 12733 8079 12767
rect 11146 12764 11152 12776
rect 11059 12736 11152 12764
rect 8021 12727 8079 12733
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 22370 12764 22376 12776
rect 22331 12736 22376 12764
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 2225 12699 2283 12705
rect 2225 12665 2237 12699
rect 2271 12696 2283 12699
rect 2961 12699 3019 12705
rect 2961 12696 2973 12699
rect 2271 12668 2973 12696
rect 2271 12665 2283 12668
rect 2225 12659 2283 12665
rect 2961 12665 2973 12668
rect 3007 12696 3019 12699
rect 3142 12696 3148 12708
rect 3007 12668 3148 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 5537 12699 5595 12705
rect 5537 12665 5549 12699
rect 5583 12696 5595 12699
rect 5994 12696 6000 12708
rect 5583 12668 6000 12696
rect 5583 12665 5595 12668
rect 5537 12659 5595 12665
rect 5994 12656 6000 12668
rect 6052 12696 6058 12708
rect 6822 12696 6828 12708
rect 6052 12668 6828 12696
rect 6052 12656 6058 12668
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 9214 12656 9220 12708
rect 9272 12696 9278 12708
rect 9309 12699 9367 12705
rect 9309 12696 9321 12699
rect 9272 12668 9321 12696
rect 9272 12656 9278 12668
rect 9309 12665 9321 12668
rect 9355 12696 9367 12699
rect 9769 12699 9827 12705
rect 9769 12696 9781 12699
rect 9355 12668 9781 12696
rect 9355 12665 9367 12668
rect 9309 12659 9367 12665
rect 9769 12665 9781 12668
rect 9815 12665 9827 12699
rect 11164 12696 11192 12724
rect 11885 12699 11943 12705
rect 11885 12696 11897 12699
rect 11164 12668 11897 12696
rect 9769 12659 9827 12665
rect 11885 12665 11897 12668
rect 11931 12665 11943 12699
rect 11885 12659 11943 12665
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 2130 12628 2136 12640
rect 1811 12600 2136 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 2130 12588 2136 12600
rect 2188 12628 2194 12640
rect 2317 12631 2375 12637
rect 2317 12628 2329 12631
rect 2188 12600 2329 12628
rect 2188 12588 2194 12600
rect 2317 12597 2329 12600
rect 2363 12597 2375 12631
rect 2317 12591 2375 12597
rect 4522 12588 4528 12640
rect 4580 12628 4586 12640
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 4580 12600 4813 12628
rect 4580 12588 4586 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8202 12628 8208 12640
rect 8159 12600 8208 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 9398 12628 9404 12640
rect 8904 12600 9404 12628
rect 8904 12588 8910 12600
rect 9398 12588 9404 12600
rect 9456 12628 9462 12640
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 9456 12600 9873 12628
rect 9456 12588 9462 12600
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10744 12600 10977 12628
rect 10744 12588 10750 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 11422 12628 11428 12640
rect 11383 12600 11428 12628
rect 10965 12591 11023 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 12989 12631 13047 12637
rect 12989 12628 13001 12631
rect 12400 12600 13001 12628
rect 12400 12588 12406 12600
rect 12989 12597 13001 12600
rect 13035 12628 13047 12631
rect 13357 12631 13415 12637
rect 13357 12628 13369 12631
rect 13035 12600 13369 12628
rect 13035 12597 13047 12600
rect 12989 12591 13047 12597
rect 13357 12597 13369 12600
rect 13403 12628 13415 12631
rect 14182 12628 14188 12640
rect 13403 12600 14188 12628
rect 13403 12597 13415 12600
rect 13357 12591 13415 12597
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 2682 12424 2688 12436
rect 1443 12396 2688 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 2958 12424 2964 12436
rect 2919 12396 2964 12424
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3418 12424 3424 12436
rect 3379 12396 3424 12424
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 5810 12424 5816 12436
rect 5771 12396 5816 12424
rect 5810 12384 5816 12396
rect 5868 12384 5874 12436
rect 6104 12396 6215 12424
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 6104 12356 6132 12396
rect 6187 12365 6215 12396
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 6972 12396 7297 12424
rect 6972 12384 6978 12396
rect 7285 12393 7297 12396
rect 7331 12393 7343 12427
rect 7285 12387 7343 12393
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 7616 12396 8033 12424
rect 7616 12384 7622 12396
rect 8021 12393 8033 12396
rect 8067 12424 8079 12427
rect 8478 12424 8484 12436
rect 8067 12396 8484 12424
rect 8067 12393 8079 12396
rect 8021 12387 8079 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 9214 12424 9220 12436
rect 8619 12396 9220 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11333 12427 11391 12433
rect 11333 12424 11345 12427
rect 11112 12396 11345 12424
rect 11112 12384 11118 12396
rect 11333 12393 11345 12396
rect 11379 12393 11391 12427
rect 11333 12387 11391 12393
rect 2924 12328 6132 12356
rect 6172 12359 6230 12365
rect 2924 12316 2930 12328
rect 6172 12325 6184 12359
rect 6218 12356 6230 12359
rect 6270 12356 6276 12368
rect 6218 12328 6276 12356
rect 6218 12325 6230 12328
rect 6172 12319 6230 12325
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 10686 12356 10692 12368
rect 9968 12328 10692 12356
rect 1762 12288 1768 12300
rect 1723 12260 1768 12288
rect 1762 12248 1768 12260
rect 1820 12248 1826 12300
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 2774 12288 2780 12300
rect 1903 12260 2780 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4212 12260 4721 12288
rect 4212 12248 4218 12260
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 4856 12260 4901 12288
rect 4856 12248 4862 12260
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 5534 12288 5540 12300
rect 5408 12260 5540 12288
rect 5408 12248 5414 12260
rect 5534 12248 5540 12260
rect 5592 12288 5598 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5592 12260 5917 12288
rect 5592 12248 5598 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 9582 12288 9588 12300
rect 9539 12260 9588 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 9968 12297 9996 12328
rect 10686 12316 10692 12328
rect 10744 12316 10750 12368
rect 9953 12291 10011 12297
rect 9953 12257 9965 12291
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10209 12291 10267 12297
rect 10209 12288 10221 12291
rect 10100 12260 10221 12288
rect 10100 12248 10106 12260
rect 10209 12257 10221 12260
rect 10255 12257 10267 12291
rect 10704 12288 10732 12316
rect 12710 12297 12716 12300
rect 12704 12288 12716 12297
rect 10704 12260 11928 12288
rect 12671 12260 12716 12288
rect 10209 12251 10267 12257
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 4816 12220 4844 12248
rect 3927 12192 4844 12220
rect 4985 12223 5043 12229
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5074 12220 5080 12232
rect 5031 12192 5080 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 10060 12220 10088 12248
rect 9171 12192 10088 12220
rect 11900 12220 11928 12260
rect 12704 12251 12716 12260
rect 12710 12248 12716 12251
rect 12768 12248 12774 12300
rect 21818 12288 21824 12300
rect 21779 12260 21824 12288
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 12342 12220 12348 12232
rect 11900 12192 12348 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 12342 12180 12348 12192
rect 12400 12220 12406 12232
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 12400 12192 12449 12220
rect 12400 12180 12406 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 4338 12152 4344 12164
rect 4299 12124 4344 12152
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12084 2651 12087
rect 2866 12084 2872 12096
rect 2639 12056 2872 12084
rect 2639 12053 2651 12056
rect 2593 12047 2651 12053
rect 2866 12044 2872 12056
rect 2924 12084 2930 12096
rect 3142 12084 3148 12096
rect 2924 12056 3148 12084
rect 2924 12044 2930 12056
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 5445 12087 5503 12093
rect 5445 12053 5457 12087
rect 5491 12084 5503 12087
rect 6546 12084 6552 12096
rect 5491 12056 6552 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 8386 12084 8392 12096
rect 8347 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11940 12056 11989 12084
rect 11940 12044 11946 12056
rect 11977 12053 11989 12056
rect 12023 12084 12035 12087
rect 12342 12084 12348 12096
rect 12023 12056 12348 12084
rect 12023 12053 12035 12056
rect 11977 12047 12035 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 13817 12087 13875 12093
rect 13817 12053 13829 12087
rect 13863 12084 13875 12087
rect 13906 12084 13912 12096
rect 13863 12056 13912 12084
rect 13863 12053 13875 12056
rect 13817 12047 13875 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 22002 12084 22008 12096
rect 21963 12056 22008 12084
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1486 11840 1492 11892
rect 1544 11880 1550 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1544 11852 1593 11880
rect 1544 11840 1550 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 1581 11843 1639 11849
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 2314 11840 2320 11892
rect 2372 11880 2378 11892
rect 2501 11883 2559 11889
rect 2501 11880 2513 11883
rect 2372 11852 2513 11880
rect 2372 11840 2378 11852
rect 2501 11849 2513 11852
rect 2547 11849 2559 11883
rect 2501 11843 2559 11849
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5500 11852 5641 11880
rect 5500 11840 5506 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 6270 11880 6276 11892
rect 6231 11852 6276 11880
rect 5629 11843 5687 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 8444 11852 10609 11880
rect 8444 11840 8450 11852
rect 10597 11849 10609 11852
rect 10643 11849 10655 11883
rect 10597 11843 10655 11849
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12710 11880 12716 11892
rect 12299 11852 12716 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 12492 11784 12537 11812
rect 12492 11772 12498 11784
rect 3050 11744 3056 11756
rect 3011 11716 3056 11744
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 4120 11716 4261 11744
rect 4120 11704 4126 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 7834 11744 7840 11756
rect 5408 11716 7840 11744
rect 5408 11704 5414 11716
rect 7834 11704 7840 11716
rect 7892 11744 7898 11756
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7892 11716 8125 11744
rect 7892 11704 7898 11716
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 10686 11744 10692 11756
rect 9456 11716 10692 11744
rect 9456 11704 9462 11716
rect 10686 11704 10692 11716
rect 10744 11744 10750 11756
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 10744 11716 11161 11744
rect 10744 11704 10750 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 11848 11716 12909 11744
rect 11848 11704 11854 11716
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13262 11744 13268 11756
rect 13127 11716 13268 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 8380 11679 8438 11685
rect 8380 11645 8392 11679
rect 8426 11676 8438 11679
rect 9416 11676 9444 11704
rect 8426 11648 9444 11676
rect 8426 11645 8438 11648
rect 8380 11639 8438 11645
rect 2409 11611 2467 11617
rect 2409 11577 2421 11611
rect 2455 11608 2467 11611
rect 2958 11608 2964 11620
rect 2455 11580 2964 11608
rect 2455 11577 2467 11580
rect 2409 11571 2467 11577
rect 2958 11568 2964 11580
rect 3016 11568 3022 11620
rect 4522 11617 4528 11620
rect 3789 11611 3847 11617
rect 3789 11577 3801 11611
rect 3835 11608 3847 11611
rect 3835 11580 4476 11608
rect 3835 11577 3847 11580
rect 3789 11571 3847 11577
rect 2866 11540 2872 11552
rect 2827 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 4154 11540 4160 11552
rect 4115 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4448 11540 4476 11580
rect 4516 11571 4528 11617
rect 4580 11608 4586 11620
rect 7653 11611 7711 11617
rect 4580 11580 4616 11608
rect 4522 11568 4528 11571
rect 4580 11568 4586 11580
rect 7653 11577 7665 11611
rect 7699 11608 7711 11611
rect 8021 11611 8079 11617
rect 8021 11608 8033 11611
rect 7699 11580 8033 11608
rect 7699 11577 7711 11580
rect 7653 11571 7711 11577
rect 8021 11577 8033 11580
rect 8067 11608 8079 11611
rect 8395 11608 8423 11639
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 10134 11676 10140 11688
rect 9916 11648 10140 11676
rect 9916 11636 9922 11648
rect 10134 11636 10140 11648
rect 10192 11676 10198 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10192 11648 10977 11676
rect 10192 11636 10198 11648
rect 10965 11645 10977 11648
rect 11011 11676 11023 11679
rect 21818 11676 21824 11688
rect 11011 11648 13032 11676
rect 21779 11648 21824 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 8478 11608 8484 11620
rect 8067 11580 8484 11608
rect 8067 11577 8079 11580
rect 8021 11571 8079 11577
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 5074 11540 5080 11552
rect 4448 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 6546 11540 6552 11552
rect 6507 11512 6552 11540
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 7098 11540 7104 11552
rect 7059 11512 7104 11540
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 8168 11512 9505 11540
rect 8168 11500 8174 11512
rect 9493 11509 9505 11512
rect 9539 11540 9551 11543
rect 9858 11540 9864 11552
rect 9539 11512 9864 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10870 11540 10876 11552
rect 10551 11512 10876 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 10870 11500 10876 11512
rect 10928 11540 10934 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10928 11512 11069 11540
rect 10928 11500 10934 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 11057 11503 11115 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12805 11543 12863 11549
rect 12805 11509 12817 11543
rect 12851 11540 12863 11543
rect 13004 11540 13032 11648
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 12851 11512 13461 11540
rect 12851 11509 12863 11512
rect 12805 11503 12863 11509
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3050 11336 3056 11348
rect 2915 11308 3056 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3050 11296 3056 11308
rect 3108 11336 3114 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3108 11308 3433 11336
rect 3108 11296 3114 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 4985 11339 5043 11345
rect 4985 11336 4997 11339
rect 4580 11308 4997 11336
rect 4580 11296 4586 11308
rect 4985 11305 4997 11308
rect 5031 11336 5043 11339
rect 5810 11336 5816 11348
rect 5031 11308 5816 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6328 11308 6837 11336
rect 6328 11296 6334 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7156 11308 7757 11336
rect 7156 11296 7162 11308
rect 7745 11305 7757 11308
rect 7791 11336 7803 11339
rect 8297 11339 8355 11345
rect 8297 11336 8309 11339
rect 7791 11308 8309 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8297 11305 8309 11308
rect 8343 11305 8355 11339
rect 8297 11299 8355 11305
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 9858 11336 9864 11348
rect 8444 11308 8489 11336
rect 9819 11308 9864 11336
rect 8444 11296 8450 11308
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 10686 11336 10692 11348
rect 10367 11308 10692 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 11112 11308 12265 11336
rect 11112 11296 11118 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12618 11336 12624 11348
rect 12579 11308 12624 11336
rect 12253 11299 12311 11305
rect 12618 11296 12624 11308
rect 12676 11336 12682 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 12676 11308 13645 11336
rect 12676 11296 12682 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 3789 11271 3847 11277
rect 3789 11268 3801 11271
rect 1452 11240 3801 11268
rect 1452 11228 1458 11240
rect 3789 11237 3801 11240
rect 3835 11268 3847 11271
rect 4433 11271 4491 11277
rect 4433 11268 4445 11271
rect 3835 11240 4445 11268
rect 3835 11237 3847 11240
rect 3789 11231 3847 11237
rect 4433 11237 4445 11240
rect 4479 11237 4491 11271
rect 4433 11231 4491 11237
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 5690 11271 5748 11277
rect 5690 11268 5702 11271
rect 5592 11240 5702 11268
rect 5592 11228 5598 11240
rect 5690 11237 5702 11240
rect 5736 11237 5748 11271
rect 5690 11231 5748 11237
rect 7469 11271 7527 11277
rect 7469 11237 7481 11271
rect 7515 11268 7527 11271
rect 7558 11268 7564 11280
rect 7515 11240 7564 11268
rect 7515 11237 7527 11240
rect 7469 11231 7527 11237
rect 7558 11228 7564 11240
rect 7616 11228 7622 11280
rect 11238 11228 11244 11280
rect 11296 11268 11302 11280
rect 13170 11268 13176 11280
rect 11296 11240 13176 11268
rect 11296 11228 11302 11240
rect 13170 11228 13176 11240
rect 13228 11228 13234 11280
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11200 1547 11203
rect 1578 11200 1584 11212
rect 1535 11172 1584 11200
rect 1535 11169 1547 11172
rect 1489 11163 1547 11169
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 1756 11203 1814 11209
rect 1756 11169 1768 11203
rect 1802 11200 1814 11203
rect 2038 11200 2044 11212
rect 1802 11172 2044 11200
rect 1802 11169 1814 11172
rect 1756 11163 1814 11169
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 4154 11200 4160 11212
rect 4115 11172 4160 11200
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 5445 11203 5503 11209
rect 5445 11200 5457 11203
rect 5408 11172 5457 11200
rect 5408 11160 5414 11172
rect 5445 11169 5457 11172
rect 5491 11169 5503 11203
rect 5445 11163 5503 11169
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10778 11200 10784 11212
rect 10459 11172 10784 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 8478 11132 8484 11144
rect 8439 11104 8484 11132
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 11422 11132 11428 11144
rect 9640 11104 11428 11132
rect 9640 11092 9646 11104
rect 11422 11092 11428 11104
rect 11480 11132 11486 11144
rect 12710 11132 12716 11144
rect 11480 11104 11744 11132
rect 12671 11104 12716 11132
rect 11480 11092 11486 11104
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 2924 11036 5396 11064
rect 2924 11024 2930 11036
rect 5258 10996 5264 11008
rect 5219 10968 5264 10996
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 5368 10996 5396 11036
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 7524 11036 7941 11064
rect 7524 11024 7530 11036
rect 7929 11033 7941 11036
rect 7975 11033 7987 11067
rect 7929 11027 7987 11033
rect 9401 11067 9459 11073
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 9490 11064 9496 11076
rect 9447 11036 9496 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 9490 11024 9496 11036
rect 9548 11064 9554 11076
rect 10042 11064 10048 11076
rect 9548 11036 10048 11064
rect 9548 11024 9554 11036
rect 10042 11024 10048 11036
rect 10100 11064 10106 11076
rect 11716 11073 11744 11104
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13262 11132 13268 11144
rect 12860 11104 12905 11132
rect 13223 11104 13268 11132
rect 12860 11092 12866 11104
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 11701 11067 11759 11073
rect 10100 11036 11100 11064
rect 10100 11024 10106 11036
rect 11072 11008 11100 11036
rect 11701 11033 11713 11067
rect 11747 11033 11759 11067
rect 11701 11027 11759 11033
rect 9033 10999 9091 11005
rect 9033 10996 9045 10999
rect 5368 10968 9045 10996
rect 9033 10965 9045 10968
rect 9079 10996 9091 10999
rect 9214 10996 9220 11008
rect 9079 10968 9220 10996
rect 9079 10965 9091 10968
rect 9033 10959 9091 10965
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 6546 10792 6552 10804
rect 6319 10764 6552 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 5626 10684 5632 10736
rect 5684 10724 5690 10736
rect 6288 10724 6316 10755
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 8846 10792 8852 10804
rect 8807 10764 8852 10792
rect 8846 10752 8852 10764
rect 8904 10752 8910 10804
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12342 10792 12348 10804
rect 12299 10764 12348 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12342 10752 12348 10764
rect 12400 10792 12406 10804
rect 12802 10792 12808 10804
rect 12400 10764 12808 10792
rect 12400 10752 12406 10764
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 5684 10696 6316 10724
rect 5684 10684 5690 10696
rect 2498 10656 2504 10668
rect 2411 10628 2504 10656
rect 2498 10616 2504 10628
rect 2556 10656 2562 10668
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 2556 10628 3249 10656
rect 2556 10616 2562 10628
rect 3237 10625 3249 10628
rect 3283 10656 3295 10659
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3283 10628 3709 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 3697 10625 3709 10628
rect 3743 10656 3755 10659
rect 4522 10656 4528 10668
rect 3743 10628 4528 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 4522 10616 4528 10628
rect 4580 10656 4586 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4580 10628 4721 10656
rect 4580 10616 4586 10628
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 6178 10656 6184 10668
rect 5767 10628 6184 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6914 10656 6920 10668
rect 6875 10628 6920 10656
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 8570 10656 8576 10668
rect 7616 10628 8576 10656
rect 7616 10616 7622 10628
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 9490 10656 9496 10668
rect 9451 10628 9496 10656
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 12986 10616 12992 10628
rect 13044 10656 13050 10668
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13044 10628 13461 10656
rect 13044 10616 13050 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 5258 10588 5264 10600
rect 4663 10560 5264 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7742 10588 7748 10600
rect 7340 10560 7748 10588
rect 7340 10548 7346 10560
rect 7742 10548 7748 10560
rect 7800 10588 7806 10600
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 7800 10560 8493 10588
rect 7800 10548 7806 10560
rect 8481 10557 8493 10560
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9766 10588 9772 10600
rect 9723 10560 9772 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 12802 10588 12808 10600
rect 12715 10560 12808 10588
rect 12802 10548 12808 10560
rect 12860 10588 12866 10600
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 12860 10560 14197 10588
rect 12860 10548 12866 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 3973 10523 4031 10529
rect 3973 10520 3985 10523
rect 1627 10492 3985 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 3973 10489 3985 10492
rect 4019 10520 4031 10523
rect 4525 10523 4583 10529
rect 4525 10520 4537 10523
rect 4019 10492 4537 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4525 10489 4537 10492
rect 4571 10489 4583 10523
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 4525 10483 4583 10489
rect 7576 10492 8401 10520
rect 7576 10464 7604 10492
rect 8389 10489 8401 10492
rect 8435 10520 8447 10523
rect 8754 10520 8760 10532
rect 8435 10492 8760 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 8754 10480 8760 10492
rect 8812 10480 8818 10532
rect 9030 10480 9036 10532
rect 9088 10520 9094 10532
rect 9309 10523 9367 10529
rect 9309 10520 9321 10523
rect 9088 10492 9321 10520
rect 9088 10480 9094 10492
rect 9309 10489 9321 10492
rect 9355 10489 9367 10523
rect 9309 10483 9367 10489
rect 9858 10480 9864 10532
rect 9916 10529 9922 10532
rect 9916 10523 9980 10529
rect 9916 10489 9934 10523
rect 9968 10489 9980 10523
rect 12894 10520 12900 10532
rect 12807 10492 12900 10520
rect 9916 10483 9980 10489
rect 9916 10480 9922 10483
rect 12894 10480 12900 10492
rect 12952 10520 12958 10532
rect 13817 10523 13875 10529
rect 13817 10520 13829 10523
rect 12952 10492 13829 10520
rect 12952 10480 12958 10492
rect 13817 10489 13829 10492
rect 13863 10489 13875 10523
rect 13817 10483 13875 10489
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2590 10452 2596 10464
rect 2551 10424 2596 10452
rect 2590 10412 2596 10424
rect 2648 10412 2654 10464
rect 2958 10452 2964 10464
rect 2919 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 3510 10452 3516 10464
rect 3099 10424 3516 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4246 10452 4252 10464
rect 4203 10424 4252 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 6604 10424 6653 10452
rect 6604 10412 6610 10424
rect 6641 10421 6653 10424
rect 6687 10452 6699 10455
rect 7282 10452 7288 10464
rect 6687 10424 7288 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7558 10452 7564 10464
rect 7519 10424 7564 10452
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7800 10424 7849 10452
rect 7800 10412 7806 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8018 10452 8024 10464
rect 7979 10424 8024 10452
rect 7837 10415 7895 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 9214 10452 9220 10464
rect 9175 10424 9220 10452
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 11422 10452 11428 10464
rect 11383 10424 11428 10452
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12710 10452 12716 10464
rect 12483 10424 12716 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12710 10412 12716 10424
rect 12768 10452 12774 10464
rect 13354 10452 13360 10464
rect 12768 10424 13360 10452
rect 12768 10412 12774 10424
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 3016 10220 5089 10248
rect 3016 10208 3022 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 5077 10211 5135 10217
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 3329 10183 3387 10189
rect 3329 10180 3341 10183
rect 2832 10152 3341 10180
rect 2832 10140 2838 10152
rect 3329 10149 3341 10152
rect 3375 10180 3387 10183
rect 4525 10183 4583 10189
rect 3375 10152 4108 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 1664 10115 1722 10121
rect 1664 10081 1676 10115
rect 1710 10112 1722 10115
rect 2498 10112 2504 10124
rect 1710 10084 2504 10112
rect 1710 10081 1722 10084
rect 1664 10075 1722 10081
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 3881 10115 3939 10121
rect 3881 10081 3893 10115
rect 3927 10112 3939 10115
rect 3970 10112 3976 10124
rect 3927 10084 3976 10112
rect 3927 10081 3939 10084
rect 3881 10075 3939 10081
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 4080 9985 4108 10152
rect 4525 10149 4537 10183
rect 4571 10180 4583 10183
rect 4614 10180 4620 10192
rect 4571 10152 4620 10180
rect 4571 10149 4583 10152
rect 4525 10143 4583 10149
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 5092 10180 5120 10211
rect 5258 10208 5264 10260
rect 5316 10248 5322 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 5316 10220 5641 10248
rect 5316 10208 5322 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 5629 10211 5687 10217
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6270 10248 6276 10260
rect 6043 10220 6276 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6270 10208 6276 10220
rect 6328 10248 6334 10260
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 6328 10220 8217 10248
rect 6328 10208 6334 10220
rect 8205 10217 8217 10220
rect 8251 10248 8263 10251
rect 8386 10248 8392 10260
rect 8251 10220 8392 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 8628 10220 9413 10248
rect 8628 10208 8634 10220
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9401 10211 9459 10217
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10686 10248 10692 10260
rect 9723 10220 10692 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 5092 10152 6592 10180
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4212 10084 4445 10112
rect 4212 10072 4218 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 5537 10115 5595 10121
rect 5537 10081 5549 10115
rect 5583 10112 5595 10115
rect 5626 10112 5632 10124
rect 5583 10084 5632 10112
rect 5583 10081 5595 10084
rect 5537 10075 5595 10081
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 6086 10112 6092 10124
rect 5999 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10112 6150 10124
rect 6454 10112 6460 10124
rect 6144 10084 6460 10112
rect 6144 10072 6150 10084
rect 6454 10072 6460 10084
rect 6512 10072 6518 10124
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4396 10016 4629 10044
rect 4396 10004 4402 10016
rect 4617 10013 4629 10016
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6564 10044 6592 10152
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 7340 10152 7880 10180
rect 7340 10140 7346 10152
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7558 10112 7564 10124
rect 6972 10084 7564 10112
rect 6972 10072 6978 10084
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 7653 10047 7711 10053
rect 6564 10016 7236 10044
rect 6273 10007 6331 10013
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9945 4123 9979
rect 6288 9976 6316 10007
rect 6546 9976 6552 9988
rect 6288 9948 6552 9976
rect 4065 9939 4123 9945
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 2777 9911 2835 9917
rect 2777 9908 2789 9911
rect 2096 9880 2789 9908
rect 2096 9868 2102 9880
rect 2777 9877 2789 9880
rect 2823 9877 2835 9911
rect 2777 9871 2835 9877
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7098 9908 7104 9920
rect 6963 9880 7104 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 7208 9917 7236 10016
rect 7653 10013 7665 10047
rect 7699 10044 7711 10047
rect 7742 10044 7748 10056
rect 7699 10016 7748 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 7852 10053 7880 10152
rect 9416 10112 9444 10211
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 13354 10248 13360 10260
rect 13315 10220 13360 10248
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 9858 10140 9864 10192
rect 9916 10180 9922 10192
rect 10045 10183 10103 10189
rect 10045 10180 10057 10183
rect 9916 10152 10057 10180
rect 9916 10140 9922 10152
rect 10045 10149 10057 10152
rect 10091 10180 10103 10183
rect 10134 10180 10140 10192
rect 10091 10152 10140 10180
rect 10091 10149 10103 10152
rect 10045 10143 10103 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 9490 10112 9496 10124
rect 9403 10084 9496 10112
rect 9490 10072 9496 10084
rect 9548 10112 9554 10124
rect 9548 10084 10364 10112
rect 9548 10072 9554 10084
rect 10336 10056 10364 10084
rect 11330 10072 11336 10124
rect 11388 10112 11394 10124
rect 11681 10115 11739 10121
rect 11681 10112 11693 10115
rect 11388 10084 11693 10112
rect 11388 10072 11394 10084
rect 11681 10081 11693 10084
rect 11727 10081 11739 10115
rect 11681 10075 11739 10081
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8202 10044 8208 10056
rect 7883 10016 8208 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10778 10044 10784 10056
rect 10739 10016 10784 10044
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 11238 9976 11244 9988
rect 9824 9948 11244 9976
rect 9824 9936 9830 9948
rect 11238 9936 11244 9948
rect 11296 9976 11302 9988
rect 11440 9976 11468 10007
rect 11296 9948 11468 9976
rect 14093 9979 14151 9985
rect 11296 9936 11302 9948
rect 14093 9945 14105 9979
rect 14139 9976 14151 9979
rect 14550 9976 14556 9988
rect 14139 9948 14556 9976
rect 14139 9945 14151 9948
rect 14093 9939 14151 9945
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 24118 9976 24124 9988
rect 19392 9948 24124 9976
rect 19392 9936 19398 9948
rect 24118 9936 24124 9948
rect 24176 9936 24182 9988
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9877 7251 9911
rect 7193 9871 7251 9877
rect 8941 9911 8999 9917
rect 8941 9877 8953 9911
rect 8987 9908 8999 9911
rect 9030 9908 9036 9920
rect 8987 9880 9036 9908
rect 8987 9877 8999 9880
rect 8941 9871 8999 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 11333 9911 11391 9917
rect 11333 9877 11345 9911
rect 11379 9908 11391 9911
rect 12158 9908 12164 9920
rect 11379 9880 12164 9908
rect 11379 9877 11391 9880
rect 11333 9871 11391 9877
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 12802 9908 12808 9920
rect 12763 9880 12808 9908
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 14274 9868 14280 9920
rect 14332 9908 14338 9920
rect 14369 9911 14427 9917
rect 14369 9908 14381 9911
rect 14332 9880 14381 9908
rect 14332 9868 14338 9880
rect 14369 9877 14381 9880
rect 14415 9877 14427 9911
rect 14369 9871 14427 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2498 9704 2504 9716
rect 1452 9676 2360 9704
rect 2459 9676 2504 9704
rect 1452 9664 1458 9676
rect 1489 9639 1547 9645
rect 1489 9605 1501 9639
rect 1535 9636 1547 9639
rect 2222 9636 2228 9648
rect 1535 9608 2228 9636
rect 1535 9605 1547 9608
rect 1489 9599 1547 9605
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 1670 9528 1676 9580
rect 1728 9568 1734 9580
rect 2038 9568 2044 9580
rect 1728 9540 2044 9568
rect 1728 9528 1734 9540
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2332 9568 2360 9676
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 4522 9704 4528 9716
rect 4483 9676 4528 9704
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 6546 9704 6552 9716
rect 5460 9676 6552 9704
rect 5350 9636 5356 9648
rect 5263 9608 5356 9636
rect 5350 9596 5356 9608
rect 5408 9636 5414 9648
rect 5460 9636 5488 9676
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 9674 9704 9680 9716
rect 9324 9676 9680 9704
rect 5408 9608 5488 9636
rect 5408 9596 5414 9608
rect 8018 9596 8024 9648
rect 8076 9636 8082 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 8076 9608 8217 9636
rect 8076 9596 8082 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 2332 9540 2728 9568
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2590 9500 2596 9512
rect 1995 9472 2596 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 2700 9500 2728 9540
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5684 9540 6009 9568
rect 5684 9528 5690 9540
rect 5997 9537 6009 9540
rect 6043 9568 6055 9571
rect 6270 9568 6276 9580
rect 6043 9540 6276 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 9324 9577 9352 9676
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 12069 9707 12127 9713
rect 12069 9704 12081 9707
rect 11296 9676 12081 9704
rect 11296 9664 11302 9676
rect 12069 9673 12081 9676
rect 12115 9673 12127 9707
rect 12069 9667 12127 9673
rect 12250 9636 12256 9648
rect 12084 9608 12256 9636
rect 12084 9580 12112 9608
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12483 9608 13768 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6788 9540 6837 9568
rect 6788 9528 6794 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 12066 9528 12072 9580
rect 12124 9528 12130 9580
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13538 9568 13544 9580
rect 13127 9540 13544 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2700 9472 3157 9500
rect 3145 9469 3157 9472
rect 3191 9500 3203 9503
rect 4890 9500 4896 9512
rect 3191 9472 4896 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 5000 9472 6561 9500
rect 3053 9435 3111 9441
rect 3053 9401 3065 9435
rect 3099 9432 3111 9435
rect 3412 9435 3470 9441
rect 3412 9432 3424 9435
rect 3099 9404 3424 9432
rect 3099 9401 3111 9404
rect 3053 9395 3111 9401
rect 3412 9401 3424 9404
rect 3458 9432 3470 9435
rect 3602 9432 3608 9444
rect 3458 9404 3608 9432
rect 3458 9401 3470 9404
rect 3412 9395 3470 9401
rect 3602 9392 3608 9404
rect 3660 9392 3666 9444
rect 5000 9432 5028 9472
rect 6549 9469 6561 9472
rect 6595 9500 6607 9503
rect 6914 9500 6920 9512
rect 6595 9472 6920 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7098 9509 7104 9512
rect 7092 9500 7104 9509
rect 7059 9472 7104 9500
rect 7092 9463 7104 9472
rect 7098 9460 7104 9463
rect 7156 9460 7162 9512
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8352 9472 8861 9500
rect 8352 9460 8358 9472
rect 8849 9469 8861 9472
rect 8895 9500 8907 9503
rect 9858 9500 9864 9512
rect 8895 9472 9864 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 12216 9472 12265 9500
rect 12216 9460 12222 9472
rect 12253 9469 12265 9472
rect 12299 9500 12311 9503
rect 12342 9500 12348 9512
rect 12299 9472 12348 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 13740 9500 13768 9608
rect 14550 9568 14556 9580
rect 14511 9540 14556 9568
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14458 9500 14464 9512
rect 13740 9472 14464 9500
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 6086 9432 6092 9444
rect 4540 9404 5028 9432
rect 5644 9404 6092 9432
rect 1854 9364 1860 9376
rect 1815 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 4540 9364 4568 9404
rect 5644 9376 5672 9404
rect 6086 9392 6092 9404
rect 6144 9392 6150 9444
rect 9490 9392 9496 9444
rect 9548 9441 9554 9444
rect 9548 9435 9612 9441
rect 9548 9401 9566 9435
rect 9600 9401 9612 9435
rect 9548 9395 9612 9401
rect 11977 9435 12035 9441
rect 11977 9401 11989 9435
rect 12023 9432 12035 9435
rect 12710 9432 12716 9444
rect 12023 9404 12716 9432
rect 12023 9401 12035 9404
rect 11977 9395 12035 9401
rect 9548 9392 9554 9395
rect 12710 9392 12716 9404
rect 12768 9432 12774 9444
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12768 9404 12909 9432
rect 12768 9392 12774 9404
rect 12897 9401 12909 9404
rect 12943 9401 12955 9435
rect 13906 9432 13912 9444
rect 13819 9404 13912 9432
rect 12897 9395 12955 9401
rect 13906 9392 13912 9404
rect 13964 9432 13970 9444
rect 14369 9435 14427 9441
rect 14369 9432 14381 9435
rect 13964 9404 14381 9432
rect 13964 9392 13970 9404
rect 14369 9401 14381 9404
rect 14415 9401 14427 9435
rect 14369 9395 14427 9401
rect 5626 9364 5632 9376
rect 2280 9336 4568 9364
rect 5587 9336 5632 9364
rect 2280 9324 2286 9336
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 9217 9367 9275 9373
rect 9217 9333 9229 9367
rect 9263 9364 9275 9367
rect 10134 9364 10140 9376
rect 9263 9336 10140 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10686 9364 10692 9376
rect 10647 9336 10692 9364
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11572 9336 11621 9364
rect 11572 9324 11578 9336
rect 11609 9333 11621 9336
rect 11655 9364 11667 9367
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 11655 9336 12817 9364
rect 11655 9333 11667 9336
rect 11609 9327 11667 9333
rect 12805 9333 12817 9336
rect 12851 9333 12863 9367
rect 13538 9364 13544 9376
rect 13499 9336 13544 9364
rect 12805 9327 12863 9333
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 13998 9364 14004 9376
rect 13959 9336 14004 9364
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 2188 9132 2237 9160
rect 2188 9120 2194 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2225 9123 2283 9129
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 2455 9132 3893 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 3881 9129 3893 9132
rect 3927 9160 3939 9163
rect 4062 9160 4068 9172
rect 3927 9132 4068 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4982 9160 4988 9172
rect 4943 9132 4988 9160
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 6549 9163 6607 9169
rect 6549 9160 6561 9163
rect 5092 9132 6561 9160
rect 1762 9052 1768 9104
rect 1820 9092 1826 9104
rect 2777 9095 2835 9101
rect 2777 9092 2789 9095
rect 1820 9064 2789 9092
rect 1820 9052 1826 9064
rect 2777 9061 2789 9064
rect 2823 9061 2835 9095
rect 3050 9092 3056 9104
rect 2963 9064 3056 9092
rect 2777 9055 2835 9061
rect 2976 8965 3004 9064
rect 3050 9052 3056 9064
rect 3108 9092 3114 9104
rect 5092 9092 5120 9132
rect 6549 9129 6561 9132
rect 6595 9129 6607 9163
rect 6549 9123 6607 9129
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 8294 9160 8300 9172
rect 8067 9132 8300 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 9217 9163 9275 9169
rect 9217 9129 9229 9163
rect 9263 9160 9275 9163
rect 9490 9160 9496 9172
rect 9263 9132 9496 9160
rect 9263 9129 9275 9132
rect 9217 9123 9275 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 11330 9160 11336 9172
rect 11291 9132 11336 9160
rect 11330 9120 11336 9132
rect 11388 9160 11394 9172
rect 12802 9160 12808 9172
rect 11388 9132 12808 9160
rect 11388 9120 11394 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13906 9160 13912 9172
rect 13867 9132 13912 9160
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 14458 9160 14464 9172
rect 14419 9132 14464 9160
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 16666 9160 16672 9172
rect 16627 9132 16672 9160
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 5534 9092 5540 9104
rect 3108 9064 5120 9092
rect 5184 9064 5540 9092
rect 3108 9052 3114 9064
rect 4890 8984 4896 9036
rect 4948 9024 4954 9036
rect 5184 9033 5212 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 7926 9092 7932 9104
rect 7852 9064 7932 9092
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 4948 8996 5181 9024
rect 4948 8984 4954 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 5436 9027 5494 9033
rect 5436 8993 5448 9027
rect 5482 9024 5494 9027
rect 6270 9024 6276 9036
rect 5482 8996 6276 9024
rect 5482 8993 5494 8996
rect 5436 8987 5494 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8925 3019 8959
rect 3510 8956 3516 8968
rect 3471 8928 3516 8956
rect 2961 8919 3019 8925
rect 2038 8848 2044 8900
rect 2096 8888 2102 8900
rect 2682 8888 2688 8900
rect 2096 8860 2688 8888
rect 2096 8848 2102 8860
rect 2682 8848 2688 8860
rect 2740 8888 2746 8900
rect 2884 8888 2912 8919
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 7650 8888 7656 8900
rect 2740 8860 2912 8888
rect 3160 8860 5028 8888
rect 7611 8860 7656 8888
rect 2740 8848 2746 8860
rect 1026 8780 1032 8832
rect 1084 8820 1090 8832
rect 3160 8820 3188 8860
rect 1084 8792 3188 8820
rect 1084 8780 1090 8792
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 3510 8820 3516 8832
rect 3292 8792 3516 8820
rect 3292 8780 3298 8792
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4614 8820 4620 8832
rect 4575 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 5000 8820 5028 8860
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 5000 8792 7205 8820
rect 7193 8789 7205 8792
rect 7239 8820 7251 8823
rect 7742 8820 7748 8832
rect 7239 8792 7748 8820
rect 7239 8789 7251 8792
rect 7193 8783 7251 8789
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 7852 8820 7880 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 10965 9095 11023 9101
rect 10965 9061 10977 9095
rect 11011 9092 11023 9095
rect 11670 9095 11728 9101
rect 11670 9092 11682 9095
rect 11011 9064 11682 9092
rect 11011 9061 11023 9064
rect 10965 9055 11023 9061
rect 11670 9061 11682 9064
rect 11716 9092 11728 9095
rect 13538 9092 13544 9104
rect 11716 9064 13544 9092
rect 11716 9061 11728 9064
rect 11670 9055 11728 9061
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 9364 8996 9505 9024
rect 9364 8984 9370 8996
rect 9493 8993 9505 8996
rect 9539 9024 9551 9027
rect 9582 9024 9588 9036
rect 9539 8996 9588 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11425 9027 11483 9033
rect 11425 9024 11437 9027
rect 11296 8996 11437 9024
rect 11296 8984 11302 8996
rect 11425 8993 11437 8996
rect 11471 9024 11483 9027
rect 13446 9024 13452 9036
rect 11471 8996 13452 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 13446 8984 13452 8996
rect 13504 9024 13510 9036
rect 14274 9024 14280 9036
rect 13504 8996 14280 9024
rect 13504 8984 13510 8996
rect 14274 8984 14280 8996
rect 14332 9024 14338 9036
rect 15562 9033 15568 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14332 8996 15301 9024
rect 14332 8984 14338 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15556 9024 15568 9033
rect 15523 8996 15568 9024
rect 15289 8987 15347 8993
rect 15556 8987 15568 8996
rect 15562 8984 15568 8987
rect 15620 8984 15626 9036
rect 7926 8916 7932 8968
rect 7984 8956 7990 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7984 8928 8125 8956
rect 7984 8916 7990 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8386 8956 8392 8968
rect 8260 8928 8392 8956
rect 8260 8916 8266 8928
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9916 8928 10149 8956
rect 9916 8916 9922 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10686 8956 10692 8968
rect 10367 8928 10692 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 9309 8891 9367 8897
rect 9309 8888 9321 8891
rect 8352 8860 9321 8888
rect 8352 8848 8358 8860
rect 9309 8857 9321 8860
rect 9355 8888 9367 8891
rect 9398 8888 9404 8900
rect 9355 8860 9404 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 12802 8888 12808 8900
rect 12715 8860 12808 8888
rect 12802 8848 12808 8860
rect 12860 8888 12866 8900
rect 14550 8888 14556 8900
rect 12860 8860 14556 8888
rect 12860 8848 12866 8860
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 8202 8820 8208 8832
rect 7852 8792 8208 8820
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 8754 8820 8760 8832
rect 8715 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 9766 8820 9772 8832
rect 9723 8792 9772 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 13446 8820 13452 8832
rect 13407 8792 13452 8820
rect 13446 8780 13452 8792
rect 13504 8820 13510 8832
rect 13725 8823 13783 8829
rect 13725 8820 13737 8823
rect 13504 8792 13737 8820
rect 13504 8780 13510 8792
rect 13725 8789 13737 8792
rect 13771 8789 13783 8823
rect 13725 8783 13783 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 3602 8616 3608 8628
rect 3515 8588 3608 8616
rect 3602 8576 3608 8588
rect 3660 8616 3666 8628
rect 5350 8616 5356 8628
rect 3660 8588 5356 8616
rect 3660 8576 3666 8588
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 6270 8616 6276 8628
rect 6183 8588 6276 8616
rect 6270 8576 6276 8588
rect 6328 8616 6334 8628
rect 8018 8616 8024 8628
rect 6328 8588 8024 8616
rect 6328 8576 6334 8588
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8478 8616 8484 8628
rect 8343 8588 8484 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 9674 8616 9680 8628
rect 9587 8588 9680 8616
rect 9674 8576 9680 8588
rect 9732 8616 9738 8628
rect 10042 8616 10048 8628
rect 9732 8588 10048 8616
rect 9732 8576 9738 8588
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 11790 8616 11796 8628
rect 10192 8588 10237 8616
rect 11751 8588 11796 8616
rect 10192 8576 10198 8588
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 4890 8548 4896 8560
rect 4851 8520 4896 8548
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 6822 8548 6828 8560
rect 6783 8520 6828 8548
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 8570 8548 8576 8560
rect 8531 8520 8576 8548
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 11974 8548 11980 8560
rect 10284 8520 11980 8548
rect 10284 8508 10290 8520
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 12621 8551 12679 8557
rect 12621 8517 12633 8551
rect 12667 8548 12679 8551
rect 13814 8548 13820 8560
rect 12667 8520 13820 8548
rect 12667 8517 12679 8520
rect 12621 8511 12679 8517
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 15194 8508 15200 8560
rect 15252 8548 15258 8560
rect 15562 8548 15568 8560
rect 15252 8520 15568 8548
rect 15252 8508 15258 8520
rect 15562 8508 15568 8520
rect 15620 8548 15626 8560
rect 16117 8551 16175 8557
rect 16117 8548 16129 8551
rect 15620 8520 16129 8548
rect 15620 8508 15626 8520
rect 16117 8517 16129 8520
rect 16163 8517 16175 8551
rect 16117 8511 16175 8517
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 2225 8483 2283 8489
rect 2225 8480 2237 8483
rect 1452 8452 2237 8480
rect 1452 8440 1458 8452
rect 2225 8449 2237 8452
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4982 8480 4988 8492
rect 4479 8452 4988 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 2240 8412 2268 8443
rect 4982 8440 4988 8452
rect 5040 8480 5046 8492
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5040 8452 5733 8480
rect 5040 8440 5046 8452
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7064 8452 7389 8480
rect 7064 8440 7070 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 8996 8452 9137 8480
rect 8996 8440 9002 8452
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11146 8480 11152 8492
rect 10827 8452 11152 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 13078 8440 13084 8492
rect 13136 8480 13142 8492
rect 13265 8483 13323 8489
rect 13265 8480 13277 8483
rect 13136 8452 13277 8480
rect 13136 8440 13142 8452
rect 13265 8449 13277 8452
rect 13311 8480 13323 8483
rect 13311 8452 14136 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 2240 8384 2636 8412
rect 2608 8356 2636 8384
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4948 8384 5089 8412
rect 4948 8372 4954 8384
rect 5077 8381 5089 8384
rect 5123 8381 5135 8415
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 5077 8375 5135 8381
rect 6564 8384 7297 8412
rect 6564 8356 6592 8384
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8904 8384 9045 8412
rect 8904 8372 8910 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 9033 8375 9091 8381
rect 10502 8372 10508 8384
rect 10560 8412 10566 8424
rect 10560 8384 10824 8412
rect 10560 8372 10566 8384
rect 10796 8356 10824 8384
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 11848 8384 13001 8412
rect 11848 8372 11854 8384
rect 12989 8381 13001 8384
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 1302 8304 1308 8356
rect 1360 8344 1366 8356
rect 2038 8344 2044 8356
rect 1360 8316 2044 8344
rect 1360 8304 1366 8316
rect 2038 8304 2044 8316
rect 2096 8304 2102 8356
rect 2130 8304 2136 8356
rect 2188 8344 2194 8356
rect 2470 8347 2528 8353
rect 2470 8344 2482 8347
rect 2188 8316 2482 8344
rect 2188 8304 2194 8316
rect 2470 8313 2482 8316
rect 2516 8344 2528 8347
rect 2516 8313 2544 8344
rect 2470 8307 2544 8313
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 1673 8279 1731 8285
rect 1673 8276 1685 8279
rect 1636 8248 1685 8276
rect 1636 8236 1642 8248
rect 1673 8245 1685 8248
rect 1719 8276 1731 8279
rect 1762 8276 1768 8288
rect 1719 8248 1768 8276
rect 1719 8245 1731 8248
rect 1673 8239 1731 8245
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 2516 8276 2544 8307
rect 2590 8304 2596 8356
rect 2648 8304 2654 8356
rect 4801 8347 4859 8353
rect 4801 8313 4813 8347
rect 4847 8344 4859 8347
rect 5258 8344 5264 8356
rect 4847 8316 5264 8344
rect 4847 8313 4859 8316
rect 4801 8307 4859 8313
rect 5258 8304 5264 8316
rect 5316 8344 5322 8356
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5316 8316 5641 8344
rect 5316 8304 5322 8316
rect 5629 8313 5641 8316
rect 5675 8313 5687 8347
rect 6546 8344 6552 8356
rect 6507 8316 6552 8344
rect 5629 8307 5687 8313
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7098 8304 7104 8356
rect 7156 8344 7162 8356
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 7156 8316 7849 8344
rect 7156 8304 7162 8316
rect 7837 8313 7849 8316
rect 7883 8344 7895 8347
rect 7926 8344 7932 8356
rect 7883 8316 7932 8344
rect 7883 8313 7895 8316
rect 7837 8307 7895 8313
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 8812 8316 8953 8344
rect 8812 8304 8818 8316
rect 8941 8313 8953 8316
rect 8987 8344 8999 8347
rect 9582 8344 9588 8356
rect 8987 8316 9588 8344
rect 8987 8313 8999 8316
rect 8941 8307 8999 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 10778 8304 10784 8356
rect 10836 8304 10842 8356
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 14108 8353 14136 8452
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 20254 8412 20260 8424
rect 14240 8384 14285 8412
rect 20215 8384 20260 8412
rect 14240 8372 14246 8384
rect 20254 8372 20260 8384
rect 20312 8412 20318 8424
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20312 8384 21005 8412
rect 20312 8372 20318 8384
rect 20993 8381 21005 8384
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 14458 8353 14464 8356
rect 12161 8347 12219 8353
rect 12161 8344 12173 8347
rect 11388 8316 12173 8344
rect 11388 8304 11394 8316
rect 12161 8313 12173 8316
rect 12207 8344 12219 8347
rect 13081 8347 13139 8353
rect 13081 8344 13093 8347
rect 12207 8316 13093 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 13081 8313 13093 8316
rect 13127 8313 13139 8347
rect 13081 8307 13139 8313
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8344 14151 8347
rect 14452 8344 14464 8353
rect 14139 8316 14464 8344
rect 14139 8313 14151 8316
rect 14093 8307 14151 8313
rect 14452 8307 14464 8316
rect 14458 8304 14464 8307
rect 14516 8304 14522 8356
rect 16666 8344 16672 8356
rect 16627 8316 16672 8344
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 20346 8304 20352 8356
rect 20404 8344 20410 8356
rect 20533 8347 20591 8353
rect 20533 8344 20545 8347
rect 20404 8316 20545 8344
rect 20404 8304 20410 8316
rect 20533 8313 20545 8316
rect 20579 8313 20591 8347
rect 20533 8307 20591 8313
rect 2682 8276 2688 8288
rect 2516 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 5166 8276 5172 8288
rect 5127 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 5537 8279 5595 8285
rect 5537 8276 5549 8279
rect 5500 8248 5549 8276
rect 5500 8236 5506 8248
rect 5537 8245 5549 8248
rect 5583 8245 5595 8279
rect 5537 8239 5595 8245
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7193 8279 7251 8285
rect 7193 8276 7205 8279
rect 6972 8248 7205 8276
rect 6972 8236 6978 8248
rect 7193 8245 7205 8248
rect 7239 8245 7251 8279
rect 7193 8239 7251 8245
rect 8110 8236 8116 8288
rect 8168 8276 8174 8288
rect 9214 8276 9220 8288
rect 8168 8248 9220 8276
rect 8168 8236 8174 8248
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 10042 8276 10048 8288
rect 9955 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8276 10106 8288
rect 10597 8279 10655 8285
rect 10597 8276 10609 8279
rect 10100 8248 10609 8276
rect 10100 8236 10106 8248
rect 10597 8245 10609 8248
rect 10643 8245 10655 8279
rect 10597 8239 10655 8245
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13446 8276 13452 8288
rect 13044 8248 13452 8276
rect 13044 8236 13050 8248
rect 13446 8236 13452 8248
rect 13504 8276 13510 8288
rect 13633 8279 13691 8285
rect 13633 8276 13645 8279
rect 13504 8248 13645 8276
rect 13504 8236 13510 8248
rect 13633 8245 13645 8248
rect 13679 8276 13691 8279
rect 14182 8276 14188 8288
rect 13679 8248 14188 8276
rect 13679 8245 13691 8248
rect 13633 8239 13691 8245
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3421 8075 3479 8081
rect 2832 8044 2877 8072
rect 2832 8032 2838 8044
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 4062 8072 4068 8084
rect 3467 8044 4068 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4798 8072 4804 8084
rect 4571 8044 4804 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 3786 8004 3792 8016
rect 3699 7976 3792 8004
rect 3786 7964 3792 7976
rect 3844 8004 3850 8016
rect 4540 8004 4568 8035
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 8662 8072 8668 8084
rect 7248 8044 8668 8072
rect 7248 8032 7254 8044
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 8849 8075 8907 8081
rect 8849 8041 8861 8075
rect 8895 8072 8907 8075
rect 8938 8072 8944 8084
rect 8895 8044 8944 8072
rect 8895 8041 8907 8044
rect 8849 8035 8907 8041
rect 8938 8032 8944 8044
rect 8996 8072 9002 8084
rect 9490 8072 9496 8084
rect 8996 8044 9496 8072
rect 8996 8032 9002 8044
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 9674 8072 9680 8084
rect 9635 8044 9680 8072
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 10686 8072 10692 8084
rect 10643 8044 10692 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 13078 8072 13084 8084
rect 13039 8044 13084 8072
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13872 8044 14105 8072
rect 13872 8032 13878 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14240 8044 14657 8072
rect 14240 8032 14246 8044
rect 14645 8041 14657 8044
rect 14691 8072 14703 8075
rect 15749 8075 15807 8081
rect 15749 8072 15761 8075
rect 14691 8044 15761 8072
rect 14691 8041 14703 8044
rect 14645 8035 14703 8041
rect 15749 8041 15761 8044
rect 15795 8072 15807 8075
rect 15838 8072 15844 8084
rect 15795 8044 15844 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 18138 8072 18144 8084
rect 18099 8044 18144 8072
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 3844 7976 4568 8004
rect 3844 7964 3850 7976
rect 5350 7964 5356 8016
rect 5408 8004 5414 8016
rect 5997 8007 6055 8013
rect 5997 8004 6009 8007
rect 5408 7976 6009 8004
rect 5408 7964 5414 7976
rect 5997 7973 6009 7976
rect 6043 7973 6055 8007
rect 8294 8004 8300 8016
rect 5997 7967 6055 7973
rect 7668 7976 8300 8004
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 1670 7945 1676 7948
rect 1664 7936 1676 7945
rect 1631 7908 1676 7936
rect 1664 7899 1676 7908
rect 1670 7896 1676 7899
rect 1728 7896 1734 7948
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5905 7939 5963 7945
rect 5905 7936 5917 7939
rect 5224 7908 5917 7936
rect 5224 7896 5230 7908
rect 5905 7905 5917 7908
rect 5951 7905 5963 7939
rect 5905 7899 5963 7905
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 7668 7945 7696 7976
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 9125 8007 9183 8013
rect 9125 8004 9137 8007
rect 8444 7976 9137 8004
rect 8444 7964 8450 7976
rect 9125 7973 9137 7976
rect 9171 7973 9183 8007
rect 9125 7967 9183 7973
rect 10229 8007 10287 8013
rect 10229 7973 10241 8007
rect 10275 8004 10287 8007
rect 10778 8004 10784 8016
rect 10275 7976 10784 8004
rect 10275 7973 10287 7976
rect 10229 7967 10287 7973
rect 10778 7964 10784 7976
rect 10836 7964 10842 8016
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11302 8007 11360 8013
rect 11302 8004 11314 8007
rect 11112 7976 11314 8004
rect 11112 7964 11118 7976
rect 11302 7973 11314 7976
rect 11348 7973 11360 8007
rect 11302 7967 11360 7973
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 7616 7908 7665 7936
rect 7616 7896 7622 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 8110 7936 8116 7948
rect 8071 7908 8116 7936
rect 7653 7899 7711 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 9456 7908 10977 7936
rect 9456 7896 9462 7908
rect 10965 7905 10977 7908
rect 11011 7936 11023 7939
rect 11606 7936 11612 7948
rect 11011 7908 11612 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 14001 7939 14059 7945
rect 14001 7936 14013 7939
rect 13320 7908 14013 7936
rect 13320 7896 13326 7908
rect 14001 7905 14013 7908
rect 14047 7936 14059 7939
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14047 7908 15301 7936
rect 14047 7905 14059 7908
rect 14001 7899 14059 7905
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 16761 7939 16819 7945
rect 16761 7936 16773 7939
rect 15896 7908 16773 7936
rect 15896 7896 15902 7908
rect 16761 7905 16773 7908
rect 16807 7905 16819 7939
rect 16761 7899 16819 7905
rect 17028 7939 17086 7945
rect 17028 7905 17040 7939
rect 17074 7936 17086 7939
rect 17310 7936 17316 7948
rect 17074 7908 17316 7936
rect 17074 7905 17086 7908
rect 17028 7899 17086 7905
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 7248 7840 8217 7868
rect 7248 7828 7254 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 3326 7760 3332 7812
rect 3384 7800 3390 7812
rect 5169 7803 5227 7809
rect 5169 7800 5181 7803
rect 3384 7772 5181 7800
rect 3384 7760 3390 7772
rect 5169 7769 5181 7772
rect 5215 7800 5227 7803
rect 5442 7800 5448 7812
rect 5215 7772 5448 7800
rect 5215 7769 5227 7772
rect 5169 7763 5227 7769
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 7377 7803 7435 7809
rect 7377 7769 7389 7803
rect 7423 7800 7435 7803
rect 7650 7800 7656 7812
rect 7423 7772 7656 7800
rect 7423 7769 7435 7772
rect 7377 7763 7435 7769
rect 7650 7760 7656 7772
rect 7708 7800 7714 7812
rect 8312 7800 8340 7831
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 11057 7871 11115 7877
rect 11057 7868 11069 7871
rect 10008 7840 11069 7868
rect 10008 7828 10014 7840
rect 11057 7837 11069 7840
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 12952 7840 14197 7868
rect 12952 7828 12958 7840
rect 14185 7837 14197 7840
rect 14231 7868 14243 7871
rect 15194 7868 15200 7880
rect 14231 7840 15200 7868
rect 14231 7837 14243 7840
rect 14185 7831 14243 7837
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 12342 7800 12348 7812
rect 7708 7772 8340 7800
rect 12255 7772 12348 7800
rect 7708 7760 7714 7772
rect 4890 7732 4896 7744
rect 4851 7704 4896 7732
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5537 7735 5595 7741
rect 5537 7701 5549 7735
rect 5583 7732 5595 7735
rect 6730 7732 6736 7744
rect 5583 7704 6736 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7466 7732 7472 7744
rect 7427 7704 7472 7732
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 7742 7732 7748 7744
rect 7703 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 12268 7732 12296 7772
rect 12342 7760 12348 7772
rect 12400 7800 12406 7812
rect 14642 7800 14648 7812
rect 12400 7772 14648 7800
rect 12400 7760 12406 7772
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 12434 7732 12440 7744
rect 10827 7704 12296 7732
rect 12395 7704 12440 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13630 7732 13636 7744
rect 13591 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 16485 7735 16543 7741
rect 16485 7701 16497 7735
rect 16531 7732 16543 7735
rect 16942 7732 16948 7744
rect 16531 7704 16948 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4801 7531 4859 7537
rect 4801 7497 4813 7531
rect 4847 7528 4859 7531
rect 5166 7528 5172 7540
rect 4847 7500 5172 7528
rect 4847 7497 4859 7500
rect 4801 7491 4859 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 8168 7500 9321 7528
rect 8168 7488 8174 7500
rect 9309 7497 9321 7500
rect 9355 7497 9367 7531
rect 12894 7528 12900 7540
rect 12855 7500 12900 7528
rect 9309 7491 9367 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13262 7528 13268 7540
rect 13223 7500 13268 7528
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 15838 7528 15844 7540
rect 15799 7500 15844 7528
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 4172 7460 4200 7488
rect 6181 7463 6239 7469
rect 6181 7460 6193 7463
rect 4172 7432 6193 7460
rect 6181 7429 6193 7432
rect 6227 7460 6239 7463
rect 7006 7460 7012 7472
rect 6227 7432 7012 7460
rect 6227 7429 6239 7432
rect 6181 7423 6239 7429
rect 7006 7420 7012 7432
rect 7064 7420 7070 7472
rect 8757 7463 8815 7469
rect 8757 7429 8769 7463
rect 8803 7460 8815 7463
rect 8803 7432 9812 7460
rect 8803 7429 8815 7432
rect 8757 7423 8815 7429
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 5166 7392 5172 7404
rect 5079 7364 5172 7392
rect 5166 7352 5172 7364
rect 5224 7392 5230 7404
rect 5350 7392 5356 7404
rect 5224 7364 5356 7392
rect 5224 7352 5230 7364
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 9784 7401 9812 7432
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 13354 7460 13360 7472
rect 12584 7432 13360 7460
rect 12584 7420 12590 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 9769 7395 9827 7401
rect 6687 7364 7512 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 2590 7284 2596 7336
rect 2648 7324 2654 7336
rect 3050 7333 3056 7336
rect 2777 7327 2835 7333
rect 2777 7324 2789 7327
rect 2648 7296 2789 7324
rect 2648 7284 2654 7296
rect 2777 7293 2789 7296
rect 2823 7293 2835 7327
rect 3044 7324 3056 7333
rect 3011 7296 3056 7324
rect 2777 7287 2835 7293
rect 3044 7287 3056 7296
rect 3050 7284 3056 7287
rect 3108 7284 3114 7336
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6972 7296 7389 7324
rect 6972 7284 6978 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7484 7324 7512 7364
rect 9769 7361 9781 7395
rect 9815 7392 9827 7395
rect 9815 7364 9996 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 7650 7333 7656 7336
rect 7644 7324 7656 7333
rect 7484 7296 7656 7324
rect 7377 7287 7435 7293
rect 7644 7287 7656 7296
rect 2133 7259 2191 7265
rect 2133 7225 2145 7259
rect 2179 7256 2191 7259
rect 2501 7259 2559 7265
rect 2501 7256 2513 7259
rect 2179 7228 2513 7256
rect 2179 7225 2191 7228
rect 2133 7219 2191 7225
rect 2501 7225 2513 7228
rect 2547 7256 2559 7259
rect 3059 7256 3087 7284
rect 2547 7228 3087 7256
rect 7392 7256 7420 7287
rect 7650 7284 7656 7287
rect 7708 7284 7714 7336
rect 9861 7327 9919 7333
rect 9861 7293 9873 7327
rect 9907 7293 9919 7327
rect 9968 7324 9996 7364
rect 12158 7352 12164 7404
rect 12216 7392 12222 7404
rect 12986 7392 12992 7404
rect 12216 7364 12992 7392
rect 12216 7352 12222 7364
rect 12986 7352 12992 7364
rect 13044 7392 13050 7404
rect 16942 7392 16948 7404
rect 13044 7364 13400 7392
rect 16903 7364 16948 7392
rect 13044 7352 13050 7364
rect 10128 7327 10186 7333
rect 10128 7324 10140 7327
rect 9968 7296 10140 7324
rect 9861 7287 9919 7293
rect 10128 7293 10140 7296
rect 10174 7324 10186 7327
rect 10686 7324 10692 7336
rect 10174 7296 10692 7324
rect 10174 7293 10186 7296
rect 10128 7287 10186 7293
rect 8202 7256 8208 7268
rect 7392 7228 8208 7256
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 8202 7216 8208 7228
rect 8260 7216 8266 7268
rect 9876 7256 9904 7287
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 13372 7333 13400 7364
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13613 7327 13671 7333
rect 13613 7324 13625 7327
rect 13504 7296 13625 7324
rect 13504 7284 13510 7296
rect 13613 7293 13625 7296
rect 13659 7293 13671 7327
rect 19702 7324 19708 7336
rect 19663 7296 19708 7324
rect 13613 7287 13671 7293
rect 19702 7284 19708 7296
rect 19760 7324 19766 7336
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 19760 7296 20453 7324
rect 19760 7284 19766 7296
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 9950 7256 9956 7268
rect 9876 7228 9956 7256
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 16206 7256 16212 7268
rect 16167 7228 16212 7256
rect 16206 7216 16212 7228
rect 16264 7256 16270 7268
rect 16853 7259 16911 7265
rect 16853 7256 16865 7259
rect 16264 7228 16865 7256
rect 16264 7216 16270 7228
rect 16853 7225 16865 7228
rect 16899 7225 16911 7259
rect 16853 7219 16911 7225
rect 19981 7259 20039 7265
rect 19981 7225 19993 7259
rect 20027 7256 20039 7259
rect 20714 7256 20720 7268
rect 20027 7228 20720 7256
rect 20027 7225 20039 7228
rect 19981 7219 20039 7225
rect 20714 7216 20720 7228
rect 20772 7216 20778 7268
rect 5261 7191 5319 7197
rect 5261 7157 5273 7191
rect 5307 7188 5319 7191
rect 5442 7188 5448 7200
rect 5307 7160 5448 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 5721 7191 5779 7197
rect 5721 7188 5733 7191
rect 5592 7160 5733 7188
rect 5592 7148 5598 7160
rect 5721 7157 5733 7160
rect 5767 7188 5779 7191
rect 6086 7188 6092 7200
rect 5767 7160 6092 7188
rect 5767 7157 5779 7160
rect 5721 7151 5779 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 11112 7160 11253 7188
rect 11112 7148 11118 7160
rect 11241 7157 11253 7160
rect 11287 7188 11299 7191
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11287 7160 11805 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 11793 7151 11851 7157
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 13998 7188 14004 7200
rect 12299 7160 14004 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 16393 7191 16451 7197
rect 16393 7157 16405 7191
rect 16439 7188 16451 7191
rect 16574 7188 16580 7200
rect 16439 7160 16580 7188
rect 16439 7157 16451 7160
rect 16393 7151 16451 7157
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 16758 7188 16764 7200
rect 16719 7160 16764 7188
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 17310 7148 17316 7200
rect 17368 7188 17374 7200
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 17368 7160 17417 7188
rect 17368 7148 17374 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17405 7151 17463 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1670 6984 1676 6996
rect 1631 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 3786 6984 3792 6996
rect 3747 6956 3792 6984
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 6089 6987 6147 6993
rect 4948 6956 5580 6984
rect 4948 6944 4954 6956
rect 5353 6919 5411 6925
rect 5353 6885 5365 6919
rect 5399 6916 5411 6919
rect 5442 6916 5448 6928
rect 5399 6888 5448 6916
rect 5399 6885 5411 6888
rect 5353 6879 5411 6885
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 2740 6820 2789 6848
rect 2740 6808 2746 6820
rect 2777 6817 2789 6820
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 2869 6851 2927 6857
rect 2869 6817 2881 6851
rect 2915 6848 2927 6851
rect 3050 6848 3056 6860
rect 2915 6820 3056 6848
rect 2915 6817 2927 6820
rect 2869 6811 2927 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 5552 6848 5580 6956
rect 6089 6953 6101 6987
rect 6135 6984 6147 6987
rect 7558 6984 7564 6996
rect 6135 6956 7564 6984
rect 6135 6953 6147 6956
rect 6089 6947 6147 6953
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 7708 6956 8217 6984
rect 7708 6944 7714 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 11606 6984 11612 6996
rect 11567 6956 11612 6984
rect 8205 6947 8263 6953
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 13446 6984 13452 6996
rect 13407 6956 13452 6984
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14001 6987 14059 6993
rect 14001 6984 14013 6987
rect 13872 6956 14013 6984
rect 13872 6944 13878 6956
rect 14001 6953 14013 6956
rect 14047 6953 14059 6987
rect 14001 6947 14059 6953
rect 7466 6916 7472 6928
rect 6840 6888 7472 6916
rect 6638 6848 6644 6860
rect 5552 6820 6644 6848
rect 6638 6808 6644 6820
rect 6696 6848 6702 6860
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 6696 6820 6745 6848
rect 6696 6808 6702 6820
rect 6733 6817 6745 6820
rect 6779 6848 6791 6851
rect 6840 6848 6868 6888
rect 7466 6876 7472 6888
rect 7524 6876 7530 6928
rect 10594 6876 10600 6928
rect 10652 6916 10658 6928
rect 10870 6916 10876 6928
rect 10652 6888 10876 6916
rect 10652 6876 10658 6888
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 11330 6916 11336 6928
rect 10980 6888 11336 6916
rect 6779 6820 6868 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 6914 6808 6920 6860
rect 6972 6808 6978 6860
rect 7092 6851 7150 6857
rect 7092 6817 7104 6851
rect 7138 6848 7150 6851
rect 7374 6848 7380 6860
rect 7138 6820 7380 6848
rect 7138 6817 7150 6820
rect 7092 6811 7150 6817
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 8846 6848 8852 6860
rect 8807 6820 8852 6848
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 9306 6848 9312 6860
rect 9267 6820 9312 6848
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 2958 6780 2964 6792
rect 2919 6752 2964 6780
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5408 6752 5457 6780
rect 5408 6740 5414 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 6825 6783 6883 6789
rect 5592 6752 5637 6780
rect 5592 6740 5598 6752
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 6932 6780 6960 6808
rect 6871 6752 6960 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 2406 6712 2412 6724
rect 2367 6684 2412 6712
rect 2406 6672 2412 6684
rect 2464 6672 2470 6724
rect 4985 6715 5043 6721
rect 4985 6681 4997 6715
rect 5031 6712 5043 6715
rect 6365 6715 6423 6721
rect 6365 6712 6377 6715
rect 5031 6684 6377 6712
rect 5031 6681 5043 6684
rect 4985 6675 5043 6681
rect 6365 6681 6377 6684
rect 6411 6712 6423 6715
rect 6730 6712 6736 6724
rect 6411 6684 6736 6712
rect 6411 6681 6423 6684
rect 6365 6675 6423 6681
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 2038 6644 2044 6656
rect 1999 6616 2044 6644
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 4614 6644 4620 6656
rect 4387 6616 4620 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 5258 6644 5264 6656
rect 4939 6616 5264 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 5258 6604 5264 6616
rect 5316 6644 5322 6656
rect 6549 6647 6607 6653
rect 6549 6644 6561 6647
rect 5316 6616 6561 6644
rect 5316 6604 5322 6616
rect 6549 6613 6561 6616
rect 6595 6644 6607 6647
rect 6840 6644 6868 6743
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10980 6789 11008 6888
rect 11330 6876 11336 6888
rect 11388 6876 11394 6928
rect 12336 6919 12394 6925
rect 12336 6885 12348 6919
rect 12382 6916 12394 6919
rect 12434 6916 12440 6928
rect 12382 6888 12440 6916
rect 12382 6885 12394 6888
rect 12336 6879 12394 6885
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 16758 6916 16764 6928
rect 16592 6888 16764 6916
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 12023 6820 12081 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12069 6817 12081 6820
rect 12115 6848 12127 6851
rect 12158 6848 12164 6860
rect 12115 6820 12164 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14700 6820 14749 6848
rect 14700 6808 14706 6820
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 15378 6848 15384 6860
rect 15339 6820 15384 6848
rect 14737 6811 14795 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6848 16543 6851
rect 16592 6848 16620 6888
rect 16758 6876 16764 6888
rect 16816 6916 16822 6928
rect 17862 6916 17868 6928
rect 16816 6888 17868 6916
rect 16816 6876 16822 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 16531 6820 16620 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17109 6851 17167 6857
rect 17109 6848 17121 6851
rect 17000 6820 17121 6848
rect 17000 6808 17006 6820
rect 17109 6817 17121 6820
rect 17155 6817 17167 6851
rect 17109 6811 17167 6817
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20772 6820 20913 6848
rect 20772 6808 20778 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10468 6752 10977 6780
rect 10468 6740 10474 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 15654 6780 15660 6792
rect 15615 6752 15660 6780
rect 11057 6743 11115 6749
rect 9950 6672 9956 6724
rect 10008 6712 10014 6724
rect 10321 6715 10379 6721
rect 10321 6712 10333 6715
rect 10008 6684 10333 6712
rect 10008 6672 10014 6684
rect 10321 6681 10333 6684
rect 10367 6712 10379 6715
rect 10778 6712 10784 6724
rect 10367 6684 10784 6712
rect 10367 6681 10379 6684
rect 10321 6675 10379 6681
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 11072 6712 11100 6743
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 16850 6780 16856 6792
rect 16811 6752 16856 6780
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 10928 6684 11100 6712
rect 10928 6672 10934 6684
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 14461 6715 14519 6721
rect 14461 6712 14473 6715
rect 14056 6684 14473 6712
rect 14056 6672 14062 6684
rect 14461 6681 14473 6684
rect 14507 6712 14519 6715
rect 14553 6715 14611 6721
rect 14553 6712 14565 6715
rect 14507 6684 14565 6712
rect 14507 6681 14519 6684
rect 14461 6675 14519 6681
rect 14553 6681 14565 6684
rect 14599 6712 14611 6715
rect 16868 6712 16896 6740
rect 14599 6684 16896 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 10502 6644 10508 6656
rect 6595 6616 6868 6644
rect 10463 6616 10508 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 17494 6604 17500 6656
rect 17552 6644 17558 6656
rect 18233 6647 18291 6653
rect 18233 6644 18245 6647
rect 17552 6616 18245 6644
rect 17552 6604 17558 6616
rect 18233 6613 18245 6616
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 21085 6647 21143 6653
rect 21085 6613 21097 6647
rect 21131 6644 21143 6647
rect 21634 6644 21640 6656
rect 21131 6616 21640 6644
rect 21131 6613 21143 6616
rect 21085 6607 21143 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3016 6412 3341 6440
rect 3016 6400 3022 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 5350 6440 5356 6452
rect 5311 6412 5356 6440
rect 3329 6403 3387 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5629 6443 5687 6449
rect 5629 6440 5641 6443
rect 5500 6412 5641 6440
rect 5500 6400 5506 6412
rect 5629 6409 5641 6412
rect 5675 6409 5687 6443
rect 5629 6403 5687 6409
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9548 6412 9781 6440
rect 9548 6400 9554 6412
rect 9769 6409 9781 6412
rect 9815 6409 9827 6443
rect 9769 6403 9827 6409
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10652 6412 10885 6440
rect 10652 6400 10658 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 11480 6412 12081 6440
rect 11480 6400 11486 6412
rect 12069 6409 12081 6412
rect 12115 6440 12127 6443
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 12115 6412 12173 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12492 6412 12537 6440
rect 12492 6400 12498 6412
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15436 6412 16037 6440
rect 15436 6400 15442 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17313 6443 17371 6449
rect 17313 6440 17325 6443
rect 17000 6412 17325 6440
rect 17000 6400 17006 6412
rect 17313 6409 17325 6412
rect 17359 6440 17371 6443
rect 17402 6440 17408 6452
rect 17359 6412 17408 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20772 6412 20913 6440
rect 20772 6400 20778 6412
rect 20901 6409 20913 6412
rect 20947 6409 20959 6443
rect 20901 6403 20959 6409
rect 11885 6375 11943 6381
rect 11885 6341 11897 6375
rect 11931 6372 11943 6375
rect 12342 6372 12348 6384
rect 11931 6344 12348 6372
rect 11931 6341 11943 6344
rect 11885 6335 11943 6341
rect 12342 6332 12348 6344
rect 12400 6372 12406 6384
rect 12400 6344 13032 6372
rect 12400 6332 12406 6344
rect 13004 6316 13032 6344
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 2096 6276 2513 6304
rect 2096 6264 2102 6276
rect 2501 6273 2513 6276
rect 2547 6304 2559 6307
rect 2774 6304 2780 6316
rect 2547 6276 2780 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4338 6304 4344 6316
rect 4203 6276 4344 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 4764 6276 4813 6304
rect 4764 6264 4770 6276
rect 4801 6273 4813 6276
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6319 6276 6653 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 6641 6273 6653 6276
rect 6687 6304 6699 6307
rect 6822 6304 6828 6316
rect 6687 6276 6828 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6822 6264 6828 6276
rect 6880 6304 6886 6316
rect 7374 6304 7380 6316
rect 6880 6276 7380 6304
rect 6880 6264 6886 6276
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 8352 6276 8401 6304
rect 8352 6264 8358 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 12894 6304 12900 6316
rect 12855 6276 12900 6304
rect 8389 6267 8447 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13044 6276 13137 6304
rect 13044 6264 13050 6276
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 14056 6276 14105 6304
rect 14056 6264 14062 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17920 6276 18061 6304
rect 17920 6264 17926 6276
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 1728 6208 2329 6236
rect 1728 6196 1734 6208
rect 2317 6205 2329 6208
rect 2363 6236 2375 6239
rect 3418 6236 3424 6248
rect 2363 6208 3424 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4617 6239 4675 6245
rect 4617 6236 4629 6239
rect 4304 6208 4629 6236
rect 4304 6196 4310 6208
rect 4617 6205 4629 6208
rect 4663 6205 4675 6239
rect 4617 6199 4675 6205
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6788 6208 7205 6236
rect 6788 6196 6794 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6236 12127 6239
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12115 6208 12817 6236
rect 12115 6205 12127 6208
rect 12069 6199 12127 6205
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12912 6236 12940 6264
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 12912 6208 13461 6236
rect 12805 6199 12863 6205
rect 13449 6205 13461 6208
rect 13495 6205 13507 6239
rect 14360 6239 14418 6245
rect 14360 6236 14372 6239
rect 13449 6199 13507 6205
rect 14292 6208 14372 6236
rect 14292 6180 14320 6208
rect 14360 6205 14372 6208
rect 14406 6236 14418 6239
rect 14734 6236 14740 6248
rect 14406 6208 14740 6236
rect 14406 6205 14418 6208
rect 14360 6199 14418 6205
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 16577 6239 16635 6245
rect 16577 6236 16589 6239
rect 16408 6208 16589 6236
rect 3697 6171 3755 6177
rect 3697 6168 3709 6171
rect 2608 6140 3709 6168
rect 2608 6112 2636 6140
rect 3697 6137 3709 6140
rect 3743 6137 3755 6171
rect 5442 6168 5448 6180
rect 3697 6131 3755 6137
rect 4264 6140 5448 6168
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1452 6072 1593 6100
rect 1452 6060 1458 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1581 6063 1639 6069
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2409 6103 2467 6109
rect 2409 6069 2421 6103
rect 2455 6100 2467 6103
rect 2590 6100 2596 6112
rect 2455 6072 2596 6100
rect 2455 6069 2467 6072
rect 2409 6063 2467 6069
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 3050 6100 3056 6112
rect 3011 6072 3056 6100
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 4264 6109 4292 6140
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 6972 6140 7297 6168
rect 6972 6128 6978 6140
rect 7285 6137 7297 6140
rect 7331 6168 7343 6171
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7331 6140 7849 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 7837 6131 7895 6137
rect 8297 6171 8355 6177
rect 8297 6137 8309 6171
rect 8343 6168 8355 6171
rect 8570 6168 8576 6180
rect 8343 6140 8576 6168
rect 8343 6137 8355 6140
rect 8297 6131 8355 6137
rect 8570 6128 8576 6140
rect 8628 6177 8634 6180
rect 8628 6171 8692 6177
rect 8628 6137 8646 6171
rect 8680 6137 8692 6171
rect 8628 6131 8692 6137
rect 8628 6128 8634 6131
rect 10410 6128 10416 6180
rect 10468 6128 10474 6180
rect 11330 6168 11336 6180
rect 11291 6140 11336 6168
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 14001 6171 14059 6177
rect 14001 6137 14013 6171
rect 14047 6168 14059 6171
rect 14274 6168 14280 6180
rect 14047 6140 14280 6168
rect 14047 6137 14059 6140
rect 14001 6131 14059 6137
rect 14274 6128 14280 6140
rect 14332 6128 14338 6180
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4396 6072 4721 6100
rect 4396 6060 4402 6072
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 4709 6063 4767 6069
rect 6825 6103 6883 6109
rect 6825 6069 6837 6103
rect 6871 6100 6883 6103
rect 7558 6100 7564 6112
rect 6871 6072 7564 6100
rect 6871 6069 6883 6072
rect 6825 6063 6883 6069
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10428 6100 10456 6128
rect 16408 6112 16436 6208
rect 16577 6205 16589 6208
rect 16623 6205 16635 6239
rect 16577 6199 16635 6205
rect 16758 6196 16764 6248
rect 16816 6236 16822 6248
rect 19153 6239 19211 6245
rect 19153 6236 19165 6239
rect 16816 6208 19165 6236
rect 16816 6196 16822 6208
rect 19153 6205 19165 6208
rect 19199 6236 19211 6239
rect 19889 6239 19947 6245
rect 19889 6236 19901 6239
rect 19199 6208 19901 6236
rect 19199 6205 19211 6208
rect 19153 6199 19211 6205
rect 19889 6205 19901 6208
rect 19935 6205 19947 6239
rect 19889 6199 19947 6205
rect 16853 6171 16911 6177
rect 16853 6137 16865 6171
rect 16899 6168 16911 6171
rect 17586 6168 17592 6180
rect 16899 6140 17592 6168
rect 16899 6137 16911 6140
rect 16853 6131 16911 6137
rect 17586 6128 17592 6140
rect 17644 6128 17650 6180
rect 19426 6168 19432 6180
rect 19387 6140 19432 6168
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 9916 6072 10517 6100
rect 9916 6060 9922 6072
rect 10505 6069 10517 6072
rect 10551 6069 10563 6103
rect 15470 6100 15476 6112
rect 15431 6072 15476 6100
rect 10505 6063 10563 6069
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 16390 6100 16396 6112
rect 16351 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 17000 6072 17785 6100
rect 17000 6060 17006 6072
rect 17773 6069 17785 6072
rect 17819 6100 17831 6103
rect 18138 6100 18144 6112
rect 17819 6072 18144 6100
rect 17819 6069 17831 6072
rect 17773 6063 17831 6069
rect 18138 6060 18144 6072
rect 18196 6100 18202 6112
rect 18509 6103 18567 6109
rect 18509 6100 18521 6103
rect 18196 6072 18521 6100
rect 18196 6060 18202 6072
rect 18509 6069 18521 6072
rect 18555 6069 18567 6103
rect 18509 6063 18567 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1397 5899 1455 5905
rect 1397 5865 1409 5899
rect 1443 5896 1455 5899
rect 1670 5896 1676 5908
rect 1443 5868 1676 5896
rect 1443 5865 1455 5868
rect 1397 5859 1455 5865
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 1854 5896 1860 5908
rect 1815 5868 1860 5896
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3786 5896 3792 5908
rect 3747 5868 3792 5896
rect 3786 5856 3792 5868
rect 3844 5896 3850 5908
rect 4062 5896 4068 5908
rect 3844 5868 4068 5896
rect 3844 5856 3850 5868
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 6822 5896 6828 5908
rect 6783 5868 6828 5896
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7929 5899 7987 5905
rect 7929 5865 7941 5899
rect 7975 5896 7987 5899
rect 8846 5896 8852 5908
rect 7975 5868 8852 5896
rect 7975 5865 7987 5868
rect 7929 5859 7987 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 9674 5896 9680 5908
rect 9635 5868 9680 5896
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5896 10655 5899
rect 10870 5896 10876 5908
rect 10643 5868 10876 5896
rect 10643 5865 10655 5868
rect 10597 5859 10655 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 12986 5896 12992 5908
rect 12943 5868 12992 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13446 5896 13452 5908
rect 13311 5868 13452 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 13630 5896 13636 5908
rect 13591 5868 13636 5896
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 13998 5896 14004 5908
rect 13780 5868 14004 5896
rect 13780 5856 13786 5868
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14642 5896 14648 5908
rect 14603 5868 14648 5896
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 16574 5896 16580 5908
rect 16535 5868 16580 5896
rect 16574 5856 16580 5868
rect 16632 5896 16638 5908
rect 17129 5899 17187 5905
rect 17129 5896 17141 5899
rect 16632 5868 17141 5896
rect 16632 5856 16638 5868
rect 17129 5865 17141 5868
rect 17175 5865 17187 5899
rect 17129 5859 17187 5865
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 18325 5899 18383 5905
rect 18325 5896 18337 5899
rect 17276 5868 18337 5896
rect 17276 5856 17282 5868
rect 18325 5865 18337 5868
rect 18371 5865 18383 5899
rect 18325 5859 18383 5865
rect 1118 5788 1124 5840
rect 1176 5828 1182 5840
rect 2409 5831 2467 5837
rect 2409 5828 2421 5831
rect 1176 5800 2421 5828
rect 1176 5788 1182 5800
rect 2409 5797 2421 5800
rect 2455 5828 2467 5831
rect 2682 5828 2688 5840
rect 2455 5800 2688 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 2682 5788 2688 5800
rect 2740 5788 2746 5840
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 8754 5828 8760 5840
rect 8444 5800 8760 5828
rect 8444 5788 8450 5800
rect 8754 5788 8760 5800
rect 8812 5828 8818 5840
rect 11146 5837 11152 5840
rect 8941 5831 8999 5837
rect 8941 5828 8953 5831
rect 8812 5800 8953 5828
rect 8812 5788 8818 5800
rect 8941 5797 8953 5800
rect 8987 5828 8999 5831
rect 9309 5831 9367 5837
rect 9309 5828 9321 5831
rect 8987 5800 9321 5828
rect 8987 5797 8999 5800
rect 8941 5791 8999 5797
rect 9309 5797 9321 5800
rect 9355 5797 9367 5831
rect 11140 5828 11152 5837
rect 11107 5800 11152 5828
rect 9309 5791 9367 5797
rect 11140 5791 11152 5800
rect 11146 5788 11152 5791
rect 11204 5788 11210 5840
rect 18785 5831 18843 5837
rect 18785 5797 18797 5831
rect 18831 5828 18843 5831
rect 18874 5828 18880 5840
rect 18831 5800 18880 5828
rect 18831 5797 18843 5800
rect 18785 5791 18843 5797
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1765 5763 1823 5769
rect 1765 5760 1777 5763
rect 1452 5732 1777 5760
rect 1452 5720 1458 5732
rect 1765 5729 1777 5732
rect 1811 5729 1823 5763
rect 1765 5723 1823 5729
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5760 4951 5763
rect 5534 5760 5540 5772
rect 4939 5732 5540 5760
rect 4939 5729 4951 5732
rect 4893 5723 4951 5729
rect 5534 5720 5540 5732
rect 5592 5760 5598 5772
rect 5712 5763 5770 5769
rect 5712 5760 5724 5763
rect 5592 5732 5724 5760
rect 5592 5720 5598 5732
rect 5712 5729 5724 5732
rect 5758 5760 5770 5763
rect 6270 5760 6276 5772
rect 5758 5732 6276 5760
rect 5758 5729 5770 5732
rect 5712 5723 5770 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 8294 5760 8300 5772
rect 8255 5732 8300 5760
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 18012 5732 18705 5760
rect 18012 5720 18018 5732
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2056 5556 2084 5655
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5316 5664 5457 5692
rect 5316 5652 5322 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 5445 5655 5503 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8570 5692 8576 5704
rect 8531 5664 8576 5692
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 10778 5692 10784 5704
rect 10275 5664 10784 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 10778 5652 10784 5664
rect 10836 5692 10842 5704
rect 10873 5695 10931 5701
rect 10873 5692 10885 5695
rect 10836 5664 10885 5692
rect 10836 5652 10842 5664
rect 10873 5661 10885 5664
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13872 5664 14105 5692
rect 13872 5652 13878 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14274 5692 14280 5704
rect 14235 5664 14280 5692
rect 14093 5655 14151 5661
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 17310 5692 17316 5704
rect 17271 5664 17316 5692
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 7837 5627 7895 5633
rect 7837 5593 7849 5627
rect 7883 5624 7895 5627
rect 8588 5624 8616 5652
rect 16758 5624 16764 5636
rect 7883 5596 8616 5624
rect 16719 5596 16764 5624
rect 7883 5593 7895 5596
rect 7837 5587 7895 5593
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 17402 5584 17408 5636
rect 17460 5624 17466 5636
rect 18892 5624 18920 5655
rect 19334 5624 19340 5636
rect 17460 5596 19340 5624
rect 17460 5584 17466 5596
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 2004 5528 2881 5556
rect 2004 5516 2010 5528
rect 2869 5525 2881 5528
rect 2915 5556 2927 5559
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 2915 5528 3157 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3145 5525 3157 5528
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 5261 5559 5319 5565
rect 5261 5525 5273 5559
rect 5307 5556 5319 5559
rect 5350 5556 5356 5568
rect 5307 5528 5356 5556
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7469 5559 7527 5565
rect 7469 5525 7481 5559
rect 7515 5556 7527 5559
rect 8202 5556 8208 5568
rect 7515 5528 8208 5556
rect 7515 5525 7527 5528
rect 7469 5519 7527 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 11882 5516 11888 5568
rect 11940 5556 11946 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 11940 5528 12265 5556
rect 11940 5516 11946 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12253 5519 12311 5525
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 18012 5528 18061 5556
rect 18012 5516 18018 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1673 5355 1731 5361
rect 1673 5321 1685 5355
rect 1719 5352 1731 5355
rect 1854 5352 1860 5364
rect 1719 5324 1860 5352
rect 1719 5321 1731 5324
rect 1673 5315 1731 5321
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 2832 5324 3249 5352
rect 2832 5312 2838 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 5166 5352 5172 5364
rect 5127 5324 5172 5352
rect 3237 5315 3295 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 6638 5352 6644 5364
rect 6599 5324 6644 5352
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 7374 5352 7380 5364
rect 7335 5324 7380 5352
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 9490 5352 9496 5364
rect 9447 5324 9496 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10873 5355 10931 5361
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 11146 5352 11152 5364
rect 10919 5324 11152 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 11146 5312 11152 5324
rect 11204 5352 11210 5364
rect 11425 5355 11483 5361
rect 11425 5352 11437 5355
rect 11204 5324 11437 5352
rect 11204 5312 11210 5324
rect 11425 5321 11437 5324
rect 11471 5321 11483 5355
rect 13630 5352 13636 5364
rect 13591 5324 13636 5352
rect 11425 5315 11483 5321
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 14093 5355 14151 5361
rect 14093 5321 14105 5355
rect 14139 5352 14151 5355
rect 14274 5352 14280 5364
rect 14139 5324 14280 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14792 5324 14933 5352
rect 14792 5312 14798 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 16945 5355 17003 5361
rect 16945 5321 16957 5355
rect 16991 5352 17003 5355
rect 17310 5352 17316 5364
rect 16991 5324 17316 5352
rect 16991 5321 17003 5324
rect 16945 5315 17003 5321
rect 2958 5244 2964 5296
rect 3016 5284 3022 5296
rect 3142 5284 3148 5296
rect 3016 5256 3148 5284
rect 3016 5244 3022 5256
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 4982 5216 4988 5228
rect 4755 5188 4988 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 4982 5176 4988 5188
rect 5040 5216 5046 5228
rect 5534 5216 5540 5228
rect 5040 5188 5540 5216
rect 5040 5176 5046 5188
rect 5534 5176 5540 5188
rect 5592 5216 5598 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5592 5188 5733 5216
rect 5592 5176 5598 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6822 5216 6828 5228
rect 6052 5188 6828 5216
rect 6052 5176 6058 5188
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 8938 5216 8944 5228
rect 8619 5188 8944 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 9508 5216 9536 5312
rect 12437 5287 12495 5293
rect 12437 5253 12449 5287
rect 12483 5284 12495 5287
rect 13722 5284 13728 5296
rect 12483 5256 13728 5284
rect 12483 5253 12495 5256
rect 12437 5247 12495 5253
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 9508 5188 9628 5216
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5117 1915 5151
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 1857 5111 1915 5117
rect 5000 5120 5641 5148
rect 1486 5040 1492 5092
rect 1544 5080 1550 5092
rect 1872 5080 1900 5111
rect 1544 5052 1900 5080
rect 1544 5040 1550 5052
rect 1872 5012 1900 5052
rect 1946 5040 1952 5092
rect 2004 5080 2010 5092
rect 2102 5083 2160 5089
rect 2102 5080 2114 5083
rect 2004 5052 2114 5080
rect 2004 5040 2010 5052
rect 2102 5049 2114 5052
rect 2148 5049 2160 5083
rect 2102 5043 2160 5049
rect 5000 5024 5028 5120
rect 5629 5117 5641 5120
rect 5675 5148 5687 5151
rect 6454 5148 6460 5160
rect 5675 5120 6460 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 8386 5148 8392 5160
rect 7760 5120 8392 5148
rect 7760 5089 7788 5120
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5117 9551 5151
rect 9600 5148 9628 5188
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12768 5188 12909 5216
rect 12768 5176 12774 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13446 5216 13452 5228
rect 13127 5188 13452 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 9749 5151 9807 5157
rect 9749 5148 9761 5151
rect 9600 5120 9761 5148
rect 9493 5111 9551 5117
rect 9749 5117 9761 5120
rect 9795 5117 9807 5151
rect 14182 5148 14188 5160
rect 14143 5120 14188 5148
rect 9749 5111 9807 5117
rect 7745 5083 7803 5089
rect 7745 5080 7757 5083
rect 5552 5052 7757 5080
rect 3142 5012 3148 5024
rect 1872 4984 3148 5012
rect 3142 4972 3148 4984
rect 3200 5012 3206 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3200 4984 3801 5012
rect 3200 4972 3206 4984
rect 3789 4981 3801 4984
rect 3835 5012 3847 5015
rect 4249 5015 4307 5021
rect 4249 5012 4261 5015
rect 3835 4984 4261 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 4249 4981 4261 4984
rect 4295 4981 4307 5015
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 4249 4975 4307 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 5552 5021 5580 5052
rect 7745 5049 7757 5052
rect 7791 5049 7803 5083
rect 9508 5080 9536 5111
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 14936 5148 14964 5315
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 17402 5312 17408 5364
rect 17460 5352 17466 5364
rect 17460 5324 17505 5352
rect 17460 5312 17466 5324
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19392 5324 19441 5352
rect 19392 5312 19398 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 14936 5120 15853 5148
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 16132 5148 16160 5179
rect 16577 5151 16635 5157
rect 16577 5148 16589 5151
rect 16132 5120 16589 5148
rect 15841 5111 15899 5117
rect 16577 5117 16589 5120
rect 16623 5148 16635 5151
rect 16850 5148 16856 5160
rect 16623 5120 16856 5148
rect 16623 5117 16635 5120
rect 16577 5111 16635 5117
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 17770 5148 17776 5160
rect 17731 5120 17776 5148
rect 17770 5108 17776 5120
rect 17828 5108 17834 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 18138 5148 18144 5160
rect 18095 5120 18144 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18138 5108 18144 5120
rect 18196 5108 18202 5160
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 19484 5120 20545 5148
rect 19484 5108 19490 5120
rect 20533 5117 20545 5120
rect 20579 5148 20591 5151
rect 21085 5151 21143 5157
rect 21085 5148 21097 5151
rect 20579 5120 21097 5148
rect 20579 5117 20591 5120
rect 20533 5111 20591 5117
rect 21085 5117 21097 5120
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 10778 5080 10784 5092
rect 9508 5052 10784 5080
rect 7745 5043 7803 5049
rect 10778 5040 10784 5052
rect 10836 5040 10842 5092
rect 12253 5083 12311 5089
rect 12253 5049 12265 5083
rect 12299 5080 12311 5083
rect 12342 5080 12348 5092
rect 12299 5052 12348 5080
rect 12299 5049 12311 5052
rect 12253 5043 12311 5049
rect 12342 5040 12348 5052
rect 12400 5080 12406 5092
rect 12710 5080 12716 5092
rect 12400 5052 12716 5080
rect 12400 5040 12406 5052
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 14458 5080 14464 5092
rect 14419 5052 14464 5080
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 15933 5083 15991 5089
rect 15933 5080 15945 5083
rect 15304 5052 15945 5080
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5408 4984 5549 5012
rect 5408 4972 5414 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 5537 4975 5595 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6914 5012 6920 5024
rect 6875 4984 6920 5012
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 7926 5012 7932 5024
rect 7887 4984 7932 5012
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8389 5015 8447 5021
rect 8389 4981 8401 5015
rect 8435 5012 8447 5015
rect 8570 5012 8576 5024
rect 8435 4984 8576 5012
rect 8435 4981 8447 4984
rect 8389 4975 8447 4981
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 8938 5012 8944 5024
rect 8899 4984 8944 5012
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 9640 4984 11805 5012
rect 9640 4972 9646 4984
rect 11793 4981 11805 4984
rect 11839 5012 11851 5015
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 11839 4984 12817 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 12805 4975 12863 4981
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 15304 5021 15332 5052
rect 15933 5049 15945 5052
rect 15979 5049 15991 5083
rect 15933 5043 15991 5049
rect 17954 5040 17960 5092
rect 18012 5080 18018 5092
rect 18294 5083 18352 5089
rect 18294 5080 18306 5083
rect 18012 5052 18306 5080
rect 18012 5040 18018 5052
rect 18294 5049 18306 5052
rect 18340 5049 18352 5083
rect 18294 5043 18352 5049
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 15068 4984 15301 5012
rect 15068 4972 15074 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 5012 15531 5015
rect 17494 5012 17500 5024
rect 15519 4984 17500 5012
rect 15519 4981 15531 4984
rect 15473 4975 15531 4981
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 20717 5015 20775 5021
rect 20717 4981 20729 5015
rect 20763 5012 20775 5015
rect 22094 5012 22100 5024
rect 20763 4984 22100 5012
rect 20763 4981 20775 4984
rect 20717 4975 20775 4981
rect 22094 4972 22100 4984
rect 22152 4972 22158 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 5994 4768 6000 4820
rect 6052 4808 6058 4820
rect 6178 4808 6184 4820
rect 6052 4780 6184 4808
rect 6052 4768 6058 4780
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 6270 4768 6276 4820
rect 6328 4808 6334 4820
rect 6641 4811 6699 4817
rect 6641 4808 6653 4811
rect 6328 4780 6653 4808
rect 6328 4768 6334 4780
rect 6641 4777 6653 4780
rect 6687 4777 6699 4811
rect 6641 4771 6699 4777
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 8570 4808 8576 4820
rect 7607 4780 8576 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 8570 4768 8576 4780
rect 8628 4808 8634 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 8628 4780 9689 4808
rect 8628 4768 8634 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 13722 4808 13728 4820
rect 13683 4780 13728 4808
rect 9677 4771 9735 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 16025 4811 16083 4817
rect 16025 4808 16037 4811
rect 15436 4780 16037 4808
rect 15436 4768 15442 4780
rect 16025 4777 16037 4780
rect 16071 4777 16083 4811
rect 16025 4771 16083 4777
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 17218 4808 17224 4820
rect 16715 4780 17224 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 18138 4768 18144 4820
rect 18196 4808 18202 4820
rect 19061 4811 19119 4817
rect 19061 4808 19073 4811
rect 18196 4780 19073 4808
rect 18196 4768 18202 4780
rect 19061 4777 19073 4780
rect 19107 4777 19119 4811
rect 19061 4771 19119 4777
rect 4338 4700 4344 4752
rect 4396 4740 4402 4752
rect 4396 4712 6684 4740
rect 4396 4700 4402 4712
rect 1486 4672 1492 4684
rect 1447 4644 1492 4672
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 1756 4675 1814 4681
rect 1756 4641 1768 4675
rect 1802 4672 1814 4675
rect 2222 4672 2228 4684
rect 1802 4644 2228 4672
rect 1802 4641 1814 4644
rect 1756 4635 1814 4641
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 5534 4681 5540 4684
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 4212 4644 5273 4672
rect 4212 4632 4218 4644
rect 5261 4641 5273 4644
rect 5307 4641 5319 4675
rect 5528 4672 5540 4681
rect 5495 4644 5540 4672
rect 5261 4635 5319 4641
rect 5528 4635 5540 4644
rect 5534 4632 5540 4635
rect 5592 4632 5598 4684
rect 6656 4672 6684 4712
rect 7742 4700 7748 4752
rect 7800 4740 7806 4752
rect 7837 4743 7895 4749
rect 7837 4740 7849 4743
rect 7800 4712 7849 4740
rect 7800 4700 7806 4712
rect 7837 4709 7849 4712
rect 7883 4740 7895 4743
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 7883 4712 8401 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 8389 4709 8401 4712
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 8754 4700 8760 4752
rect 8812 4740 8818 4752
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 8812 4712 9045 4740
rect 8812 4700 8818 4712
rect 9033 4709 9045 4712
rect 9079 4709 9091 4743
rect 15010 4740 15016 4752
rect 9033 4703 9091 4709
rect 9324 4712 15016 4740
rect 8478 4672 8484 4684
rect 6656 4644 8484 4672
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9324 4672 9352 4712
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 15105 4743 15163 4749
rect 15105 4709 15117 4743
rect 15151 4740 15163 4743
rect 15470 4740 15476 4752
rect 15151 4712 15476 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 15470 4700 15476 4712
rect 15528 4740 15534 4752
rect 18156 4740 18184 4768
rect 15528 4712 18184 4740
rect 15528 4700 15534 4712
rect 9490 4672 9496 4684
rect 8904 4644 9352 4672
rect 9403 4644 9496 4672
rect 8904 4632 8910 4644
rect 9490 4632 9496 4644
rect 9548 4672 9554 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9548 4644 10057 4672
rect 9548 4632 9554 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 10778 4632 10784 4684
rect 10836 4672 10842 4684
rect 11882 4681 11888 4684
rect 10873 4675 10931 4681
rect 10873 4672 10885 4675
rect 10836 4644 10885 4672
rect 10836 4632 10842 4644
rect 10873 4641 10885 4644
rect 10919 4672 10931 4675
rect 11876 4672 11888 4681
rect 10919 4644 11652 4672
rect 11843 4644 11888 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 11624 4616 11652 4644
rect 11876 4635 11888 4644
rect 11882 4632 11888 4635
rect 11940 4632 11946 4684
rect 14093 4675 14151 4681
rect 14093 4641 14105 4675
rect 14139 4672 14151 4675
rect 14458 4672 14464 4684
rect 14139 4644 14464 4672
rect 14139 4641 14151 4644
rect 14093 4635 14151 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 16776 4681 16804 4712
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 15252 4644 15301 4672
rect 15252 4632 15258 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 16761 4675 16819 4681
rect 16761 4641 16773 4675
rect 16807 4641 16819 4675
rect 16761 4635 16819 4641
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 17017 4675 17075 4681
rect 17017 4672 17029 4675
rect 16908 4644 17029 4672
rect 16908 4632 16914 4644
rect 17017 4641 17029 4644
rect 17063 4641 17075 4675
rect 17017 4635 17075 4641
rect 17586 4632 17592 4684
rect 17644 4672 17650 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 17644 4644 19257 4672
rect 17644 4632 17650 4644
rect 19245 4641 19257 4644
rect 19291 4672 19303 4675
rect 19334 4672 19340 4684
rect 19291 4644 19340 4672
rect 19291 4641 19303 4644
rect 19245 4635 19303 4641
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 21082 4672 21088 4684
rect 20947 4644 21088 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21082 4632 21088 4644
rect 21140 4632 21146 4684
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 8202 4496 8208 4548
rect 8260 4536 8266 4548
rect 8680 4536 8708 4567
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9732 4576 10149 4604
rect 9732 4564 9738 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10962 4604 10968 4616
rect 10367 4576 10968 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 15565 4607 15623 4613
rect 15565 4573 15577 4607
rect 15611 4604 15623 4607
rect 16206 4604 16212 4616
rect 15611 4576 16212 4604
rect 15611 4573 15623 4576
rect 15565 4567 15623 4573
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 9858 4536 9864 4548
rect 8260 4508 9864 4536
rect 8260 4496 8266 4508
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 12986 4536 12992 4548
rect 12947 4508 12992 4536
rect 12986 4496 12992 4508
rect 13044 4496 13050 4548
rect 14182 4536 14188 4548
rect 13096 4508 14188 4536
rect 1854 4428 1860 4480
rect 1912 4468 1918 4480
rect 2869 4471 2927 4477
rect 2869 4468 2881 4471
rect 1912 4440 2881 4468
rect 1912 4428 1918 4440
rect 2869 4437 2881 4440
rect 2915 4437 2927 4471
rect 2869 4431 2927 4437
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 3200 4440 3433 4468
rect 3200 4428 3206 4440
rect 3421 4437 3433 4440
rect 3467 4468 3479 4471
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3467 4440 3801 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3789 4437 3801 4440
rect 3835 4468 3847 4471
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 3835 4440 4261 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4249 4437 4261 4440
rect 4295 4468 4307 4471
rect 4617 4471 4675 4477
rect 4617 4468 4629 4471
rect 4295 4440 4629 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 4617 4437 4629 4440
rect 4663 4468 4675 4471
rect 5077 4471 5135 4477
rect 5077 4468 5089 4471
rect 4663 4440 5089 4468
rect 4663 4437 4675 4440
rect 4617 4431 4675 4437
rect 5077 4437 5089 4440
rect 5123 4468 5135 4471
rect 5258 4468 5264 4480
rect 5123 4440 5264 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 8018 4468 8024 4480
rect 7979 4440 8024 4468
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 13096 4468 13124 4508
rect 14182 4496 14188 4508
rect 14240 4536 14246 4548
rect 14645 4539 14703 4545
rect 14645 4536 14657 4539
rect 14240 4508 14657 4536
rect 14240 4496 14246 4508
rect 14645 4505 14657 4508
rect 14691 4505 14703 4539
rect 14645 4499 14703 4505
rect 14274 4468 14280 4480
rect 8444 4440 13124 4468
rect 14235 4440 14280 4468
rect 8444 4428 8450 4440
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18141 4471 18199 4477
rect 18141 4468 18153 4471
rect 18012 4440 18153 4468
rect 18012 4428 18018 4440
rect 18141 4437 18153 4440
rect 18187 4437 18199 4471
rect 18141 4431 18199 4437
rect 18785 4471 18843 4477
rect 18785 4437 18797 4471
rect 18831 4468 18843 4471
rect 18874 4468 18880 4480
rect 18831 4440 18880 4468
rect 18831 4437 18843 4440
rect 18785 4431 18843 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 19426 4468 19432 4480
rect 19387 4440 19432 4468
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 19886 4468 19892 4480
rect 19847 4440 19892 4468
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 20990 4428 20996 4480
rect 21048 4468 21054 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 21048 4440 21097 4468
rect 21048 4428 21054 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3053 4267 3111 4273
rect 3053 4264 3065 4267
rect 2832 4236 3065 4264
rect 2832 4224 2838 4236
rect 3053 4233 3065 4236
rect 3099 4233 3111 4267
rect 3053 4227 3111 4233
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4128 2286 4140
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2280 4100 2697 4128
rect 2280 4088 2286 4100
rect 2685 4097 2697 4100
rect 2731 4128 2743 4131
rect 2958 4128 2964 4140
rect 2731 4100 2964 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3068 4128 3096 4227
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 8386 4264 8392 4276
rect 7616 4236 8392 4264
rect 7616 4224 7622 4236
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8757 4267 8815 4273
rect 8757 4264 8769 4267
rect 8536 4236 8769 4264
rect 8536 4224 8542 4236
rect 8757 4233 8769 4236
rect 8803 4233 8815 4267
rect 8757 4227 8815 4233
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9548 4236 9781 4264
rect 9548 4224 9554 4236
rect 9769 4233 9781 4236
rect 9815 4233 9827 4267
rect 10870 4264 10876 4276
rect 10831 4236 10876 4264
rect 9769 4227 9827 4233
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 14458 4264 14464 4276
rect 14419 4236 14464 4264
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 5353 4199 5411 4205
rect 5353 4165 5365 4199
rect 5399 4196 5411 4199
rect 5534 4196 5540 4208
rect 5399 4168 5540 4196
rect 5399 4165 5411 4168
rect 5353 4159 5411 4165
rect 5534 4156 5540 4168
rect 5592 4196 5598 4208
rect 9677 4199 9735 4205
rect 5592 4168 6868 4196
rect 5592 4156 5598 4168
rect 3068 4100 3372 4128
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 2314 4060 2320 4072
rect 2179 4032 2320 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 2314 4020 2320 4032
rect 2372 4020 2378 4072
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 3200 4032 3249 4060
rect 3200 4020 3206 4032
rect 3237 4029 3249 4032
rect 3283 4029 3295 4063
rect 3344 4060 3372 4100
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 6840 4128 6868 4168
rect 9677 4165 9689 4199
rect 9723 4196 9735 4199
rect 10042 4196 10048 4208
rect 9723 4168 10048 4196
rect 9723 4165 9735 4168
rect 9677 4159 9735 4165
rect 5316 4100 6776 4128
rect 6840 4100 6960 4128
rect 5316 4088 5322 4100
rect 3493 4063 3551 4069
rect 3493 4060 3505 4063
rect 3344 4032 3505 4060
rect 3237 4023 3295 4029
rect 3493 4029 3505 4032
rect 3539 4029 3551 4063
rect 3493 4023 3551 4029
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 5592 4032 6193 4060
rect 5592 4020 5598 4032
rect 6181 4029 6193 4032
rect 6227 4060 6239 4063
rect 6546 4060 6552 4072
rect 6227 4032 6552 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6748 4060 6776 4100
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6748 4032 6837 4060
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6932 4060 6960 4100
rect 9784 4060 9812 4168
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 9916 4100 10425 4128
rect 9916 4088 9922 4100
rect 10413 4097 10425 4100
rect 10459 4128 10471 4131
rect 10888 4128 10916 4224
rect 15286 4196 15292 4208
rect 15120 4168 15292 4196
rect 10459 4100 10916 4128
rect 12253 4131 12311 4137
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 15013 4131 15071 4137
rect 12299 4100 12572 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 6932 4032 8248 4060
rect 9784 4032 10241 4060
rect 6825 4023 6883 4029
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 6748 3964 7082 3992
rect 6748 3936 6776 3964
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7070 3955 7128 3961
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 2038 3924 2044 3936
rect 1999 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5592 3896 5641 3924
rect 5592 3884 5598 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 6730 3924 6736 3936
rect 6687 3896 6736 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 8220 3933 8248 4032
rect 10229 4029 10241 4032
rect 10275 4060 10287 4063
rect 10686 4060 10692 4072
rect 10275 4032 10692 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12544 4060 12572 4100
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 15120 4128 15148 4168
rect 15286 4156 15292 4168
rect 15344 4156 15350 4208
rect 19426 4196 19432 4208
rect 17880 4168 18644 4196
rect 17880 4140 17908 4168
rect 15470 4128 15476 4140
rect 15059 4100 15148 4128
rect 15431 4100 15476 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17862 4128 17868 4140
rect 17543 4100 17868 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18616 4137 18644 4168
rect 19352 4168 19432 4196
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19352 4128 19380 4168
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 19886 4156 19892 4208
rect 19944 4196 19950 4208
rect 19944 4168 20208 4196
rect 19944 4156 19950 4168
rect 19518 4128 19524 4140
rect 18840 4100 19380 4128
rect 19479 4100 19524 4128
rect 18840 4088 18846 4100
rect 19518 4088 19524 4100
rect 19576 4128 19582 4140
rect 20180 4137 20208 4168
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19576 4100 20085 4128
rect 19576 4088 19582 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 20165 4131 20223 4137
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 12704 4063 12762 4069
rect 12704 4060 12716 4063
rect 12544 4032 12716 4060
rect 12437 4023 12495 4029
rect 12704 4029 12716 4032
rect 12750 4060 12762 4063
rect 12986 4060 12992 4072
rect 12750 4032 12992 4060
rect 12750 4029 12762 4032
rect 12704 4023 12762 4029
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3992 9367 3995
rect 12452 3992 12480 4023
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 17586 4020 17592 4072
rect 17644 4060 17650 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 17644 4032 18521 4060
rect 17644 4020 17650 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 19058 4060 19064 4072
rect 19019 4032 19064 4060
rect 18509 4023 18567 4029
rect 19058 4020 19064 4032
rect 19116 4060 19122 4072
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19116 4032 19993 4060
rect 19116 4020 19122 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 21177 4063 21235 4069
rect 21177 4060 21189 4063
rect 20772 4032 21189 4060
rect 20772 4020 20778 4032
rect 21177 4029 21189 4032
rect 21223 4060 21235 4063
rect 21729 4063 21787 4069
rect 21729 4060 21741 4063
rect 21223 4032 21741 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21729 4029 21741 4032
rect 21775 4029 21787 4063
rect 21729 4023 21787 4029
rect 13262 3992 13268 4004
rect 9355 3964 10180 3992
rect 12452 3964 13268 3992
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 10152 3936 10180 3964
rect 13262 3952 13268 3964
rect 13320 3952 13326 4004
rect 15381 3995 15439 4001
rect 15381 3961 15393 3995
rect 15427 3992 15439 3995
rect 15718 3995 15776 4001
rect 15718 3992 15730 3995
rect 15427 3964 15730 3992
rect 15427 3961 15439 3964
rect 15381 3955 15439 3961
rect 15718 3961 15730 3964
rect 15764 3992 15776 3995
rect 16022 3992 16028 4004
rect 15764 3964 16028 3992
rect 15764 3961 15776 3964
rect 15718 3955 15776 3961
rect 16022 3952 16028 3964
rect 16080 3992 16086 4004
rect 16666 3992 16672 4004
rect 16080 3964 16672 3992
rect 16080 3952 16086 3964
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 17865 3995 17923 4001
rect 17865 3961 17877 3995
rect 17911 3992 17923 3995
rect 18414 3992 18420 4004
rect 17911 3964 18420 3992
rect 17911 3961 17923 3964
rect 17865 3955 17923 3961
rect 18414 3952 18420 3964
rect 18472 3952 18478 4004
rect 20438 3952 20444 4004
rect 20496 3992 20502 4004
rect 22278 3992 22284 4004
rect 20496 3964 21404 3992
rect 22239 3964 22284 3992
rect 20496 3952 20502 3964
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3893 8263 3927
rect 10134 3924 10140 3936
rect 10095 3896 10140 3924
rect 8205 3887 8263 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 11112 3896 11161 3924
rect 11112 3884 11118 3896
rect 11149 3893 11161 3896
rect 11195 3893 11207 3927
rect 11330 3924 11336 3936
rect 11291 3896 11336 3924
rect 11149 3887 11207 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13596 3896 13829 3924
rect 13596 3884 13602 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 13817 3887 13875 3893
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19576 3896 19625 3924
rect 19576 3884 19582 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 20993 3927 21051 3933
rect 20993 3893 21005 3927
rect 21039 3924 21051 3927
rect 21082 3924 21088 3936
rect 21039 3896 21088 3924
rect 21039 3893 21051 3896
rect 20993 3887 21051 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 21376 3933 21404 3964
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3893 21419 3927
rect 21361 3887 21419 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 2777 3723 2835 3729
rect 2777 3720 2789 3723
rect 2464 3692 2789 3720
rect 2464 3680 2470 3692
rect 2777 3689 2789 3692
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 7837 3723 7895 3729
rect 7837 3689 7849 3723
rect 7883 3720 7895 3723
rect 8202 3720 8208 3732
rect 7883 3692 8208 3720
rect 7883 3689 7895 3692
rect 7837 3683 7895 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8812 3692 8953 3720
rect 8812 3680 8818 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9582 3720 9588 3732
rect 9539 3692 9588 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 12158 3720 12164 3732
rect 12119 3692 12164 3720
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 16666 3720 16672 3732
rect 16627 3692 16672 3720
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 16850 3680 16856 3732
rect 16908 3720 16914 3732
rect 17221 3723 17279 3729
rect 17221 3720 17233 3723
rect 16908 3692 17233 3720
rect 16908 3680 16914 3692
rect 17221 3689 17233 3692
rect 17267 3689 17279 3723
rect 17221 3683 17279 3689
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 17460 3692 18460 3720
rect 17460 3680 17466 3692
rect 1765 3655 1823 3661
rect 1765 3621 1777 3655
rect 1811 3652 1823 3655
rect 2314 3652 2320 3664
rect 1811 3624 2320 3652
rect 1811 3621 1823 3624
rect 1765 3615 1823 3621
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 2682 3652 2688 3664
rect 2643 3624 2688 3652
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 8386 3652 8392 3664
rect 8347 3624 8392 3652
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 9858 3612 9864 3664
rect 9916 3661 9922 3664
rect 9916 3655 9980 3661
rect 9916 3621 9934 3655
rect 9968 3621 9980 3655
rect 9916 3615 9980 3621
rect 9916 3612 9922 3615
rect 17494 3612 17500 3664
rect 17552 3652 17558 3664
rect 17589 3655 17647 3661
rect 17589 3652 17601 3655
rect 17552 3624 17601 3652
rect 17552 3612 17558 3624
rect 17589 3621 17601 3624
rect 17635 3621 17647 3655
rect 17589 3615 17647 3621
rect 2038 3544 2044 3596
rect 2096 3584 2102 3596
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 2096 3556 2145 3584
rect 2096 3544 2102 3556
rect 2133 3553 2145 3556
rect 2179 3584 2191 3587
rect 3418 3584 3424 3596
rect 2179 3556 3424 3584
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5316 3556 5457 3584
rect 5316 3544 5322 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5712 3587 5770 3593
rect 5712 3553 5724 3587
rect 5758 3584 5770 3587
rect 6270 3584 6276 3596
rect 5758 3556 6276 3584
rect 5758 3553 5770 3556
rect 5712 3547 5770 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 7469 3587 7527 3593
rect 7469 3553 7481 3587
rect 7515 3584 7527 3587
rect 8297 3587 8355 3593
rect 8297 3584 8309 3587
rect 7515 3556 8309 3584
rect 7515 3553 7527 3556
rect 7469 3547 7527 3553
rect 8297 3553 8309 3556
rect 8343 3584 8355 3587
rect 9677 3587 9735 3593
rect 8343 3556 9076 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 2958 3516 2964 3528
rect 2871 3488 2964 3516
rect 2958 3476 2964 3488
rect 3016 3516 3022 3528
rect 3145 3519 3203 3525
rect 3145 3516 3157 3519
rect 3016 3488 3157 3516
rect 3016 3476 3022 3488
rect 3145 3485 3157 3488
rect 3191 3485 3203 3519
rect 4430 3516 4436 3528
rect 4391 3488 4436 3516
rect 3145 3479 3203 3485
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 2317 3451 2375 3457
rect 2317 3417 2329 3451
rect 2363 3448 2375 3451
rect 2498 3448 2504 3460
rect 2363 3420 2504 3448
rect 2363 3417 2375 3420
rect 2317 3411 2375 3417
rect 2498 3408 2504 3420
rect 2556 3448 2562 3460
rect 3697 3451 3755 3457
rect 3697 3448 3709 3451
rect 2556 3420 3709 3448
rect 2556 3408 2562 3420
rect 3697 3417 3709 3420
rect 3743 3417 3755 3451
rect 3697 3411 3755 3417
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 7929 3451 7987 3457
rect 7929 3448 7941 3451
rect 6512 3420 7941 3448
rect 6512 3408 6518 3420
rect 7929 3417 7941 3420
rect 7975 3417 7987 3451
rect 7929 3411 7987 3417
rect 3145 3383 3203 3389
rect 3145 3349 3157 3383
rect 3191 3380 3203 3383
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3191 3352 3433 3380
rect 3191 3349 3203 3352
rect 3145 3343 3203 3349
rect 3421 3349 3433 3352
rect 3467 3380 3479 3383
rect 3970 3380 3976 3392
rect 3467 3352 3976 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 5261 3383 5319 3389
rect 5261 3349 5273 3383
rect 5307 3380 5319 3383
rect 6472 3380 6500 3408
rect 5307 3352 6500 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 6825 3383 6883 3389
rect 6825 3380 6837 3383
rect 6788 3352 6837 3380
rect 6788 3340 6794 3352
rect 6825 3349 6837 3352
rect 6871 3349 6883 3383
rect 9048 3380 9076 3556
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 11606 3584 11612 3596
rect 9723 3556 11612 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 12526 3584 12532 3596
rect 12487 3556 12532 3584
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 13906 3584 13912 3596
rect 13867 3556 13912 3584
rect 13906 3544 13912 3556
rect 13964 3584 13970 3596
rect 14645 3587 14703 3593
rect 14645 3584 14657 3587
rect 13964 3556 14657 3584
rect 13964 3544 13970 3556
rect 14645 3553 14657 3556
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 15105 3587 15163 3593
rect 15105 3584 15117 3587
rect 14792 3556 15117 3584
rect 14792 3544 14798 3556
rect 15105 3553 15117 3556
rect 15151 3584 15163 3587
rect 15556 3587 15614 3593
rect 15556 3584 15568 3587
rect 15151 3556 15568 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15556 3553 15568 3556
rect 15602 3584 15614 3587
rect 16390 3584 16396 3596
rect 15602 3556 16396 3584
rect 15602 3553 15614 3556
rect 15556 3547 15614 3553
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 11848 3488 12633 3516
rect 11848 3476 11854 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 14090 3516 14096 3528
rect 12768 3488 12813 3516
rect 14051 3488 14096 3516
rect 12768 3476 12774 3488
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 18230 3516 18236 3528
rect 18191 3488 18236 3516
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 18432 3525 18460 3692
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 18877 3723 18935 3729
rect 18877 3720 18889 3723
rect 18564 3692 18889 3720
rect 18564 3680 18570 3692
rect 18877 3689 18889 3692
rect 18923 3720 18935 3723
rect 19518 3720 19524 3732
rect 18923 3692 19524 3720
rect 18923 3689 18935 3692
rect 18877 3683 18935 3689
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 20073 3655 20131 3661
rect 20073 3652 20085 3655
rect 19484 3624 20085 3652
rect 19484 3612 19490 3624
rect 20073 3621 20085 3624
rect 20119 3621 20131 3655
rect 20073 3615 20131 3621
rect 19337 3587 19395 3593
rect 19337 3553 19349 3587
rect 19383 3553 19395 3587
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 19337 3547 19395 3553
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 11606 3408 11612 3460
rect 11664 3448 11670 3460
rect 11701 3451 11759 3457
rect 11701 3448 11713 3451
rect 11664 3420 11713 3448
rect 11664 3408 11670 3420
rect 11701 3417 11713 3420
rect 11747 3448 11759 3451
rect 12069 3451 12127 3457
rect 12069 3448 12081 3451
rect 11747 3420 12081 3448
rect 11747 3417 11759 3420
rect 11701 3411 11759 3417
rect 12069 3417 12081 3420
rect 12115 3448 12127 3451
rect 13262 3448 13268 3460
rect 12115 3420 13268 3448
rect 12115 3417 12127 3420
rect 12069 3411 12127 3417
rect 13262 3408 13268 3420
rect 13320 3448 13326 3460
rect 13633 3451 13691 3457
rect 13633 3448 13645 3451
rect 13320 3420 13645 3448
rect 13320 3408 13326 3420
rect 13633 3417 13645 3420
rect 13679 3448 13691 3451
rect 15304 3448 15332 3476
rect 13679 3420 15332 3448
rect 17773 3451 17831 3457
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 17773 3417 17785 3451
rect 17819 3448 17831 3451
rect 19352 3448 19380 3547
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 22002 3584 22008 3596
rect 21963 3556 22008 3584
rect 22002 3544 22008 3556
rect 22060 3544 22066 3596
rect 24026 3584 24032 3596
rect 23987 3556 24032 3584
rect 24026 3544 24032 3556
rect 24084 3544 24090 3596
rect 19610 3516 19616 3528
rect 19571 3488 19616 3516
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 19426 3448 19432 3460
rect 17819 3420 19432 3448
rect 17819 3417 17831 3420
rect 17773 3411 17831 3417
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 9674 3380 9680 3392
rect 9048 3352 9680 3380
rect 6825 3343 6883 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 11054 3380 11060 3392
rect 11015 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 20772 3352 21097 3380
rect 20772 3340 20778 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 22189 3383 22247 3389
rect 22189 3380 22201 3383
rect 21600 3352 22201 3380
rect 21600 3340 21606 3352
rect 22189 3349 22201 3352
rect 22235 3349 22247 3383
rect 24210 3380 24216 3392
rect 24171 3352 24216 3380
rect 22189 3343 22247 3349
rect 24210 3340 24216 3352
rect 24268 3340 24274 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 3970 3176 3976 3188
rect 3931 3148 3976 3176
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 4488 3148 6561 3176
rect 4488 3136 4494 3148
rect 6549 3145 6561 3148
rect 6595 3176 6607 3179
rect 8021 3179 8079 3185
rect 6595 3148 6960 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 5166 3108 5172 3120
rect 5127 3080 5172 3108
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 6825 3111 6883 3117
rect 6825 3108 6837 3111
rect 5552 3080 6837 3108
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 5552 2984 5580 3080
rect 6825 3077 6837 3080
rect 6871 3077 6883 3111
rect 6825 3071 6883 3077
rect 5718 3040 5724 3052
rect 5679 3012 5724 3040
rect 5718 3000 5724 3012
rect 5776 3040 5782 3052
rect 6730 3040 6736 3052
rect 5776 3012 6736 3040
rect 5776 3000 5782 3012
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 3142 2972 3148 2984
rect 2639 2944 3148 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 3142 2932 3148 2944
rect 3200 2972 3206 2984
rect 4338 2972 4344 2984
rect 3200 2944 4344 2972
rect 3200 2932 3206 2944
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 5534 2972 5540 2984
rect 5495 2944 5540 2972
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 6454 2972 6460 2984
rect 5675 2944 6460 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 6932 2972 6960 3148
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8478 3176 8484 3188
rect 8067 3148 8484 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 8036 3040 8064 3139
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9916 3148 10609 3176
rect 9916 3136 9922 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11238 3176 11244 3188
rect 11195 3148 11244 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12526 3176 12532 3188
rect 12299 3148 12532 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 12710 3176 12716 3188
rect 12671 3148 12716 3176
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 14645 3179 14703 3185
rect 14645 3145 14657 3179
rect 14691 3176 14703 3179
rect 14734 3176 14740 3188
rect 14691 3148 14740 3176
rect 14691 3145 14703 3148
rect 14645 3139 14703 3145
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 15562 3176 15568 3188
rect 15523 3148 15568 3176
rect 15562 3136 15568 3148
rect 15620 3176 15626 3188
rect 17402 3176 17408 3188
rect 15620 3148 16252 3176
rect 17363 3148 17408 3176
rect 15620 3136 15626 3148
rect 9766 3068 9772 3120
rect 9824 3108 9830 3120
rect 10045 3111 10103 3117
rect 10045 3108 10057 3111
rect 9824 3080 10057 3108
rect 9824 3068 9830 3080
rect 10045 3077 10057 3080
rect 10091 3077 10103 3111
rect 11422 3108 11428 3120
rect 11383 3080 11428 3108
rect 10045 3071 10103 3077
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 7515 3012 8064 3040
rect 8573 3043 8631 3049
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8619 3012 8800 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 6932 2944 7205 2972
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 1210 2864 1216 2916
rect 1268 2904 1274 2916
rect 2041 2907 2099 2913
rect 2041 2904 2053 2907
rect 1268 2876 2053 2904
rect 1268 2864 1274 2876
rect 2041 2873 2053 2876
rect 2087 2904 2099 2907
rect 2682 2904 2688 2916
rect 2087 2876 2688 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 2682 2864 2688 2876
rect 2740 2864 2746 2916
rect 2860 2907 2918 2913
rect 2860 2873 2872 2907
rect 2906 2904 2918 2907
rect 3050 2904 3056 2916
rect 2906 2876 3056 2904
rect 2906 2873 2918 2876
rect 2860 2867 2918 2873
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 5718 2904 5724 2916
rect 5123 2876 5724 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 6270 2904 6276 2916
rect 6183 2876 6276 2904
rect 6270 2864 6276 2876
rect 6328 2904 6334 2916
rect 7484 2904 7512 3003
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2941 8723 2975
rect 8772 2972 8800 3012
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 12728 3040 12756 3136
rect 15289 3111 15347 3117
rect 15289 3077 15301 3111
rect 15335 3108 15347 3111
rect 15746 3108 15752 3120
rect 15335 3080 15752 3108
rect 15335 3077 15347 3080
rect 15289 3071 15347 3077
rect 15746 3068 15752 3080
rect 15804 3108 15810 3120
rect 15804 3080 16160 3108
rect 15804 3068 15810 3080
rect 11112 3012 12756 3040
rect 13173 3043 13231 3049
rect 11112 3000 11118 3012
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13219 3012 13400 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 8938 2981 8944 2984
rect 8932 2972 8944 2981
rect 8772 2944 8944 2972
rect 8665 2935 8723 2941
rect 8932 2935 8944 2944
rect 6328 2876 7512 2904
rect 8680 2904 8708 2935
rect 8938 2932 8944 2935
rect 8996 2932 9002 2984
rect 11238 2972 11244 2984
rect 11199 2944 11244 2972
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 13262 2972 13268 2984
rect 13223 2944 13268 2972
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13372 2972 13400 3012
rect 13538 2981 13544 2984
rect 13532 2972 13544 2981
rect 13372 2944 13544 2972
rect 13532 2935 13544 2944
rect 13538 2932 13544 2935
rect 13596 2932 13602 2984
rect 16132 2981 16160 3080
rect 16224 3049 16252 3148
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 17865 3179 17923 3185
rect 17865 3145 17877 3179
rect 17911 3176 17923 3179
rect 18138 3176 18144 3188
rect 17911 3148 18144 3176
rect 17911 3145 17923 3148
rect 17865 3139 17923 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 18380 3148 19441 3176
rect 18380 3136 18386 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 20806 3176 20812 3188
rect 20767 3148 20812 3176
rect 19429 3139 19487 3145
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21637 3179 21695 3185
rect 21637 3176 21649 3179
rect 20956 3148 21649 3176
rect 20956 3136 20962 3148
rect 21637 3145 21649 3148
rect 21683 3145 21695 3179
rect 22002 3176 22008 3188
rect 21963 3148 22008 3176
rect 21637 3139 21695 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23566 3176 23572 3188
rect 23523 3148 23572 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 24213 3179 24271 3185
rect 24213 3176 24225 3179
rect 24084 3148 24225 3176
rect 24084 3136 24090 3148
rect 24213 3145 24225 3148
rect 24259 3145 24271 3179
rect 24213 3139 24271 3145
rect 18049 3111 18107 3117
rect 18049 3077 18061 3111
rect 18095 3108 18107 3111
rect 19334 3108 19340 3120
rect 18095 3080 19340 3108
rect 18095 3077 18107 3080
rect 18049 3071 18107 3077
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 16209 3043 16267 3049
rect 16209 3009 16221 3043
rect 16255 3009 16267 3043
rect 16390 3040 16396 3052
rect 16303 3012 16396 3040
rect 16209 3003 16267 3009
rect 16390 3000 16396 3012
rect 16448 3040 16454 3052
rect 16761 3043 16819 3049
rect 16761 3040 16773 3043
rect 16448 3012 16773 3040
rect 16448 3000 16454 3012
rect 16761 3009 16773 3012
rect 16807 3009 16819 3043
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 16761 3003 16819 3009
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18690 3040 18696 3052
rect 18603 3012 18696 3040
rect 18690 3000 18696 3012
rect 18748 3040 18754 3052
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 18748 3012 19073 3040
rect 18748 3000 18754 3012
rect 19061 3009 19073 3012
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3040 21235 3043
rect 22020 3040 22048 3136
rect 23198 3068 23204 3120
rect 23256 3108 23262 3120
rect 23845 3111 23903 3117
rect 23845 3108 23857 3111
rect 23256 3080 23857 3108
rect 23256 3068 23262 3080
rect 23845 3077 23857 3080
rect 23891 3077 23903 3111
rect 23845 3071 23903 3077
rect 21223 3012 22048 3040
rect 21223 3009 21235 3012
rect 21177 3003 21235 3009
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 18012 2944 18429 2972
rect 18012 2932 18018 2944
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2972 19671 2975
rect 19978 2972 19984 2984
rect 19659 2944 19984 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 19978 2932 19984 2944
rect 20036 2972 20042 2984
rect 20349 2975 20407 2981
rect 20349 2972 20361 2975
rect 20036 2944 20361 2972
rect 20036 2932 20042 2944
rect 20349 2941 20361 2944
rect 20395 2941 20407 2975
rect 20349 2935 20407 2941
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 20864 2944 20913 2972
rect 20864 2932 20870 2944
rect 20901 2941 20913 2944
rect 20947 2941 20959 2975
rect 22186 2972 22192 2984
rect 22147 2944 22192 2972
rect 20901 2935 20959 2941
rect 22186 2932 22192 2944
rect 22244 2972 22250 2984
rect 22741 2975 22799 2981
rect 22741 2972 22753 2975
rect 22244 2944 22753 2972
rect 22244 2932 22250 2944
rect 22741 2941 22753 2944
rect 22787 2941 22799 2975
rect 22741 2935 22799 2941
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23624 2944 23673 2972
rect 23624 2932 23630 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 8754 2904 8760 2916
rect 8680 2876 8760 2904
rect 6328 2864 6334 2876
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 19889 2907 19947 2913
rect 19889 2873 19901 2907
rect 19935 2904 19947 2907
rect 20622 2904 20628 2916
rect 19935 2876 20628 2904
rect 19935 2873 19947 2876
rect 19889 2867 19947 2873
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 256 2808 2329 2836
rect 256 2796 262 2808
rect 2317 2805 2329 2808
rect 2363 2836 2375 2839
rect 2406 2836 2412 2848
rect 2363 2808 2412 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 6288 2836 6316 2864
rect 4755 2808 6316 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 6546 2796 6552 2848
rect 6604 2836 6610 2848
rect 7285 2839 7343 2845
rect 7285 2836 7297 2839
rect 6604 2808 7297 2836
rect 6604 2796 6610 2808
rect 7285 2805 7297 2808
rect 7331 2805 7343 2839
rect 7285 2799 7343 2805
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 9122 2836 9128 2848
rect 8536 2808 9128 2836
rect 8536 2796 8542 2808
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 15746 2836 15752 2848
rect 15707 2808 15752 2836
rect 15746 2796 15752 2808
rect 15804 2796 15810 2848
rect 20162 2796 20168 2848
rect 20220 2836 20226 2848
rect 22373 2839 22431 2845
rect 22373 2836 22385 2839
rect 20220 2808 22385 2836
rect 20220 2796 20226 2808
rect 22373 2805 22385 2808
rect 22419 2805 22431 2839
rect 22373 2799 22431 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2222 2632 2228 2644
rect 1995 2604 2228 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2498 2632 2504 2644
rect 2459 2604 2504 2632
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 6270 2632 6276 2644
rect 5767 2604 6276 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 9214 2632 9220 2644
rect 9175 2604 9220 2632
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 9769 2635 9827 2641
rect 9769 2632 9781 2635
rect 9732 2604 9781 2632
rect 9732 2592 9738 2604
rect 9769 2601 9781 2604
rect 9815 2601 9827 2635
rect 9769 2595 9827 2601
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 10008 2604 10241 2632
rect 10008 2592 10014 2604
rect 10229 2601 10241 2604
rect 10275 2632 10287 2635
rect 10686 2632 10692 2644
rect 10275 2604 10692 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11330 2632 11336 2644
rect 11291 2604 11336 2632
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13722 2632 13728 2644
rect 13683 2604 13728 2632
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 15746 2592 15752 2644
rect 15804 2632 15810 2644
rect 15933 2635 15991 2641
rect 15933 2632 15945 2635
rect 15804 2604 15945 2632
rect 15804 2592 15810 2604
rect 15933 2601 15945 2604
rect 15979 2632 15991 2635
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 15979 2604 16497 2632
rect 15979 2601 15991 2604
rect 15933 2595 15991 2601
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 16485 2595 16543 2601
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 18012 2604 18061 2632
rect 18012 2592 18018 2604
rect 18049 2601 18061 2604
rect 18095 2601 18107 2635
rect 19426 2632 19432 2644
rect 19387 2604 19432 2632
rect 18049 2595 18107 2601
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 24762 2632 24768 2644
rect 24723 2604 24768 2632
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 1670 2524 1676 2576
rect 1728 2564 1734 2576
rect 4614 2573 4620 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 1728 2536 2421 2564
rect 1728 2524 1734 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 2409 2527 2467 2533
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4608 2564 4620 2573
rect 3927 2536 4620 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4608 2527 4620 2536
rect 4614 2524 4620 2527
rect 4672 2524 4678 2576
rect 9232 2564 9260 2592
rect 10134 2564 10140 2576
rect 9232 2536 10140 2564
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 4338 2496 4344 2508
rect 4299 2468 4344 2496
rect 4338 2456 4344 2468
rect 4396 2456 4402 2508
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 6733 2499 6791 2505
rect 6733 2496 6745 2499
rect 6696 2468 6745 2496
rect 6696 2456 6702 2468
rect 6733 2465 6745 2468
rect 6779 2496 6791 2499
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6779 2468 7297 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7285 2465 7297 2468
rect 7331 2496 7343 2499
rect 7558 2496 7564 2508
rect 7331 2468 7564 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 11348 2496 11376 2592
rect 15378 2524 15384 2576
rect 15436 2564 15442 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 15436 2536 16865 2564
rect 15436 2524 15442 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 19889 2567 19947 2573
rect 19889 2533 19901 2567
rect 19935 2564 19947 2567
rect 20530 2564 20536 2576
rect 19935 2536 20536 2564
rect 19935 2533 19947 2536
rect 19889 2527 19947 2533
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 21082 2524 21088 2576
rect 21140 2564 21146 2576
rect 21453 2567 21511 2573
rect 21453 2564 21465 2567
rect 21140 2536 21465 2564
rect 21140 2524 21146 2536
rect 21453 2533 21465 2536
rect 21499 2533 21511 2567
rect 21453 2527 21511 2533
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 8067 2468 10456 2496
rect 11348 2468 11437 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 2682 2428 2688 2440
rect 2595 2400 2688 2428
rect 2682 2388 2688 2400
rect 2740 2428 2746 2440
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 2740 2400 3433 2428
rect 2740 2388 2746 2400
rect 3421 2397 3433 2400
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 7190 2428 7196 2440
rect 6411 2400 7196 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 7190 2388 7196 2400
rect 7248 2428 7254 2440
rect 7374 2428 7380 2440
rect 7248 2400 7380 2428
rect 7248 2388 7254 2400
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 8036 2428 8064 2459
rect 8662 2428 8668 2440
rect 7524 2400 8064 2428
rect 8623 2400 8668 2428
rect 7524 2388 7530 2400
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 10428 2437 10456 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12492 2468 13001 2496
rect 12492 2456 12498 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2496 14151 2499
rect 14182 2496 14188 2508
rect 14139 2468 14188 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 15194 2496 15200 2508
rect 15155 2468 15200 2496
rect 15194 2456 15200 2468
rect 15252 2496 15258 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15252 2468 15853 2496
rect 15252 2456 15258 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 16206 2456 16212 2508
rect 16264 2496 16270 2508
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 16264 2468 17049 2496
rect 16264 2456 16270 2468
rect 17037 2465 17049 2468
rect 17083 2496 17095 2499
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17083 2468 17601 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 18322 2496 18328 2508
rect 18283 2468 18328 2496
rect 17589 2459 17647 2465
rect 18322 2456 18328 2468
rect 18380 2496 18386 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18380 2468 19073 2496
rect 18380 2456 18386 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19613 2499 19671 2505
rect 19613 2496 19625 2499
rect 19392 2468 19625 2496
rect 19392 2456 19398 2468
rect 19613 2465 19625 2468
rect 19659 2496 19671 2499
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 19659 2468 20361 2496
rect 19659 2465 19671 2468
rect 19613 2459 19671 2465
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 20349 2459 20407 2465
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21913 2499 21971 2505
rect 21913 2496 21925 2499
rect 21232 2468 21925 2496
rect 21232 2456 21238 2468
rect 21913 2465 21925 2468
rect 21959 2465 21971 2499
rect 22462 2496 22468 2508
rect 22423 2468 22468 2496
rect 21913 2459 21971 2465
rect 22462 2456 22468 2468
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 10459 2400 10793 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10781 2397 10793 2400
rect 10827 2397 10839 2431
rect 12066 2428 12072 2440
rect 11979 2400 12072 2428
rect 10781 2391 10839 2397
rect 12066 2388 12072 2400
rect 12124 2428 12130 2440
rect 13078 2428 13084 2440
rect 12124 2400 13084 2428
rect 12124 2388 12130 2400
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 13722 2428 13728 2440
rect 13311 2400 13728 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 16022 2428 16028 2440
rect 14967 2400 16028 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 18506 2428 18512 2440
rect 18467 2400 18512 2428
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 2041 2363 2099 2369
rect 2041 2329 2053 2363
rect 2087 2360 2099 2363
rect 2590 2360 2596 2372
rect 2087 2332 2596 2360
rect 2087 2329 2099 2332
rect 2041 2323 2099 2329
rect 2590 2320 2596 2332
rect 2648 2320 2654 2372
rect 6917 2363 6975 2369
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 8297 2363 8355 2369
rect 8297 2360 8309 2363
rect 6963 2332 8309 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 8297 2329 8309 2332
rect 8343 2360 8355 2363
rect 8386 2360 8392 2372
rect 8343 2332 8392 2360
rect 8343 2329 8355 2332
rect 8297 2323 8355 2329
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 15470 2360 15476 2372
rect 12492 2332 12537 2360
rect 15431 2332 15476 2360
rect 12492 2320 12498 2332
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17221 2363 17279 2369
rect 17221 2360 17233 2363
rect 16172 2332 17233 2360
rect 16172 2320 16178 2332
rect 17221 2329 17233 2332
rect 17267 2329 17279 2363
rect 17221 2323 17279 2329
rect 9398 2252 9404 2304
rect 9456 2292 9462 2304
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 9456 2264 9505 2292
rect 9456 2252 9462 2264
rect 9493 2261 9505 2264
rect 9539 2292 9551 2295
rect 9950 2292 9956 2304
rect 9539 2264 9956 2292
rect 9539 2261 9551 2264
rect 9493 2255 9551 2261
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 14369 2295 14427 2301
rect 14369 2261 14381 2295
rect 14415 2292 14427 2295
rect 15378 2292 15384 2304
rect 14415 2264 15384 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 15378 2252 15384 2264
rect 15436 2252 15442 2304
rect 22646 2292 22652 2304
rect 22607 2264 22652 2292
rect 22646 2252 22652 2264
rect 22704 2252 22710 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 11974 1980 11980 2032
rect 12032 2020 12038 2032
rect 14918 2020 14924 2032
rect 12032 1992 14924 2020
rect 12032 1980 12038 1992
rect 14918 1980 14924 1992
rect 14976 1980 14982 2032
rect 23474 1980 23480 2032
rect 23532 2020 23538 2032
rect 24302 2020 24308 2032
rect 23532 1992 24308 2020
rect 23532 1980 23538 1992
rect 24302 1980 24308 1992
rect 24360 1980 24366 2032
rect 6730 552 6736 604
rect 6788 592 6794 604
rect 6822 592 6828 604
rect 6788 564 6828 592
rect 6788 552 6794 564
rect 6822 552 6828 564
rect 6880 552 6886 604
rect 7834 552 7840 604
rect 7892 592 7898 604
rect 8110 592 8116 604
rect 7892 564 8116 592
rect 7892 552 7898 564
rect 8110 552 8116 564
rect 8168 552 8174 604
rect 12158 552 12164 604
rect 12216 592 12222 604
rect 12250 592 12256 604
rect 12216 564 12256 592
rect 12216 552 12222 564
rect 12250 552 12256 564
rect 12308 552 12314 604
rect 13814 552 13820 604
rect 13872 592 13878 604
rect 13906 592 13912 604
rect 13872 564 13912 592
rect 13872 552 13878 564
rect 13906 552 13912 564
rect 13964 552 13970 604
rect 24946 552 24952 604
rect 25004 592 25010 604
rect 25406 592 25412 604
rect 25004 564 25412 592
rect 25004 552 25010 564
rect 25406 552 25412 564
rect 25464 552 25470 604
rect 26234 552 26240 604
rect 26292 592 26298 604
rect 27062 592 27068 604
rect 26292 564 27068 592
rect 26292 552 26298 564
rect 27062 552 27068 564
rect 27120 552 27126 604
<< via1 >>
rect 3240 26324 3292 26376
rect 10048 26324 10100 26376
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 1584 25483 1636 25492
rect 1584 25449 1593 25483
rect 1593 25449 1627 25483
rect 1627 25449 1636 25483
rect 1584 25440 1636 25449
rect 2596 25304 2648 25356
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 1952 24599 2004 24608
rect 1952 24565 1961 24599
rect 1961 24565 1995 24599
rect 1995 24565 2004 24599
rect 1952 24556 2004 24565
rect 2596 24556 2648 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 2688 24395 2740 24404
rect 2688 24361 2697 24395
rect 2697 24361 2731 24395
rect 2731 24361 2740 24395
rect 2688 24352 2740 24361
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 2504 24259 2556 24268
rect 2504 24225 2513 24259
rect 2513 24225 2547 24259
rect 2547 24225 2556 24259
rect 2504 24216 2556 24225
rect 1676 24012 1728 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1400 23808 1452 23860
rect 1860 23808 1912 23860
rect 2504 23808 2556 23860
rect 3148 23851 3200 23860
rect 3148 23817 3157 23851
rect 3157 23817 3191 23851
rect 3191 23817 3200 23851
rect 3148 23808 3200 23817
rect 7012 23851 7064 23860
rect 7012 23817 7021 23851
rect 7021 23817 7055 23851
rect 7055 23817 7064 23851
rect 7012 23808 7064 23817
rect 20996 23808 21048 23860
rect 1676 23647 1728 23656
rect 1676 23613 1685 23647
rect 1685 23613 1719 23647
rect 1719 23613 1728 23647
rect 1676 23604 1728 23613
rect 7472 23579 7524 23588
rect 7472 23545 7481 23579
rect 7481 23545 7515 23579
rect 7515 23545 7524 23579
rect 7472 23536 7524 23545
rect 3608 23511 3660 23520
rect 3608 23477 3617 23511
rect 3617 23477 3651 23511
rect 3651 23477 3660 23511
rect 3608 23468 3660 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 4160 23264 4212 23316
rect 1952 23239 2004 23248
rect 1952 23205 1961 23239
rect 1961 23205 1995 23239
rect 1995 23205 2004 23239
rect 1952 23196 2004 23205
rect 2780 23128 2832 23180
rect 3976 23128 4028 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 3056 22763 3108 22772
rect 3056 22729 3065 22763
rect 3065 22729 3099 22763
rect 3099 22729 3108 22763
rect 3056 22720 3108 22729
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 3148 22516 3200 22568
rect 2412 22491 2464 22500
rect 2412 22457 2421 22491
rect 2421 22457 2455 22491
rect 2455 22457 2464 22491
rect 2412 22448 2464 22457
rect 2780 22423 2832 22432
rect 2780 22389 2789 22423
rect 2789 22389 2823 22423
rect 2823 22389 2832 22423
rect 2780 22380 2832 22389
rect 3976 22380 4028 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 3976 22108 4028 22160
rect 8024 22040 8076 22092
rect 2964 21972 3016 22024
rect 3976 21972 4028 22024
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 4252 21947 4304 21956
rect 4252 21913 4261 21947
rect 4261 21913 4295 21947
rect 4295 21913 4304 21947
rect 4252 21904 4304 21913
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 4436 21675 4488 21684
rect 4436 21641 4445 21675
rect 4445 21641 4479 21675
rect 4479 21641 4488 21675
rect 4436 21632 4488 21641
rect 3148 21539 3200 21548
rect 3148 21505 3157 21539
rect 3157 21505 3191 21539
rect 3191 21505 3200 21539
rect 3148 21496 3200 21505
rect 1952 21403 2004 21412
rect 1952 21369 1961 21403
rect 1961 21369 1995 21403
rect 1995 21369 2004 21403
rect 1952 21360 2004 21369
rect 4252 21471 4304 21480
rect 4252 21437 4261 21471
rect 4261 21437 4295 21471
rect 4295 21437 4304 21471
rect 4252 21428 4304 21437
rect 2504 21335 2556 21344
rect 2504 21301 2513 21335
rect 2513 21301 2547 21335
rect 2547 21301 2556 21335
rect 2504 21292 2556 21301
rect 2964 21292 3016 21344
rect 3792 21335 3844 21344
rect 3792 21301 3801 21335
rect 3801 21301 3835 21335
rect 3835 21301 3844 21335
rect 3792 21292 3844 21301
rect 3976 21292 4028 21344
rect 8024 21335 8076 21344
rect 8024 21301 8033 21335
rect 8033 21301 8067 21335
rect 8067 21301 8076 21335
rect 8024 21292 8076 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 3516 21088 3568 21140
rect 9680 21131 9732 21140
rect 9680 21097 9689 21131
rect 9689 21097 9723 21131
rect 9723 21097 9732 21131
rect 9680 21088 9732 21097
rect 11336 21131 11388 21140
rect 11336 21097 11345 21131
rect 11345 21097 11379 21131
rect 11379 21097 11388 21131
rect 11336 21088 11388 21097
rect 3976 21020 4028 21072
rect 6276 21063 6328 21072
rect 6276 21029 6285 21063
rect 6285 21029 6319 21063
rect 6319 21029 6328 21063
rect 6276 21020 6328 21029
rect 12348 21020 12400 21072
rect 2320 20952 2372 21004
rect 2872 20995 2924 21004
rect 2872 20961 2881 20995
rect 2881 20961 2915 20995
rect 2915 20961 2924 20995
rect 2872 20952 2924 20961
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 4068 20952 4120 20961
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 9680 20952 9732 21004
rect 11980 20952 12032 21004
rect 10140 20927 10192 20936
rect 10140 20893 10149 20927
rect 10149 20893 10183 20927
rect 10183 20893 10192 20927
rect 10140 20884 10192 20893
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 11520 20816 11572 20868
rect 3056 20791 3108 20800
rect 3056 20757 3065 20791
rect 3065 20757 3099 20791
rect 3099 20757 3108 20791
rect 3056 20748 3108 20757
rect 7564 20748 7616 20800
rect 12440 20791 12492 20800
rect 12440 20757 12449 20791
rect 12449 20757 12483 20791
rect 12483 20757 12492 20791
rect 12440 20748 12492 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 4252 20587 4304 20596
rect 4252 20553 4261 20587
rect 4261 20553 4295 20587
rect 4295 20553 4304 20587
rect 4252 20544 4304 20553
rect 9680 20544 9732 20596
rect 11980 20544 12032 20596
rect 6000 20476 6052 20528
rect 2872 20408 2924 20460
rect 7564 20451 7616 20460
rect 7564 20417 7573 20451
rect 7573 20417 7607 20451
rect 7607 20417 7616 20451
rect 7564 20408 7616 20417
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 9496 20383 9548 20392
rect 2412 20204 2464 20256
rect 9496 20349 9505 20383
rect 9505 20349 9539 20383
rect 9539 20349 9548 20383
rect 9496 20340 9548 20349
rect 6920 20272 6972 20324
rect 10232 20340 10284 20392
rect 11520 20383 11572 20392
rect 11520 20349 11529 20383
rect 11529 20349 11563 20383
rect 11563 20349 11572 20383
rect 11520 20340 11572 20349
rect 9772 20315 9824 20324
rect 9772 20281 9806 20315
rect 9806 20281 9824 20315
rect 9772 20272 9824 20281
rect 3332 20204 3384 20256
rect 4068 20204 4120 20256
rect 6184 20204 6236 20256
rect 7472 20247 7524 20256
rect 7472 20213 7481 20247
rect 7481 20213 7515 20247
rect 7515 20213 7524 20247
rect 7472 20204 7524 20213
rect 12164 20272 12216 20324
rect 10692 20204 10744 20256
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 5540 20043 5592 20052
rect 5540 20009 5549 20043
rect 5549 20009 5583 20043
rect 5583 20009 5592 20043
rect 5540 20000 5592 20009
rect 6000 20043 6052 20052
rect 6000 20009 6009 20043
rect 6009 20009 6043 20043
rect 6043 20009 6052 20043
rect 6000 20000 6052 20009
rect 7564 20000 7616 20052
rect 8116 20000 8168 20052
rect 9680 20043 9732 20052
rect 9680 20009 9689 20043
rect 9689 20009 9723 20043
rect 9723 20009 9732 20043
rect 9680 20000 9732 20009
rect 10140 20043 10192 20052
rect 10140 20009 10149 20043
rect 10149 20009 10183 20043
rect 10183 20009 10192 20043
rect 10140 20000 10192 20009
rect 10692 20043 10744 20052
rect 10692 20009 10701 20043
rect 10701 20009 10735 20043
rect 10735 20009 10744 20043
rect 10692 20000 10744 20009
rect 12164 20043 12216 20052
rect 12164 20009 12173 20043
rect 12173 20009 12207 20043
rect 12207 20009 12216 20043
rect 12164 20000 12216 20009
rect 1492 19907 1544 19916
rect 1492 19873 1501 19907
rect 1501 19873 1535 19907
rect 1535 19873 1544 19907
rect 1492 19864 1544 19873
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 4068 19907 4120 19916
rect 2780 19864 2832 19873
rect 4068 19873 4077 19907
rect 4077 19873 4111 19907
rect 4111 19873 4120 19907
rect 4068 19864 4120 19873
rect 5448 19864 5500 19916
rect 7380 19907 7432 19916
rect 7380 19873 7414 19907
rect 7414 19873 7432 19907
rect 7380 19864 7432 19873
rect 7104 19839 7156 19848
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 7104 19796 7156 19805
rect 10692 19796 10744 19848
rect 2320 19703 2372 19712
rect 2320 19669 2329 19703
rect 2329 19669 2363 19703
rect 2363 19669 2372 19703
rect 2320 19660 2372 19669
rect 2964 19703 3016 19712
rect 2964 19669 2973 19703
rect 2973 19669 3007 19703
rect 3007 19669 3016 19703
rect 2964 19660 3016 19669
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 4896 19703 4948 19712
rect 4896 19669 4905 19703
rect 4905 19669 4939 19703
rect 4939 19669 4948 19703
rect 4896 19660 4948 19669
rect 8300 19660 8352 19712
rect 9496 19660 9548 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 3332 19499 3384 19508
rect 2780 19456 2832 19465
rect 3332 19465 3341 19499
rect 3341 19465 3375 19499
rect 3375 19465 3384 19499
rect 3332 19456 3384 19465
rect 8116 19499 8168 19508
rect 8116 19465 8125 19499
rect 8125 19465 8159 19499
rect 8159 19465 8168 19499
rect 8116 19456 8168 19465
rect 10140 19456 10192 19508
rect 12348 19456 12400 19508
rect 12532 19456 12584 19508
rect 3424 19320 3476 19372
rect 3792 19363 3844 19372
rect 3792 19329 3801 19363
rect 3801 19329 3835 19363
rect 3835 19329 3844 19363
rect 3792 19320 3844 19329
rect 3976 19363 4028 19372
rect 3976 19329 3985 19363
rect 3985 19329 4019 19363
rect 4019 19329 4028 19363
rect 3976 19320 4028 19329
rect 6920 19320 6972 19372
rect 4804 19252 4856 19304
rect 5540 19252 5592 19304
rect 8300 19295 8352 19304
rect 8300 19261 8309 19295
rect 8309 19261 8343 19295
rect 8343 19261 8352 19295
rect 8300 19252 8352 19261
rect 9772 19320 9824 19372
rect 12164 19320 12216 19372
rect 12624 19320 12676 19372
rect 2780 19184 2832 19236
rect 4160 19184 4212 19236
rect 2504 19116 2556 19168
rect 2596 19116 2648 19168
rect 4068 19116 4120 19168
rect 4436 19159 4488 19168
rect 4436 19125 4445 19159
rect 4445 19125 4479 19159
rect 4479 19125 4488 19159
rect 4436 19116 4488 19125
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 4896 19116 4948 19168
rect 6736 19116 6788 19168
rect 7104 19116 7156 19168
rect 7380 19116 7432 19168
rect 8668 19116 8720 19168
rect 9128 19116 9180 19168
rect 11336 19116 11388 19168
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 14372 19116 14424 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1492 18912 1544 18964
rect 2228 18955 2280 18964
rect 2228 18921 2237 18955
rect 2237 18921 2271 18955
rect 2271 18921 2280 18955
rect 2228 18912 2280 18921
rect 2964 18955 3016 18964
rect 2964 18921 2973 18955
rect 2973 18921 3007 18955
rect 3007 18921 3016 18955
rect 2964 18912 3016 18921
rect 7196 18955 7248 18964
rect 7196 18921 7205 18955
rect 7205 18921 7239 18955
rect 7239 18921 7248 18955
rect 7196 18912 7248 18921
rect 9772 18912 9824 18964
rect 12624 18955 12676 18964
rect 12624 18921 12633 18955
rect 12633 18921 12667 18955
rect 12667 18921 12676 18955
rect 12624 18912 12676 18921
rect 3976 18844 4028 18896
rect 5172 18844 5224 18896
rect 6920 18844 6972 18896
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 2780 18776 2832 18785
rect 3240 18776 3292 18828
rect 3884 18776 3936 18828
rect 4712 18819 4764 18828
rect 4712 18785 4721 18819
rect 4721 18785 4755 18819
rect 4755 18785 4764 18819
rect 4712 18776 4764 18785
rect 6184 18776 6236 18828
rect 10968 18819 11020 18828
rect 10968 18785 11002 18819
rect 11002 18785 11020 18819
rect 10968 18776 11020 18785
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 7748 18751 7800 18760
rect 7748 18717 7757 18751
rect 7757 18717 7791 18751
rect 7791 18717 7800 18751
rect 7748 18708 7800 18717
rect 10692 18751 10744 18760
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 2688 18615 2740 18624
rect 2688 18581 2697 18615
rect 2697 18581 2731 18615
rect 2731 18581 2740 18615
rect 2688 18572 2740 18581
rect 6092 18615 6144 18624
rect 6092 18581 6101 18615
rect 6101 18581 6135 18615
rect 6135 18581 6144 18615
rect 6092 18572 6144 18581
rect 6736 18615 6788 18624
rect 6736 18581 6745 18615
rect 6745 18581 6779 18615
rect 6779 18581 6788 18615
rect 6736 18572 6788 18581
rect 6920 18572 6972 18624
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 9680 18572 9732 18624
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2872 18411 2924 18420
rect 2872 18377 2881 18411
rect 2881 18377 2915 18411
rect 2915 18377 2924 18411
rect 2872 18368 2924 18377
rect 3240 18411 3292 18420
rect 3240 18377 3249 18411
rect 3249 18377 3283 18411
rect 3283 18377 3292 18411
rect 3240 18368 3292 18377
rect 6184 18368 6236 18420
rect 7472 18368 7524 18420
rect 8668 18411 8720 18420
rect 8668 18377 8677 18411
rect 8677 18377 8711 18411
rect 8711 18377 8720 18411
rect 8668 18368 8720 18377
rect 9220 18411 9272 18420
rect 9220 18377 9229 18411
rect 9229 18377 9263 18411
rect 9263 18377 9272 18411
rect 9220 18368 9272 18377
rect 12440 18368 12492 18420
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 1768 18164 1820 18216
rect 2780 18164 2832 18216
rect 3884 18164 3936 18216
rect 4068 18139 4120 18148
rect 4068 18105 4080 18139
rect 4080 18105 4120 18139
rect 4068 18096 4120 18105
rect 1768 18028 1820 18080
rect 2320 18028 2372 18080
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 5816 18071 5868 18080
rect 5816 18037 5825 18071
rect 5825 18037 5859 18071
rect 5859 18037 5868 18071
rect 5816 18028 5868 18037
rect 6920 18028 6972 18080
rect 8024 18071 8076 18080
rect 8024 18037 8033 18071
rect 8033 18037 8067 18071
rect 8067 18037 8076 18071
rect 8024 18028 8076 18037
rect 9588 18071 9640 18080
rect 9588 18037 9597 18071
rect 9597 18037 9631 18071
rect 9631 18037 9640 18071
rect 9588 18028 9640 18037
rect 11520 18232 11572 18284
rect 10968 18028 11020 18080
rect 11152 18071 11204 18080
rect 11152 18037 11161 18071
rect 11161 18037 11195 18071
rect 11195 18037 11204 18071
rect 11152 18028 11204 18037
rect 11244 18071 11296 18080
rect 11244 18037 11253 18071
rect 11253 18037 11287 18071
rect 11287 18037 11296 18071
rect 11244 18028 11296 18037
rect 11520 18028 11572 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2780 17824 2832 17876
rect 3792 17824 3844 17876
rect 5172 17867 5224 17876
rect 4160 17756 4212 17808
rect 2044 17688 2096 17740
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 7288 17824 7340 17876
rect 7748 17867 7800 17876
rect 7748 17833 7757 17867
rect 7757 17833 7791 17867
rect 7791 17833 7800 17867
rect 7748 17824 7800 17833
rect 9680 17824 9732 17876
rect 11060 17824 11112 17876
rect 6092 17799 6144 17808
rect 6092 17765 6126 17799
rect 6126 17765 6144 17799
rect 6092 17756 6144 17765
rect 5172 17688 5224 17740
rect 9036 17688 9088 17740
rect 2320 17663 2372 17672
rect 2320 17629 2329 17663
rect 2329 17629 2363 17663
rect 2363 17629 2372 17663
rect 2320 17620 2372 17629
rect 2136 17552 2188 17604
rect 4344 17620 4396 17672
rect 4620 17663 4672 17672
rect 4620 17629 4629 17663
rect 4629 17629 4663 17663
rect 4663 17629 4672 17663
rect 5816 17663 5868 17672
rect 4620 17620 4672 17629
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 8300 17663 8352 17672
rect 8300 17629 8309 17663
rect 8309 17629 8343 17663
rect 8343 17629 8352 17663
rect 8300 17620 8352 17629
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 1860 17527 1912 17536
rect 1860 17493 1869 17527
rect 1869 17493 1903 17527
rect 1903 17493 1912 17527
rect 1860 17484 1912 17493
rect 5448 17484 5500 17536
rect 5540 17484 5592 17536
rect 6736 17484 6788 17536
rect 7380 17484 7432 17536
rect 8208 17484 8260 17536
rect 9496 17484 9548 17536
rect 10692 17620 10744 17672
rect 12440 17756 12492 17808
rect 11520 17688 11572 17740
rect 10784 17527 10836 17536
rect 10784 17493 10793 17527
rect 10793 17493 10827 17527
rect 10827 17493 10836 17527
rect 10784 17484 10836 17493
rect 11152 17484 11204 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 4620 17280 4672 17332
rect 6092 17280 6144 17332
rect 9680 17280 9732 17332
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 1676 17144 1728 17196
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 9496 17187 9548 17196
rect 2596 17076 2648 17128
rect 3884 17076 3936 17128
rect 5540 17076 5592 17128
rect 9496 17153 9505 17187
rect 9505 17153 9539 17187
rect 9539 17153 9548 17187
rect 9496 17144 9548 17153
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 7288 17119 7340 17128
rect 7288 17085 7322 17119
rect 7322 17085 7340 17119
rect 3056 17051 3108 17060
rect 3056 17017 3065 17051
rect 3065 17017 3099 17051
rect 3099 17017 3108 17051
rect 3056 17008 3108 17017
rect 1676 16940 1728 16992
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 2136 16940 2188 16992
rect 5172 16983 5224 16992
rect 5172 16949 5181 16983
rect 5181 16949 5215 16983
rect 5215 16949 5224 16983
rect 5172 16940 5224 16949
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 7288 17076 7340 17085
rect 10784 17008 10836 17060
rect 12624 17008 12676 17060
rect 7288 16940 7340 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2412 16779 2464 16788
rect 2412 16745 2421 16779
rect 2421 16745 2455 16779
rect 2455 16745 2464 16779
rect 2412 16736 2464 16745
rect 4252 16736 4304 16788
rect 5448 16736 5500 16788
rect 6828 16736 6880 16788
rect 7564 16736 7616 16788
rect 9128 16736 9180 16788
rect 10140 16736 10192 16788
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 2688 16668 2740 16720
rect 3792 16711 3844 16720
rect 3792 16677 3801 16711
rect 3801 16677 3835 16711
rect 3835 16677 3844 16711
rect 3792 16668 3844 16677
rect 4896 16668 4948 16720
rect 6092 16668 6144 16720
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 2136 16600 2188 16652
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 3516 16643 3568 16652
rect 2780 16600 2832 16609
rect 3516 16609 3525 16643
rect 3525 16609 3559 16643
rect 3559 16609 3568 16643
rect 3516 16600 3568 16609
rect 4344 16643 4396 16652
rect 4344 16609 4353 16643
rect 4353 16609 4387 16643
rect 4387 16609 4396 16643
rect 4344 16600 4396 16609
rect 4528 16600 4580 16652
rect 6000 16600 6052 16652
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 8392 16668 8444 16720
rect 12440 16668 12492 16720
rect 2688 16532 2740 16584
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 6644 16575 6696 16584
rect 6644 16541 6653 16575
rect 6653 16541 6687 16575
rect 6687 16541 6696 16575
rect 6644 16532 6696 16541
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 8024 16532 8076 16584
rect 11888 16600 11940 16652
rect 9496 16532 9548 16584
rect 9956 16532 10008 16584
rect 6092 16396 6144 16448
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 7288 16396 7340 16405
rect 7932 16439 7984 16448
rect 7932 16405 7941 16439
rect 7941 16405 7975 16439
rect 7975 16405 7984 16439
rect 7932 16396 7984 16405
rect 9404 16439 9456 16448
rect 9404 16405 9413 16439
rect 9413 16405 9447 16439
rect 9447 16405 9456 16439
rect 9404 16396 9456 16405
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 10968 16396 11020 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2688 16192 2740 16244
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 7564 16235 7616 16244
rect 7564 16201 7573 16235
rect 7573 16201 7607 16235
rect 7607 16201 7616 16235
rect 7564 16192 7616 16201
rect 10692 16192 10744 16244
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 12440 16192 12492 16244
rect 10232 16124 10284 16176
rect 6000 16056 6052 16108
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 10784 16056 10836 16108
rect 1768 15988 1820 16040
rect 2596 15988 2648 16040
rect 2688 15920 2740 15972
rect 8116 15988 8168 16040
rect 8576 15988 8628 16040
rect 9588 15988 9640 16040
rect 6644 15920 6696 15972
rect 7196 15920 7248 15972
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 5264 15852 5316 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 8024 15852 8076 15904
rect 8852 15852 8904 15904
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10876 15895 10928 15904
rect 10876 15861 10885 15895
rect 10885 15861 10919 15895
rect 10919 15861 10928 15895
rect 10876 15852 10928 15861
rect 10968 15895 11020 15904
rect 10968 15861 10977 15895
rect 10977 15861 11011 15895
rect 11011 15861 11020 15895
rect 10968 15852 11020 15861
rect 11152 15852 11204 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1400 15648 1452 15700
rect 1860 15648 1912 15700
rect 6736 15691 6788 15700
rect 6736 15657 6745 15691
rect 6745 15657 6779 15691
rect 6779 15657 6788 15691
rect 6736 15648 6788 15657
rect 7472 15691 7524 15700
rect 7472 15657 7481 15691
rect 7481 15657 7515 15691
rect 7515 15657 7524 15691
rect 7472 15648 7524 15657
rect 7932 15691 7984 15700
rect 7932 15657 7941 15691
rect 7941 15657 7975 15691
rect 7975 15657 7984 15691
rect 7932 15648 7984 15657
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 10876 15648 10928 15700
rect 11888 15648 11940 15700
rect 12992 15648 13044 15700
rect 14004 15691 14056 15700
rect 14004 15657 14013 15691
rect 14013 15657 14047 15691
rect 14047 15657 14056 15691
rect 14004 15648 14056 15657
rect 1676 15580 1728 15632
rect 7656 15580 7708 15632
rect 8208 15580 8260 15632
rect 11152 15580 11204 15632
rect 4988 15555 5040 15564
rect 4988 15521 5022 15555
rect 5022 15521 5040 15555
rect 4988 15512 5040 15521
rect 3424 15444 3476 15496
rect 3884 15487 3936 15496
rect 3884 15453 3893 15487
rect 3893 15453 3927 15487
rect 3927 15453 3936 15487
rect 3884 15444 3936 15453
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 2688 15419 2740 15428
rect 2688 15385 2697 15419
rect 2697 15385 2731 15419
rect 2731 15385 2740 15419
rect 2688 15376 2740 15385
rect 4252 15376 4304 15428
rect 2780 15308 2832 15360
rect 5356 15308 5408 15360
rect 6920 15308 6972 15360
rect 9312 15512 9364 15564
rect 9680 15512 9732 15564
rect 10876 15512 10928 15564
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 8576 15444 8628 15496
rect 7288 15376 7340 15428
rect 8208 15376 8260 15428
rect 8852 15351 8904 15360
rect 8852 15317 8861 15351
rect 8861 15317 8895 15351
rect 8895 15317 8904 15351
rect 8852 15308 8904 15317
rect 9036 15308 9088 15360
rect 9404 15308 9456 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 3516 15104 3568 15156
rect 7656 15147 7708 15156
rect 7656 15113 7665 15147
rect 7665 15113 7699 15147
rect 7699 15113 7708 15147
rect 7656 15104 7708 15113
rect 8116 15104 8168 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 10140 15104 10192 15156
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 6552 15079 6604 15088
rect 6552 15045 6561 15079
rect 6561 15045 6595 15079
rect 6595 15045 6604 15079
rect 6552 15036 6604 15045
rect 14004 15036 14056 15088
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 4252 14968 4304 15020
rect 4620 14968 4672 15020
rect 5356 14968 5408 15020
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 12440 14968 12492 15020
rect 12992 15011 13044 15020
rect 1768 14900 1820 14952
rect 2412 14875 2464 14884
rect 2412 14841 2421 14875
rect 2421 14841 2455 14875
rect 2455 14841 2464 14875
rect 2412 14832 2464 14841
rect 4896 14900 4948 14952
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 8852 14900 8904 14952
rect 4804 14832 4856 14884
rect 5724 14875 5776 14884
rect 5724 14841 5733 14875
rect 5733 14841 5767 14875
rect 5767 14841 5776 14875
rect 5724 14832 5776 14841
rect 9588 14832 9640 14884
rect 10140 14832 10192 14884
rect 11888 14875 11940 14884
rect 11888 14841 11897 14875
rect 11897 14841 11931 14875
rect 11931 14841 11940 14875
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 11888 14832 11940 14841
rect 14096 14832 14148 14884
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 12164 14764 12216 14773
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 13912 14764 13964 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1400 14603 1452 14612
rect 1400 14569 1409 14603
rect 1409 14569 1443 14603
rect 1443 14569 1452 14603
rect 1400 14560 1452 14569
rect 1676 14560 1728 14612
rect 2412 14560 2464 14612
rect 2872 14560 2924 14612
rect 4068 14560 4120 14612
rect 4620 14603 4672 14612
rect 4620 14569 4629 14603
rect 4629 14569 4663 14603
rect 4663 14569 4672 14603
rect 4620 14560 4672 14569
rect 4988 14560 5040 14612
rect 7932 14560 7984 14612
rect 8852 14603 8904 14612
rect 8852 14569 8861 14603
rect 8861 14569 8895 14603
rect 8895 14569 8904 14603
rect 8852 14560 8904 14569
rect 9496 14560 9548 14612
rect 10140 14560 10192 14612
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 14004 14603 14056 14612
rect 12440 14560 12492 14569
rect 14004 14569 14013 14603
rect 14013 14569 14047 14603
rect 14047 14569 14056 14603
rect 14004 14560 14056 14569
rect 2136 14492 2188 14544
rect 2688 14492 2740 14544
rect 11060 14492 11112 14544
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 4160 14424 4212 14476
rect 5540 14467 5592 14476
rect 5540 14433 5574 14467
rect 5574 14433 5592 14467
rect 5540 14424 5592 14433
rect 7288 14424 7340 14476
rect 10968 14424 11020 14476
rect 11704 14424 11756 14476
rect 23388 14467 23440 14476
rect 23388 14433 23397 14467
rect 23397 14433 23431 14467
rect 23431 14433 23440 14467
rect 23388 14424 23440 14433
rect 2044 14356 2096 14408
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3056 14356 3108 14365
rect 4712 14356 4764 14408
rect 5172 14356 5224 14408
rect 7380 14356 7432 14408
rect 5080 14288 5132 14340
rect 7748 14331 7800 14340
rect 7748 14297 7757 14331
rect 7757 14297 7791 14331
rect 7791 14297 7800 14331
rect 7748 14288 7800 14297
rect 7840 14288 7892 14340
rect 10876 14356 10928 14408
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 9680 14220 9732 14272
rect 24952 14220 25004 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2872 14016 2924 14068
rect 11060 14016 11112 14068
rect 23388 14059 23440 14068
rect 23388 14025 23397 14059
rect 23397 14025 23431 14059
rect 23431 14025 23440 14059
rect 23388 14016 23440 14025
rect 2044 13991 2096 14000
rect 2044 13957 2053 13991
rect 2053 13957 2087 13991
rect 2087 13957 2096 13991
rect 2044 13948 2096 13957
rect 3424 13948 3476 14000
rect 4436 13948 4488 14000
rect 7288 13948 7340 14000
rect 10692 13948 10744 14000
rect 13452 13948 13504 14000
rect 24860 13948 24912 14000
rect 8116 13923 8168 13932
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2688 13812 2740 13864
rect 2872 13812 2924 13864
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 11704 13880 11756 13932
rect 5448 13812 5500 13864
rect 4988 13787 5040 13796
rect 4988 13753 4997 13787
rect 4997 13753 5031 13787
rect 5031 13753 5040 13787
rect 6552 13812 6604 13864
rect 6920 13812 6972 13864
rect 7380 13812 7432 13864
rect 8852 13812 8904 13864
rect 10876 13812 10928 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 10968 13787 11020 13796
rect 4988 13744 5040 13753
rect 10968 13753 10977 13787
rect 10977 13753 11011 13787
rect 11011 13753 11020 13787
rect 10968 13744 11020 13753
rect 2688 13676 2740 13728
rect 3056 13676 3108 13728
rect 4436 13676 4488 13728
rect 5264 13676 5316 13728
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 6460 13719 6512 13728
rect 6460 13685 6469 13719
rect 6469 13685 6503 13719
rect 6503 13685 6512 13719
rect 6460 13676 6512 13685
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 11704 13719 11756 13728
rect 11704 13685 11713 13719
rect 11713 13685 11747 13719
rect 11747 13685 11756 13719
rect 11704 13676 11756 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 5724 13472 5776 13524
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 9680 13472 9732 13524
rect 11704 13472 11756 13524
rect 2596 13404 2648 13456
rect 3056 13404 3108 13456
rect 5264 13447 5316 13456
rect 5264 13413 5273 13447
rect 5273 13413 5307 13447
rect 5307 13413 5316 13447
rect 5264 13404 5316 13413
rect 6368 13404 6420 13456
rect 7656 13404 7708 13456
rect 8576 13404 8628 13456
rect 1584 13336 1636 13388
rect 2136 13336 2188 13388
rect 2780 13336 2832 13388
rect 5172 13336 5224 13388
rect 6000 13336 6052 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 11428 13404 11480 13456
rect 10784 13336 10836 13388
rect 22376 13379 22428 13388
rect 22376 13345 22385 13379
rect 22385 13345 22419 13379
rect 22419 13345 22428 13379
rect 22376 13336 22428 13345
rect 5356 13268 5408 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 7840 13200 7892 13252
rect 1768 13132 1820 13184
rect 2596 13132 2648 13184
rect 3976 13132 4028 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7932 13175 7984 13184
rect 7932 13141 7941 13175
rect 7941 13141 7975 13175
rect 7975 13141 7984 13175
rect 7932 13132 7984 13141
rect 9404 13175 9456 13184
rect 9404 13141 9413 13175
rect 9413 13141 9447 13175
rect 9447 13141 9456 13175
rect 9404 13132 9456 13141
rect 9772 13132 9824 13184
rect 11888 13132 11940 13184
rect 23480 13132 23532 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 2136 12928 2188 12980
rect 2872 12860 2924 12912
rect 4068 12928 4120 12980
rect 5540 12928 5592 12980
rect 6092 12928 6144 12980
rect 6552 12971 6604 12980
rect 6552 12937 6561 12971
rect 6561 12937 6595 12971
rect 6595 12937 6604 12971
rect 6552 12928 6604 12937
rect 7012 12928 7064 12980
rect 8576 12928 8628 12980
rect 8852 12928 8904 12980
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 5080 12860 5132 12912
rect 8300 12860 8352 12912
rect 10784 12903 10836 12912
rect 8116 12792 8168 12844
rect 9680 12792 9732 12844
rect 10784 12869 10793 12903
rect 10793 12869 10827 12903
rect 10827 12869 10836 12903
rect 10784 12860 10836 12869
rect 10968 12860 11020 12912
rect 11888 12792 11940 12844
rect 3516 12724 3568 12776
rect 5816 12724 5868 12776
rect 6460 12724 6512 12776
rect 7472 12724 7524 12776
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 22376 12767 22428 12776
rect 22376 12733 22385 12767
rect 22385 12733 22419 12767
rect 22419 12733 22428 12767
rect 22376 12724 22428 12733
rect 3148 12656 3200 12708
rect 6000 12656 6052 12708
rect 6828 12656 6880 12708
rect 9220 12656 9272 12708
rect 2136 12588 2188 12640
rect 4528 12588 4580 12640
rect 8208 12588 8260 12640
rect 8852 12588 8904 12640
rect 9404 12588 9456 12640
rect 10692 12588 10744 12640
rect 11428 12631 11480 12640
rect 11428 12597 11437 12631
rect 11437 12597 11471 12631
rect 11471 12597 11480 12631
rect 11428 12588 11480 12597
rect 12348 12588 12400 12640
rect 14188 12588 14240 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2688 12384 2740 12436
rect 2964 12427 3016 12436
rect 2964 12393 2973 12427
rect 2973 12393 3007 12427
rect 3007 12393 3016 12427
rect 2964 12384 3016 12393
rect 3424 12427 3476 12436
rect 3424 12393 3433 12427
rect 3433 12393 3467 12427
rect 3467 12393 3476 12427
rect 3424 12384 3476 12393
rect 5816 12427 5868 12436
rect 5816 12393 5825 12427
rect 5825 12393 5859 12427
rect 5859 12393 5868 12427
rect 5816 12384 5868 12393
rect 2872 12316 2924 12368
rect 6920 12384 6972 12436
rect 7564 12384 7616 12436
rect 8484 12384 8536 12436
rect 9220 12384 9272 12436
rect 11060 12384 11112 12436
rect 6276 12316 6328 12368
rect 1768 12291 1820 12300
rect 1768 12257 1777 12291
rect 1777 12257 1811 12291
rect 1811 12257 1820 12291
rect 1768 12248 1820 12257
rect 2780 12248 2832 12300
rect 4160 12248 4212 12300
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 5356 12248 5408 12300
rect 5540 12248 5592 12300
rect 9588 12248 9640 12300
rect 10692 12316 10744 12368
rect 10048 12248 10100 12300
rect 12716 12291 12768 12300
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 5080 12180 5132 12232
rect 12716 12257 12750 12291
rect 12750 12257 12768 12291
rect 12716 12248 12768 12257
rect 21824 12291 21876 12300
rect 21824 12257 21833 12291
rect 21833 12257 21867 12291
rect 21867 12257 21876 12291
rect 21824 12248 21876 12257
rect 12348 12180 12400 12232
rect 4344 12155 4396 12164
rect 4344 12121 4353 12155
rect 4353 12121 4387 12155
rect 4387 12121 4396 12155
rect 4344 12112 4396 12121
rect 2872 12044 2924 12096
rect 3148 12044 3200 12096
rect 6552 12044 6604 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 11888 12044 11940 12096
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 13912 12044 13964 12096
rect 22008 12087 22060 12096
rect 22008 12053 22017 12087
rect 22017 12053 22051 12087
rect 22051 12053 22060 12087
rect 22008 12044 22060 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1492 11840 1544 11892
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 2320 11840 2372 11892
rect 5448 11840 5500 11892
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 8392 11840 8444 11892
rect 12716 11840 12768 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 12440 11815 12492 11824
rect 12440 11781 12449 11815
rect 12449 11781 12483 11815
rect 12483 11781 12492 11815
rect 12440 11772 12492 11781
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 4068 11704 4120 11756
rect 5356 11704 5408 11756
rect 7840 11704 7892 11756
rect 9404 11704 9456 11756
rect 10692 11704 10744 11756
rect 11796 11704 11848 11756
rect 13268 11704 13320 11756
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 2964 11611 3016 11620
rect 2964 11577 2973 11611
rect 2973 11577 3007 11611
rect 3007 11577 3016 11611
rect 2964 11568 3016 11577
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 4528 11611 4580 11620
rect 4528 11577 4562 11611
rect 4562 11577 4580 11611
rect 4528 11568 4580 11577
rect 9864 11636 9916 11688
rect 10140 11679 10192 11688
rect 10140 11645 10149 11679
rect 10149 11645 10183 11679
rect 10183 11645 10192 11679
rect 10140 11636 10192 11645
rect 21824 11679 21876 11688
rect 8484 11568 8536 11620
rect 5080 11500 5132 11552
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 7104 11543 7156 11552
rect 7104 11509 7113 11543
rect 7113 11509 7147 11543
rect 7147 11509 7156 11543
rect 7104 11500 7156 11509
rect 8116 11500 8168 11552
rect 9864 11500 9916 11552
rect 10876 11500 10928 11552
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3056 11296 3108 11348
rect 4528 11296 4580 11348
rect 5816 11296 5868 11348
rect 6276 11296 6328 11348
rect 7104 11296 7156 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 9864 11339 9916 11348
rect 8392 11296 8444 11305
rect 9864 11305 9873 11339
rect 9873 11305 9907 11339
rect 9907 11305 9916 11339
rect 9864 11296 9916 11305
rect 10692 11296 10744 11348
rect 11060 11296 11112 11348
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 1400 11228 1452 11280
rect 5540 11228 5592 11280
rect 7564 11228 7616 11280
rect 11244 11228 11296 11280
rect 13176 11228 13228 11280
rect 1584 11160 1636 11212
rect 2044 11160 2096 11212
rect 4160 11203 4212 11212
rect 4160 11169 4169 11203
rect 4169 11169 4203 11203
rect 4203 11169 4212 11203
rect 4160 11160 4212 11169
rect 5356 11160 5408 11212
rect 10784 11160 10836 11212
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 9588 11092 9640 11144
rect 11428 11092 11480 11144
rect 12716 11135 12768 11144
rect 2872 11024 2924 11076
rect 5264 10999 5316 11008
rect 5264 10965 5273 10999
rect 5273 10965 5307 10999
rect 5307 10965 5316 10999
rect 5264 10956 5316 10965
rect 7472 11024 7524 11076
rect 9496 11024 9548 11076
rect 10048 11024 10100 11076
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 13268 11135 13320 11144
rect 12808 11092 12860 11101
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 9220 10956 9272 11008
rect 11060 10956 11112 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 5632 10684 5684 10736
rect 6552 10752 6604 10804
rect 8852 10795 8904 10804
rect 8852 10761 8861 10795
rect 8861 10761 8895 10795
rect 8895 10761 8904 10795
rect 8852 10752 8904 10761
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 12348 10752 12400 10804
rect 12808 10752 12860 10804
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 4528 10616 4580 10668
rect 6184 10616 6236 10668
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7564 10616 7616 10668
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 5264 10548 5316 10600
rect 7288 10548 7340 10600
rect 7748 10548 7800 10600
rect 9772 10548 9824 10600
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 8760 10480 8812 10532
rect 9036 10480 9088 10532
rect 9864 10480 9916 10532
rect 12900 10523 12952 10532
rect 12900 10489 12909 10523
rect 12909 10489 12943 10523
rect 12943 10489 12952 10523
rect 12900 10480 12952 10489
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 3516 10412 3568 10464
rect 4252 10412 4304 10464
rect 6552 10412 6604 10464
rect 7288 10412 7340 10464
rect 7564 10455 7616 10464
rect 7564 10421 7573 10455
rect 7573 10421 7607 10455
rect 7607 10421 7616 10455
rect 7564 10412 7616 10421
rect 7748 10412 7800 10464
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 11428 10455 11480 10464
rect 11428 10421 11437 10455
rect 11437 10421 11471 10455
rect 11471 10421 11480 10455
rect 11428 10412 11480 10421
rect 12716 10412 12768 10464
rect 13360 10412 13412 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2964 10208 3016 10260
rect 2780 10140 2832 10192
rect 2504 10072 2556 10124
rect 3976 10072 4028 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 4620 10140 4672 10192
rect 5264 10208 5316 10260
rect 6276 10208 6328 10260
rect 8392 10208 8444 10260
rect 8576 10208 8628 10260
rect 4160 10072 4212 10124
rect 5632 10072 5684 10124
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 6460 10072 6512 10124
rect 4344 10004 4396 10056
rect 7288 10140 7340 10192
rect 6920 10072 6972 10124
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 6552 9936 6604 9988
rect 2044 9868 2096 9920
rect 7104 9868 7156 9920
rect 7748 10004 7800 10056
rect 10692 10208 10744 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 9864 10140 9916 10192
rect 10140 10140 10192 10192
rect 9496 10072 9548 10124
rect 11336 10072 11388 10124
rect 8208 10004 8260 10056
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 9772 9936 9824 9988
rect 11244 9936 11296 9988
rect 14556 9936 14608 9988
rect 19340 9936 19392 9988
rect 24124 9936 24176 9988
rect 9036 9868 9088 9920
rect 12164 9868 12216 9920
rect 12808 9911 12860 9920
rect 12808 9877 12817 9911
rect 12817 9877 12851 9911
rect 12851 9877 12860 9911
rect 12808 9868 12860 9877
rect 14280 9868 14332 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1400 9664 1452 9716
rect 2504 9707 2556 9716
rect 2228 9596 2280 9648
rect 1676 9528 1728 9580
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2504 9673 2513 9707
rect 2513 9673 2547 9707
rect 2547 9673 2556 9707
rect 2504 9664 2556 9673
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 5356 9639 5408 9648
rect 5356 9605 5365 9639
rect 5365 9605 5399 9639
rect 5399 9605 5408 9639
rect 6552 9664 6604 9716
rect 5356 9596 5408 9605
rect 8024 9596 8076 9648
rect 2596 9460 2648 9512
rect 5632 9528 5684 9580
rect 6276 9528 6328 9580
rect 6736 9528 6788 9580
rect 9680 9664 9732 9716
rect 11244 9664 11296 9716
rect 12256 9596 12308 9648
rect 12072 9528 12124 9580
rect 13544 9528 13596 9580
rect 4896 9460 4948 9512
rect 3608 9392 3660 9444
rect 6920 9460 6972 9512
rect 7104 9503 7156 9512
rect 7104 9469 7138 9503
rect 7138 9469 7156 9503
rect 7104 9460 7156 9469
rect 8300 9460 8352 9512
rect 9864 9460 9916 9512
rect 12164 9460 12216 9512
rect 12348 9460 12400 9512
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 1860 9367 1912 9376
rect 1860 9333 1869 9367
rect 1869 9333 1903 9367
rect 1903 9333 1912 9367
rect 1860 9324 1912 9333
rect 2228 9324 2280 9376
rect 6092 9392 6144 9444
rect 9496 9392 9548 9444
rect 12716 9392 12768 9444
rect 13912 9435 13964 9444
rect 13912 9401 13921 9435
rect 13921 9401 13955 9435
rect 13955 9401 13964 9435
rect 13912 9392 13964 9401
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 10140 9324 10192 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11520 9324 11572 9376
rect 13544 9367 13596 9376
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 2136 9120 2188 9172
rect 4068 9120 4120 9172
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 1768 9052 1820 9104
rect 3056 9052 3108 9104
rect 8300 9120 8352 9172
rect 9496 9120 9548 9172
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 12808 9120 12860 9172
rect 13912 9163 13964 9172
rect 13912 9129 13921 9163
rect 13921 9129 13955 9163
rect 13955 9129 13964 9163
rect 13912 9120 13964 9129
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 4896 8984 4948 9036
rect 5540 9052 5592 9104
rect 6276 8984 6328 9036
rect 3516 8959 3568 8968
rect 2044 8848 2096 8900
rect 2688 8848 2740 8900
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 7656 8891 7708 8900
rect 1032 8780 1084 8832
rect 3240 8780 3292 8832
rect 3516 8780 3568 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 4620 8823 4672 8832
rect 4620 8789 4629 8823
rect 4629 8789 4663 8823
rect 4663 8789 4672 8823
rect 4620 8780 4672 8789
rect 7656 8857 7665 8891
rect 7665 8857 7699 8891
rect 7699 8857 7708 8891
rect 7656 8848 7708 8857
rect 7748 8780 7800 8832
rect 7932 9052 7984 9104
rect 13544 9052 13596 9104
rect 9312 8984 9364 9036
rect 9588 8984 9640 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 11244 8984 11296 9036
rect 13452 8984 13504 9036
rect 14280 8984 14332 9036
rect 15568 9027 15620 9036
rect 15568 8993 15602 9027
rect 15602 8993 15620 9027
rect 15568 8984 15620 8993
rect 7932 8916 7984 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8392 8916 8444 8968
rect 9864 8916 9916 8968
rect 10692 8916 10744 8968
rect 8300 8848 8352 8900
rect 9404 8848 9456 8900
rect 12808 8891 12860 8900
rect 12808 8857 12817 8891
rect 12817 8857 12851 8891
rect 12851 8857 12860 8891
rect 12808 8848 12860 8857
rect 14556 8848 14608 8900
rect 8208 8780 8260 8832
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 9772 8780 9824 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 5356 8576 5408 8628
rect 6276 8619 6328 8628
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 8024 8576 8076 8628
rect 8484 8576 8536 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 10048 8576 10100 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 11796 8619 11848 8628
rect 10140 8576 10192 8585
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 4896 8551 4948 8560
rect 4896 8517 4905 8551
rect 4905 8517 4939 8551
rect 4939 8517 4948 8551
rect 4896 8508 4948 8517
rect 6828 8551 6880 8560
rect 6828 8517 6837 8551
rect 6837 8517 6871 8551
rect 6871 8517 6880 8551
rect 6828 8508 6880 8517
rect 8576 8551 8628 8560
rect 8576 8517 8585 8551
rect 8585 8517 8619 8551
rect 8619 8517 8628 8551
rect 8576 8508 8628 8517
rect 10232 8508 10284 8560
rect 11980 8508 12032 8560
rect 13820 8508 13872 8560
rect 15200 8508 15252 8560
rect 15568 8551 15620 8560
rect 15568 8517 15577 8551
rect 15577 8517 15611 8551
rect 15611 8517 15620 8551
rect 15568 8508 15620 8517
rect 1400 8440 1452 8492
rect 4988 8440 5040 8492
rect 7012 8440 7064 8492
rect 8944 8440 8996 8492
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 13084 8440 13136 8492
rect 4896 8372 4948 8424
rect 8852 8372 8904 8424
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11796 8372 11848 8424
rect 1308 8304 1360 8356
rect 2044 8347 2096 8356
rect 2044 8313 2053 8347
rect 2053 8313 2087 8347
rect 2087 8313 2096 8347
rect 2044 8304 2096 8313
rect 2136 8304 2188 8356
rect 1584 8236 1636 8288
rect 1768 8236 1820 8288
rect 2596 8304 2648 8356
rect 5264 8304 5316 8356
rect 6552 8347 6604 8356
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 7104 8304 7156 8356
rect 7932 8304 7984 8356
rect 8760 8304 8812 8356
rect 9588 8304 9640 8356
rect 10784 8304 10836 8356
rect 11336 8304 11388 8356
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 20260 8415 20312 8424
rect 14188 8372 14240 8381
rect 20260 8381 20269 8415
rect 20269 8381 20303 8415
rect 20303 8381 20312 8415
rect 20260 8372 20312 8381
rect 14464 8347 14516 8356
rect 14464 8313 14498 8347
rect 14498 8313 14516 8347
rect 14464 8304 14516 8313
rect 16672 8347 16724 8356
rect 16672 8313 16681 8347
rect 16681 8313 16715 8347
rect 16715 8313 16724 8347
rect 16672 8304 16724 8313
rect 20352 8304 20404 8356
rect 2688 8236 2740 8288
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 5448 8236 5500 8288
rect 6920 8236 6972 8288
rect 8116 8236 8168 8288
rect 9220 8236 9272 8288
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 12992 8236 13044 8288
rect 13452 8236 13504 8288
rect 14188 8236 14240 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 4068 8032 4120 8084
rect 3792 8007 3844 8016
rect 3792 7973 3801 8007
rect 3801 7973 3835 8007
rect 3835 7973 3844 8007
rect 4804 8032 4856 8084
rect 7196 8032 7248 8084
rect 8668 8032 8720 8084
rect 8944 8032 8996 8084
rect 9496 8032 9548 8084
rect 9680 8075 9732 8084
rect 9680 8041 9689 8075
rect 9689 8041 9723 8075
rect 9723 8041 9732 8075
rect 9680 8032 9732 8041
rect 10692 8032 10744 8084
rect 13084 8075 13136 8084
rect 13084 8041 13093 8075
rect 13093 8041 13127 8075
rect 13127 8041 13136 8075
rect 13084 8032 13136 8041
rect 13820 8032 13872 8084
rect 14188 8032 14240 8084
rect 15844 8032 15896 8084
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 3792 7964 3844 7973
rect 5356 7964 5408 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 1676 7939 1728 7948
rect 1676 7905 1710 7939
rect 1710 7905 1728 7939
rect 1676 7896 1728 7905
rect 5172 7896 5224 7948
rect 7564 7896 7616 7948
rect 8300 7964 8352 8016
rect 8392 7964 8444 8016
rect 10784 7964 10836 8016
rect 11060 7964 11112 8016
rect 8116 7939 8168 7948
rect 8116 7905 8125 7939
rect 8125 7905 8159 7939
rect 8159 7905 8168 7939
rect 8116 7896 8168 7905
rect 9404 7896 9456 7948
rect 11612 7896 11664 7948
rect 13268 7896 13320 7948
rect 15844 7896 15896 7948
rect 17316 7896 17368 7948
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 7196 7828 7248 7880
rect 3332 7760 3384 7812
rect 5448 7760 5500 7812
rect 7656 7760 7708 7812
rect 9956 7828 10008 7880
rect 12900 7828 12952 7880
rect 15200 7828 15252 7880
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 4896 7692 4948 7701
rect 6736 7692 6788 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 12348 7760 12400 7812
rect 14648 7760 14700 7812
rect 12440 7735 12492 7744
rect 12440 7701 12449 7735
rect 12449 7701 12483 7735
rect 12483 7701 12492 7735
rect 12440 7692 12492 7701
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 16948 7692 17000 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 5172 7488 5224 7540
rect 8116 7488 8168 7540
rect 12900 7531 12952 7540
rect 12900 7497 12909 7531
rect 12909 7497 12943 7531
rect 12943 7497 12952 7531
rect 12900 7488 12952 7497
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 15844 7531 15896 7540
rect 15844 7497 15853 7531
rect 15853 7497 15887 7531
rect 15887 7497 15896 7531
rect 15844 7488 15896 7497
rect 7012 7420 7064 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5356 7352 5408 7404
rect 12532 7420 12584 7472
rect 13360 7420 13412 7472
rect 2596 7284 2648 7336
rect 3056 7327 3108 7336
rect 3056 7293 3090 7327
rect 3090 7293 3108 7327
rect 3056 7284 3108 7293
rect 6920 7284 6972 7336
rect 7656 7327 7708 7336
rect 7656 7293 7690 7327
rect 7690 7293 7708 7327
rect 7656 7284 7708 7293
rect 12164 7352 12216 7404
rect 12992 7352 13044 7404
rect 16948 7395 17000 7404
rect 8208 7216 8260 7268
rect 10692 7284 10744 7336
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 13452 7284 13504 7336
rect 19708 7327 19760 7336
rect 19708 7293 19717 7327
rect 19717 7293 19751 7327
rect 19751 7293 19760 7327
rect 19708 7284 19760 7293
rect 9956 7216 10008 7268
rect 16212 7259 16264 7268
rect 16212 7225 16221 7259
rect 16221 7225 16255 7259
rect 16255 7225 16264 7259
rect 16212 7216 16264 7225
rect 20720 7216 20772 7268
rect 5448 7148 5500 7200
rect 5540 7148 5592 7200
rect 6092 7148 6144 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 11060 7148 11112 7200
rect 14004 7148 14056 7200
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 16580 7148 16632 7200
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 17316 7148 17368 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 4896 6944 4948 6996
rect 5448 6876 5500 6928
rect 2688 6808 2740 6860
rect 3056 6808 3108 6860
rect 7564 6944 7616 6996
rect 7656 6944 7708 6996
rect 11612 6987 11664 6996
rect 11612 6953 11621 6987
rect 11621 6953 11655 6987
rect 11655 6953 11664 6987
rect 11612 6944 11664 6953
rect 13452 6987 13504 6996
rect 13452 6953 13461 6987
rect 13461 6953 13495 6987
rect 13495 6953 13504 6987
rect 13452 6944 13504 6953
rect 13820 6944 13872 6996
rect 6644 6808 6696 6860
rect 7472 6876 7524 6928
rect 10600 6876 10652 6928
rect 10876 6919 10928 6928
rect 10876 6885 10885 6919
rect 10885 6885 10919 6919
rect 10919 6885 10928 6919
rect 10876 6876 10928 6885
rect 6920 6808 6972 6860
rect 7380 6808 7432 6860
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 5356 6740 5408 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 2412 6715 2464 6724
rect 2412 6681 2421 6715
rect 2421 6681 2455 6715
rect 2455 6681 2464 6715
rect 2412 6672 2464 6681
rect 6736 6672 6788 6724
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 4620 6604 4672 6656
rect 5264 6604 5316 6656
rect 10416 6740 10468 6792
rect 11336 6876 11388 6928
rect 12440 6876 12492 6928
rect 12164 6808 12216 6860
rect 14648 6808 14700 6860
rect 15384 6851 15436 6860
rect 15384 6817 15393 6851
rect 15393 6817 15427 6851
rect 15427 6817 15436 6851
rect 15384 6808 15436 6817
rect 16764 6876 16816 6928
rect 17868 6876 17920 6928
rect 16948 6808 17000 6860
rect 20720 6808 20772 6860
rect 15660 6783 15712 6792
rect 9956 6672 10008 6724
rect 10784 6672 10836 6724
rect 10876 6672 10928 6724
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 14004 6672 14056 6724
rect 10508 6647 10560 6656
rect 10508 6613 10517 6647
rect 10517 6613 10551 6647
rect 10551 6613 10560 6647
rect 10508 6604 10560 6613
rect 17500 6604 17552 6656
rect 21640 6604 21692 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2964 6400 3016 6452
rect 5356 6443 5408 6452
rect 5356 6409 5365 6443
rect 5365 6409 5399 6443
rect 5399 6409 5408 6443
rect 5356 6400 5408 6409
rect 5448 6400 5500 6452
rect 9496 6400 9548 6452
rect 10600 6400 10652 6452
rect 11428 6400 11480 6452
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 15384 6400 15436 6452
rect 16948 6400 17000 6452
rect 17408 6400 17460 6452
rect 20720 6400 20772 6452
rect 12348 6332 12400 6384
rect 2044 6264 2096 6316
rect 2780 6264 2832 6316
rect 4344 6264 4396 6316
rect 4712 6264 4764 6316
rect 6828 6264 6880 6316
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8300 6264 8352 6316
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 14004 6264 14056 6316
rect 17868 6264 17920 6316
rect 1676 6196 1728 6248
rect 3424 6196 3476 6248
rect 4252 6196 4304 6248
rect 6736 6196 6788 6248
rect 14740 6196 14792 6248
rect 1400 6060 1452 6112
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2596 6060 2648 6112
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 5448 6128 5500 6180
rect 6920 6128 6972 6180
rect 8576 6128 8628 6180
rect 10416 6128 10468 6180
rect 11336 6171 11388 6180
rect 11336 6137 11345 6171
rect 11345 6137 11379 6171
rect 11379 6137 11388 6171
rect 11336 6128 11388 6137
rect 14280 6128 14332 6180
rect 4344 6060 4396 6112
rect 7564 6060 7616 6112
rect 9864 6060 9916 6112
rect 16764 6196 16816 6248
rect 17592 6128 17644 6180
rect 19432 6171 19484 6180
rect 19432 6137 19441 6171
rect 19441 6137 19475 6171
rect 19475 6137 19484 6171
rect 19432 6128 19484 6137
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 16948 6060 17000 6112
rect 18144 6060 18196 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1676 5856 1728 5908
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 3792 5899 3844 5908
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 4068 5856 4120 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 6828 5899 6880 5908
rect 6828 5865 6837 5899
rect 6837 5865 6871 5899
rect 6871 5865 6880 5899
rect 6828 5856 6880 5865
rect 8852 5856 8904 5908
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 10876 5856 10928 5908
rect 12992 5856 13044 5908
rect 13452 5856 13504 5908
rect 13636 5899 13688 5908
rect 13636 5865 13645 5899
rect 13645 5865 13679 5899
rect 13679 5865 13688 5899
rect 13636 5856 13688 5865
rect 13728 5856 13780 5908
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 14648 5899 14700 5908
rect 14648 5865 14657 5899
rect 14657 5865 14691 5899
rect 14691 5865 14700 5899
rect 14648 5856 14700 5865
rect 16580 5899 16632 5908
rect 16580 5865 16589 5899
rect 16589 5865 16623 5899
rect 16623 5865 16632 5899
rect 16580 5856 16632 5865
rect 17224 5899 17276 5908
rect 17224 5865 17233 5899
rect 17233 5865 17267 5899
rect 17267 5865 17276 5899
rect 17224 5856 17276 5865
rect 1124 5788 1176 5840
rect 2688 5788 2740 5840
rect 8392 5788 8444 5840
rect 8760 5788 8812 5840
rect 11152 5831 11204 5840
rect 11152 5797 11186 5831
rect 11186 5797 11204 5831
rect 11152 5788 11204 5797
rect 18880 5788 18932 5840
rect 1400 5720 1452 5772
rect 5540 5720 5592 5772
rect 6276 5720 6328 5772
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 17960 5720 18012 5772
rect 1952 5516 2004 5568
rect 5264 5652 5316 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 10784 5652 10836 5704
rect 13820 5652 13872 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 16764 5627 16816 5636
rect 16764 5593 16773 5627
rect 16773 5593 16807 5627
rect 16807 5593 16816 5627
rect 16764 5584 16816 5593
rect 17408 5584 17460 5636
rect 19340 5584 19392 5636
rect 5356 5516 5408 5568
rect 8208 5516 8260 5568
rect 11888 5516 11940 5568
rect 17960 5516 18012 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1860 5312 1912 5364
rect 2780 5312 2832 5364
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 7380 5355 7432 5364
rect 7380 5321 7389 5355
rect 7389 5321 7423 5355
rect 7423 5321 7432 5355
rect 7380 5312 7432 5321
rect 9496 5312 9548 5364
rect 11152 5312 11204 5364
rect 13636 5355 13688 5364
rect 13636 5321 13645 5355
rect 13645 5321 13679 5355
rect 13679 5321 13688 5355
rect 13636 5312 13688 5321
rect 14280 5312 14332 5364
rect 14740 5312 14792 5364
rect 2964 5244 3016 5296
rect 3148 5244 3200 5296
rect 4988 5176 5040 5228
rect 5540 5176 5592 5228
rect 6000 5176 6052 5228
rect 6828 5176 6880 5228
rect 8944 5176 8996 5228
rect 13728 5244 13780 5296
rect 1492 5040 1544 5092
rect 1952 5040 2004 5092
rect 6460 5108 6512 5160
rect 8392 5108 8444 5160
rect 12716 5176 12768 5228
rect 13452 5176 13504 5228
rect 14188 5151 14240 5160
rect 3148 4972 3200 5024
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5356 4972 5408 5024
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 17316 5312 17368 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 19340 5312 19392 5364
rect 16856 5108 16908 5160
rect 17776 5151 17828 5160
rect 17776 5117 17785 5151
rect 17785 5117 17819 5151
rect 17819 5117 17828 5151
rect 17776 5108 17828 5117
rect 18144 5108 18196 5160
rect 19432 5108 19484 5160
rect 10784 5040 10836 5092
rect 12348 5040 12400 5092
rect 12716 5040 12768 5092
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 14464 5040 14516 5049
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6920 5015 6972 5024
rect 6920 4981 6929 5015
rect 6929 4981 6963 5015
rect 6963 4981 6972 5015
rect 6920 4972 6972 4981
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 8576 4972 8628 5024
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 9588 4972 9640 5024
rect 15016 4972 15068 5024
rect 17960 5040 18012 5092
rect 17500 4972 17552 5024
rect 22100 4972 22152 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 6000 4768 6052 4820
rect 6184 4768 6236 4820
rect 6276 4768 6328 4820
rect 8576 4768 8628 4820
rect 13728 4811 13780 4820
rect 13728 4777 13737 4811
rect 13737 4777 13771 4811
rect 13771 4777 13780 4811
rect 13728 4768 13780 4777
rect 15384 4768 15436 4820
rect 17224 4768 17276 4820
rect 18144 4768 18196 4820
rect 4344 4700 4396 4752
rect 1492 4675 1544 4684
rect 1492 4641 1501 4675
rect 1501 4641 1535 4675
rect 1535 4641 1544 4675
rect 1492 4632 1544 4641
rect 2228 4632 2280 4684
rect 4160 4632 4212 4684
rect 5540 4675 5592 4684
rect 5540 4641 5574 4675
rect 5574 4641 5592 4675
rect 5540 4632 5592 4641
rect 7748 4700 7800 4752
rect 8760 4700 8812 4752
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 8852 4632 8904 4684
rect 15016 4700 15068 4752
rect 15476 4700 15528 4752
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 10784 4632 10836 4684
rect 11888 4675 11940 4684
rect 11888 4641 11922 4675
rect 11922 4641 11940 4675
rect 11888 4632 11940 4641
rect 14464 4632 14516 4684
rect 15200 4632 15252 4684
rect 16856 4632 16908 4684
rect 17592 4632 17644 4684
rect 19340 4632 19392 4684
rect 21088 4632 21140 4684
rect 8208 4496 8260 4548
rect 9680 4564 9732 4616
rect 10968 4564 11020 4616
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 16212 4564 16264 4616
rect 9864 4496 9916 4548
rect 12992 4539 13044 4548
rect 12992 4505 13001 4539
rect 13001 4505 13035 4539
rect 13035 4505 13044 4539
rect 12992 4496 13044 4505
rect 1860 4428 1912 4480
rect 3148 4428 3200 4480
rect 5264 4428 5316 4480
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 8392 4428 8444 4480
rect 14188 4496 14240 4548
rect 14280 4471 14332 4480
rect 14280 4437 14289 4471
rect 14289 4437 14323 4471
rect 14323 4437 14332 4471
rect 14280 4428 14332 4437
rect 17960 4428 18012 4480
rect 18880 4428 18932 4480
rect 19432 4471 19484 4480
rect 19432 4437 19441 4471
rect 19441 4437 19475 4471
rect 19475 4437 19484 4471
rect 19432 4428 19484 4437
rect 19892 4471 19944 4480
rect 19892 4437 19901 4471
rect 19901 4437 19935 4471
rect 19935 4437 19944 4471
rect 19892 4428 19944 4437
rect 20996 4428 21048 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2780 4224 2832 4276
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 2964 4088 3016 4140
rect 7564 4224 7616 4276
rect 8392 4224 8444 4276
rect 8484 4224 8536 4276
rect 9496 4224 9548 4276
rect 10876 4267 10928 4276
rect 10876 4233 10885 4267
rect 10885 4233 10919 4267
rect 10919 4233 10928 4267
rect 10876 4224 10928 4233
rect 14464 4267 14516 4276
rect 14464 4233 14473 4267
rect 14473 4233 14507 4267
rect 14507 4233 14516 4267
rect 14464 4224 14516 4233
rect 5540 4156 5592 4208
rect 2320 4020 2372 4072
rect 3148 4020 3200 4072
rect 5264 4088 5316 4140
rect 5540 4020 5592 4072
rect 6552 4020 6604 4072
rect 10048 4156 10100 4208
rect 9864 4088 9916 4140
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 5540 3884 5592 3936
rect 6736 3884 6788 3936
rect 10692 4020 10744 4072
rect 15292 4156 15344 4208
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 17868 4088 17920 4140
rect 18788 4088 18840 4140
rect 19432 4156 19484 4208
rect 19892 4156 19944 4208
rect 19524 4131 19576 4140
rect 19524 4097 19533 4131
rect 19533 4097 19567 4131
rect 19567 4097 19576 4131
rect 19524 4088 19576 4097
rect 12992 4020 13044 4072
rect 17592 4020 17644 4072
rect 19064 4063 19116 4072
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 20720 4020 20772 4072
rect 13268 3952 13320 4004
rect 16028 3952 16080 4004
rect 16672 3952 16724 4004
rect 18420 3995 18472 4004
rect 18420 3961 18429 3995
rect 18429 3961 18463 3995
rect 18463 3961 18472 3995
rect 18420 3952 18472 3961
rect 20444 3952 20496 4004
rect 22284 3995 22336 4004
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 11060 3884 11112 3936
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 13544 3884 13596 3936
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 19524 3884 19576 3936
rect 21088 3884 21140 3936
rect 22284 3961 22293 3995
rect 22293 3961 22327 3995
rect 22327 3961 22336 3995
rect 22284 3952 22336 3961
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2412 3680 2464 3732
rect 8208 3680 8260 3732
rect 8760 3680 8812 3732
rect 9588 3680 9640 3732
rect 12164 3723 12216 3732
rect 12164 3689 12173 3723
rect 12173 3689 12207 3723
rect 12207 3689 12216 3723
rect 12164 3680 12216 3689
rect 16672 3723 16724 3732
rect 16672 3689 16681 3723
rect 16681 3689 16715 3723
rect 16715 3689 16724 3723
rect 16672 3680 16724 3689
rect 16856 3680 16908 3732
rect 17408 3680 17460 3732
rect 2320 3612 2372 3664
rect 2688 3655 2740 3664
rect 2688 3621 2697 3655
rect 2697 3621 2731 3655
rect 2731 3621 2740 3655
rect 2688 3612 2740 3621
rect 8392 3655 8444 3664
rect 8392 3621 8401 3655
rect 8401 3621 8435 3655
rect 8435 3621 8444 3655
rect 8392 3612 8444 3621
rect 9864 3612 9916 3664
rect 17500 3612 17552 3664
rect 2044 3544 2096 3596
rect 3424 3544 3476 3596
rect 5264 3544 5316 3596
rect 6276 3544 6328 3596
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 2504 3408 2556 3460
rect 6460 3408 6512 3460
rect 3976 3340 4028 3392
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 6736 3340 6788 3392
rect 11612 3544 11664 3596
rect 12532 3587 12584 3596
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 14740 3544 14792 3596
rect 16396 3544 16448 3596
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 11796 3476 11848 3528
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 14096 3519 14148 3528
rect 12716 3476 12768 3485
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 18512 3680 18564 3732
rect 19524 3680 19576 3732
rect 19432 3612 19484 3664
rect 20904 3587 20956 3596
rect 11612 3408 11664 3460
rect 13268 3451 13320 3460
rect 13268 3417 13277 3451
rect 13277 3417 13311 3451
rect 13311 3417 13320 3451
rect 13268 3408 13320 3417
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 22008 3587 22060 3596
rect 22008 3553 22017 3587
rect 22017 3553 22051 3587
rect 22051 3553 22060 3587
rect 22008 3544 22060 3553
rect 24032 3587 24084 3596
rect 24032 3553 24041 3587
rect 24041 3553 24075 3587
rect 24075 3553 24084 3587
rect 24032 3544 24084 3553
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 19432 3408 19484 3460
rect 9680 3340 9732 3392
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 20720 3340 20772 3392
rect 21548 3340 21600 3392
rect 24216 3383 24268 3392
rect 24216 3349 24225 3383
rect 24225 3349 24259 3383
rect 24259 3349 24268 3383
rect 24216 3340 24268 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 3976 3179 4028 3188
rect 3976 3145 3985 3179
rect 3985 3145 4019 3179
rect 4019 3145 4028 3179
rect 3976 3136 4028 3145
rect 4436 3136 4488 3188
rect 5172 3111 5224 3120
rect 5172 3077 5181 3111
rect 5181 3077 5215 3111
rect 5215 3077 5224 3111
rect 5172 3068 5224 3077
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6736 3000 6788 3052
rect 3148 2932 3200 2984
rect 4344 2932 4396 2984
rect 5540 2975 5592 2984
rect 5540 2941 5549 2975
rect 5549 2941 5583 2975
rect 5583 2941 5592 2975
rect 5540 2932 5592 2941
rect 6460 2932 6512 2984
rect 8484 3136 8536 3188
rect 9864 3136 9916 3188
rect 11244 3136 11296 3188
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12532 3136 12584 3188
rect 12716 3179 12768 3188
rect 12716 3145 12725 3179
rect 12725 3145 12759 3179
rect 12759 3145 12768 3179
rect 12716 3136 12768 3145
rect 14740 3136 14792 3188
rect 15568 3179 15620 3188
rect 15568 3145 15577 3179
rect 15577 3145 15611 3179
rect 15611 3145 15620 3179
rect 17408 3179 17460 3188
rect 15568 3136 15620 3145
rect 9772 3068 9824 3120
rect 11428 3111 11480 3120
rect 11428 3077 11437 3111
rect 11437 3077 11471 3111
rect 11471 3077 11480 3111
rect 11428 3068 11480 3077
rect 1216 2864 1268 2916
rect 2688 2864 2740 2916
rect 3056 2864 3108 2916
rect 5724 2864 5776 2916
rect 6276 2907 6328 2916
rect 6276 2873 6285 2907
rect 6285 2873 6319 2907
rect 6319 2873 6328 2907
rect 11060 3000 11112 3052
rect 15752 3068 15804 3120
rect 8944 2975 8996 2984
rect 8944 2941 8978 2975
rect 8978 2941 8996 2975
rect 8944 2932 8996 2941
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 13544 2975 13596 2984
rect 13544 2941 13578 2975
rect 13578 2941 13596 2975
rect 13544 2932 13596 2941
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 18144 3136 18196 3188
rect 18328 3136 18380 3188
rect 20812 3179 20864 3188
rect 20812 3145 20821 3179
rect 20821 3145 20855 3179
rect 20855 3145 20864 3179
rect 20812 3136 20864 3145
rect 20904 3136 20956 3188
rect 22008 3179 22060 3188
rect 22008 3145 22017 3179
rect 22017 3145 22051 3179
rect 22051 3145 22060 3179
rect 22008 3136 22060 3145
rect 23572 3136 23624 3188
rect 24032 3136 24084 3188
rect 19340 3068 19392 3120
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 23204 3068 23256 3120
rect 17960 2932 18012 2984
rect 19984 2932 20036 2984
rect 20812 2932 20864 2984
rect 22192 2975 22244 2984
rect 22192 2941 22201 2975
rect 22201 2941 22235 2975
rect 22235 2941 22244 2975
rect 22192 2932 22244 2941
rect 23572 2932 23624 2984
rect 6276 2864 6328 2873
rect 8760 2864 8812 2916
rect 20628 2864 20680 2916
rect 204 2796 256 2848
rect 2412 2796 2464 2848
rect 6552 2796 6604 2848
rect 8484 2796 8536 2848
rect 9128 2796 9180 2848
rect 15752 2839 15804 2848
rect 15752 2805 15761 2839
rect 15761 2805 15795 2839
rect 15795 2805 15804 2839
rect 15752 2796 15804 2805
rect 20168 2796 20220 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2228 2592 2280 2644
rect 2504 2635 2556 2644
rect 2504 2601 2513 2635
rect 2513 2601 2547 2635
rect 2547 2601 2556 2635
rect 2504 2592 2556 2601
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 6276 2592 6328 2644
rect 9220 2635 9272 2644
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 9680 2592 9732 2644
rect 9956 2592 10008 2644
rect 10692 2592 10744 2644
rect 11336 2635 11388 2644
rect 11336 2601 11345 2635
rect 11345 2601 11379 2635
rect 11379 2601 11388 2635
rect 11336 2592 11388 2601
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 13728 2635 13780 2644
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 15752 2592 15804 2644
rect 17960 2592 18012 2644
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 1676 2524 1728 2576
rect 4620 2567 4672 2576
rect 4620 2533 4654 2567
rect 4654 2533 4672 2567
rect 4620 2524 4672 2533
rect 10140 2567 10192 2576
rect 10140 2533 10149 2567
rect 10149 2533 10183 2567
rect 10183 2533 10192 2567
rect 10140 2524 10192 2533
rect 4344 2499 4396 2508
rect 4344 2465 4353 2499
rect 4353 2465 4387 2499
rect 4387 2465 4396 2499
rect 4344 2456 4396 2465
rect 6644 2456 6696 2508
rect 7564 2456 7616 2508
rect 15384 2524 15436 2576
rect 20536 2524 20588 2576
rect 21088 2524 21140 2576
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 7196 2388 7248 2440
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 8668 2431 8720 2440
rect 7472 2388 7524 2397
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 12440 2456 12492 2508
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 15200 2499 15252 2508
rect 15200 2465 15209 2499
rect 15209 2465 15243 2499
rect 15243 2465 15252 2499
rect 15200 2456 15252 2465
rect 16212 2456 16264 2508
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 19340 2456 19392 2508
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 22468 2499 22520 2508
rect 22468 2465 22477 2499
rect 22477 2465 22511 2499
rect 22511 2465 22520 2499
rect 22468 2456 22520 2465
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 13084 2431 13136 2440
rect 12072 2388 12124 2397
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 13728 2388 13780 2440
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 2596 2320 2648 2372
rect 8392 2320 8444 2372
rect 12440 2363 12492 2372
rect 12440 2329 12449 2363
rect 12449 2329 12483 2363
rect 12483 2329 12492 2363
rect 15476 2363 15528 2372
rect 12440 2320 12492 2329
rect 15476 2329 15485 2363
rect 15485 2329 15519 2363
rect 15519 2329 15528 2363
rect 15476 2320 15528 2329
rect 16120 2320 16172 2372
rect 9404 2252 9456 2304
rect 9956 2252 10008 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 15384 2252 15436 2304
rect 22652 2295 22704 2304
rect 22652 2261 22661 2295
rect 22661 2261 22695 2295
rect 22695 2261 22704 2295
rect 22652 2252 22704 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 11980 1980 12032 2032
rect 14924 1980 14976 2032
rect 23480 1980 23532 2032
rect 24308 1980 24360 2032
rect 6736 552 6788 604
rect 6828 552 6880 604
rect 7840 552 7892 604
rect 8116 552 8168 604
rect 12164 552 12216 604
rect 12256 552 12308 604
rect 13820 552 13872 604
rect 13912 552 13964 604
rect 24952 552 25004 604
rect 25412 552 25464 604
rect 26240 552 26292 604
rect 27068 552 27120 604
<< metal2 >>
rect 3238 27704 3294 27713
rect 3238 27639 3294 27648
rect 1582 26616 1638 26625
rect 1582 26551 1638 26560
rect 1596 25498 1624 26551
rect 3252 26382 3280 27639
rect 7010 27520 7066 28000
rect 20994 27520 21050 28000
rect 4158 27160 4214 27169
rect 4158 27095 4214 27104
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3146 26072 3202 26081
rect 3146 26007 3202 26016
rect 1584 25492 1636 25498
rect 1584 25434 1636 25440
rect 2686 25392 2742 25401
rect 2596 25356 2648 25362
rect 2686 25327 2742 25336
rect 2596 25298 2648 25304
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1596 24614 1624 24783
rect 2608 24614 2636 25298
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1596 24313 1624 24346
rect 1582 24304 1638 24313
rect 1400 24268 1452 24274
rect 1582 24239 1638 24248
rect 1400 24210 1452 24216
rect 1412 23866 1440 24210
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1400 23860 1452 23866
rect 1400 23802 1452 23808
rect 1688 23662 1716 24006
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1676 23656 1728 23662
rect 1676 23598 1728 23604
rect 1688 23497 1716 23598
rect 1674 23488 1730 23497
rect 1674 23423 1730 23432
rect 1872 22642 1900 23802
rect 1964 23254 1992 24550
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2516 23866 2544 24210
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 1952 23248 2004 23254
rect 1952 23190 2004 23196
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 2410 22536 2466 22545
rect 2410 22471 2412 22480
rect 2464 22471 2466 22480
rect 2412 22442 2464 22448
rect 2608 21865 2636 24550
rect 2700 24410 2728 25327
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 3160 23866 3188 26007
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3054 23760 3110 23769
rect 3054 23695 3110 23704
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 22438 2820 23122
rect 3068 22778 3096 23695
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 3620 23361 3648 23462
rect 3606 23352 3662 23361
rect 4172 23322 4200 27095
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 7024 23866 7052 27520
rect 10048 26376 10100 26382
rect 10048 26318 10100 26324
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 7470 23624 7526 23633
rect 7470 23559 7472 23568
rect 7524 23559 7526 23568
rect 7472 23530 7524 23536
rect 9218 23488 9274 23497
rect 9218 23423 9274 23432
rect 6274 23352 6330 23361
rect 3606 23287 3662 23296
rect 4160 23316 4212 23322
rect 6274 23287 6330 23296
rect 4160 23258 4212 23264
rect 4250 23216 4306 23225
rect 3976 23180 4028 23186
rect 4250 23151 4306 23160
rect 3976 23122 4028 23128
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2792 22137 2820 22374
rect 2778 22128 2834 22137
rect 2778 22063 2834 22072
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 2594 21856 2650 21865
rect 2594 21791 2650 21800
rect 1950 21448 2006 21457
rect 1950 21383 1952 21392
rect 2004 21383 2006 21392
rect 1952 21354 2004 21360
rect 2976 21350 3004 21966
rect 3160 21554 3188 22510
rect 3988 22438 4016 23122
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3988 22166 4016 22374
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3976 22024 4028 22030
rect 3514 21992 3570 22001
rect 3976 21966 4028 21972
rect 3514 21927 3570 21936
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1504 18970 1532 19858
rect 2332 19718 2360 20946
rect 2516 20505 2544 21286
rect 2976 21049 3004 21286
rect 3528 21146 3556 21927
rect 3988 21350 4016 21966
rect 4264 21962 4292 23151
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 4434 22400 4490 22409
rect 4434 22335 4490 22344
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4448 21690 4476 22335
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4252 21480 4304 21486
rect 4250 21448 4252 21457
rect 4304 21448 4306 21457
rect 4250 21383 4306 21392
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 5538 21312 5594 21321
rect 3804 21185 3832 21286
rect 3790 21176 3846 21185
rect 3516 21140 3568 21146
rect 3790 21111 3846 21120
rect 3516 21082 3568 21088
rect 3988 21078 4016 21286
rect 5538 21247 5594 21256
rect 3976 21072 4028 21078
rect 2962 21040 3018 21049
rect 2872 21004 2924 21010
rect 3976 21014 4028 21020
rect 2962 20975 3018 20984
rect 4068 21004 4120 21010
rect 2872 20946 2924 20952
rect 4068 20946 4120 20952
rect 2502 20496 2558 20505
rect 2884 20466 2912 20946
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2502 20431 2558 20440
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 3068 20369 3096 20742
rect 3054 20360 3110 20369
rect 3054 20295 3110 20304
rect 4080 20262 4108 20946
rect 4250 20904 4306 20913
rect 4250 20839 4306 20848
rect 4264 20602 4292 20839
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 4068 20256 4120 20262
rect 4120 20216 4200 20244
rect 4068 20198 4120 20204
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2332 19417 2360 19654
rect 2318 19408 2374 19417
rect 2318 19343 2374 19352
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1780 18222 1808 18702
rect 2240 18465 2268 18906
rect 2226 18456 2282 18465
rect 2226 18391 2282 18400
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1412 15706 1440 18158
rect 1768 18080 1820 18086
rect 1582 18048 1638 18057
rect 1768 18022 1820 18028
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 1582 17983 1638 17992
rect 1490 16280 1546 16289
rect 1596 16250 1624 17983
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17202 1716 17478
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1688 17105 1716 17138
rect 1674 17096 1730 17105
rect 1674 17031 1730 17040
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1490 16215 1546 16224
rect 1584 16244 1636 16250
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1398 15328 1454 15337
rect 1398 15263 1454 15272
rect 1412 14618 1440 15263
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1504 11898 1532 16215
rect 1584 16186 1636 16192
rect 1688 15638 1716 16934
rect 1780 16697 1808 18022
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1766 16688 1822 16697
rect 1766 16623 1822 16632
rect 1780 16046 1808 16623
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1872 15706 1900 17478
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1964 16658 1992 16934
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1676 15632 1728 15638
rect 1872 15609 1900 15642
rect 1676 15574 1728 15580
rect 1858 15600 1914 15609
rect 1688 15065 1716 15574
rect 1858 15535 1914 15544
rect 1674 15056 1730 15065
rect 1674 14991 1730 15000
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11286 1440 11630
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1596 11218 1624 13330
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9722 1440 9998
rect 1688 9874 1716 14554
rect 1780 13190 1808 14894
rect 1858 14784 1914 14793
rect 1858 14719 1914 14728
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1872 12986 1900 14719
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1964 12481 1992 16594
rect 2056 15162 2084 17682
rect 2332 17678 2360 18022
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2136 17604 2188 17610
rect 2136 17546 2188 17552
rect 2148 17202 2176 17546
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2148 16998 2176 17138
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2148 16658 2176 16934
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2148 14550 2176 16594
rect 2226 14920 2282 14929
rect 2226 14855 2282 14864
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 14006 2084 14350
rect 2044 14000 2096 14006
rect 2044 13942 2096 13948
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2148 13394 2176 13806
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2148 12986 2176 13330
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2136 12640 2188 12646
rect 2134 12608 2136 12617
rect 2188 12608 2190 12617
rect 2134 12543 2190 12552
rect 1950 12472 2006 12481
rect 1950 12407 2006 12416
rect 1766 12336 1822 12345
rect 1766 12271 1768 12280
rect 1820 12271 1822 12280
rect 1768 12242 1820 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 11898 2084 12174
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2056 11336 2084 11834
rect 2056 11308 2176 11336
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2056 10470 2084 11154
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2056 9926 2084 10406
rect 2044 9920 2096 9926
rect 1688 9846 1808 9874
rect 2044 9862 2096 9868
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1032 8832 1084 8838
rect 1032 8774 1084 8780
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 480 244 2790
rect 662 1864 718 1873
rect 662 1799 718 1808
rect 676 480 704 1799
rect 1044 921 1072 8774
rect 1412 8498 1440 9658
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1688 9178 1716 9522
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1780 9110 1808 9846
rect 2056 9586 2084 9862
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1860 9376 1912 9382
rect 1858 9344 1860 9353
rect 1912 9344 1914 9353
rect 1858 9279 1914 9288
rect 2148 9178 2176 11308
rect 2240 9654 2268 14855
rect 2332 11898 2360 17614
rect 2424 16794 2452 20198
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19514 2820 19858
rect 2964 19712 3016 19718
rect 2962 19680 2964 19689
rect 3016 19680 3018 19689
rect 2962 19615 3018 19624
rect 3344 19514 3372 20198
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3436 19378 3464 19654
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2516 16969 2544 19110
rect 2608 17218 2636 19110
rect 2792 18834 2820 19178
rect 2962 19136 3018 19145
rect 2962 19071 3018 19080
rect 2976 18970 3004 19071
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2870 18592 2926 18601
rect 2700 17921 2728 18566
rect 2870 18527 2926 18536
rect 2884 18426 2912 18527
rect 3252 18426 3280 18770
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2686 17912 2742 17921
rect 2792 17882 2820 18158
rect 3804 17882 3832 19314
rect 3988 18902 4016 19314
rect 4080 19174 4108 19858
rect 4172 19242 4200 20216
rect 5552 20058 5580 21247
rect 6288 21078 6316 23287
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 8036 21350 8064 22034
rect 8116 22024 8168 22030
rect 8114 21992 8116 22001
rect 8168 21992 8170 22001
rect 8114 21927 8170 21936
rect 8024 21344 8076 21350
rect 8022 21312 8024 21321
rect 8076 21312 8078 21321
rect 8022 21247 8078 21256
rect 8758 21176 8814 21185
rect 8758 21111 8814 21120
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 20534 6040 20946
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 6012 20058 6040 20470
rect 7576 20466 7604 20742
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 6920 20324 6972 20330
rect 6920 20266 6972 20272
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5460 19802 5488 19858
rect 5460 19774 5580 19802
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4908 19394 4936 19654
rect 4724 19366 4936 19394
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4068 19168 4120 19174
rect 4436 19168 4488 19174
rect 4068 19110 4120 19116
rect 4434 19136 4436 19145
rect 4488 19136 4490 19145
rect 4434 19071 4490 19080
rect 3976 18896 4028 18902
rect 3976 18838 4028 18844
rect 4724 18834 4752 19366
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4816 19174 4844 19246
rect 4908 19174 4936 19366
rect 5552 19310 5580 19774
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 3896 18222 3924 18770
rect 4250 18456 4306 18465
rect 4250 18391 4306 18400
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 2686 17847 2742 17856
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 2608 17190 2728 17218
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2502 16960 2558 16969
rect 2502 16895 2558 16904
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2608 16046 2636 17070
rect 2700 16726 2728 17190
rect 3896 17134 3924 18158
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4080 17796 4108 18090
rect 4160 17808 4212 17814
rect 4080 17768 4160 17796
rect 4160 17750 4212 17756
rect 4066 17504 4122 17513
rect 4066 17439 4122 17448
rect 3884 17128 3936 17134
rect 3238 17096 3294 17105
rect 3056 17060 3108 17066
rect 3884 17070 3936 17076
rect 3238 17031 3294 17040
rect 3056 17002 3108 17008
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2688 16584 2740 16590
rect 2792 16561 2820 16594
rect 3068 16590 3096 17002
rect 3056 16584 3108 16590
rect 2688 16526 2740 16532
rect 2778 16552 2834 16561
rect 2700 16250 2728 16526
rect 3056 16526 3108 16532
rect 2778 16487 2834 16496
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2596 16040 2648 16046
rect 2502 16008 2558 16017
rect 2596 15982 2648 15988
rect 2502 15943 2558 15952
rect 2688 15972 2740 15978
rect 2412 15904 2464 15910
rect 2410 15872 2412 15881
rect 2464 15872 2466 15881
rect 2410 15807 2466 15816
rect 2516 15042 2544 15943
rect 2688 15914 2740 15920
rect 2700 15434 2728 15914
rect 2792 15881 2820 16487
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 15042 2820 15302
rect 2424 15014 2544 15042
rect 2608 15026 2820 15042
rect 2596 15020 2820 15026
rect 2424 14890 2452 15014
rect 2648 15014 2820 15020
rect 2596 14962 2648 14968
rect 2412 14884 2464 14890
rect 2412 14826 2464 14832
rect 2424 14618 2452 14826
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 13977 2452 14214
rect 2410 13968 2466 13977
rect 2410 13903 2466 13912
rect 2608 13462 2636 14962
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2700 13870 2728 14486
rect 2884 14113 2912 14554
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 2870 14104 2926 14113
rect 2870 14039 2872 14048
rect 2924 14039 2926 14048
rect 2872 14010 2924 14016
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2700 13734 2728 13806
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2884 13530 2912 13806
rect 3068 13734 3096 14350
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 13274 2820 13330
rect 2700 13246 2820 13274
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2516 10130 2544 10610
rect 2608 10554 2636 13126
rect 2700 12442 2728 13246
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2884 12374 2912 12854
rect 2962 12472 3018 12481
rect 2962 12407 2964 12416
rect 3016 12407 3018 12416
rect 2964 12378 3016 12384
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2608 10526 2728 10554
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9722 2544 10066
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2608 9518 2636 10406
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 1768 9104 1820 9110
rect 1768 9046 1820 9052
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1308 8356 1360 8362
rect 1308 8298 1360 8304
rect 1124 5840 1176 5846
rect 1124 5782 1176 5788
rect 1030 912 1086 921
rect 1030 847 1086 856
rect 202 0 258 480
rect 662 0 718 480
rect 1136 377 1164 5782
rect 1216 2916 1268 2922
rect 1216 2858 1268 2864
rect 1228 480 1256 2858
rect 1320 1465 1348 8298
rect 1412 7954 1440 8434
rect 1780 8294 1808 9046
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 2056 8362 2084 8842
rect 2148 8362 2176 9114
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1768 8288 1820 8294
rect 2240 8242 2268 9318
rect 2608 9217 2636 9454
rect 2594 9208 2650 9217
rect 2594 9143 2650 9152
rect 2502 8936 2558 8945
rect 2700 8906 2728 10526
rect 2792 10198 2820 12242
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11558 2912 12038
rect 2962 11792 3018 11801
rect 3068 11762 3096 13398
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 12102 3188 12650
rect 3252 12481 3280 17031
rect 3792 16720 3844 16726
rect 3790 16688 3792 16697
rect 3844 16688 3846 16697
rect 3516 16652 3568 16658
rect 3790 16623 3846 16632
rect 3516 16594 3568 16600
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3436 14006 3464 15438
rect 3528 15162 3556 16594
rect 3974 16008 4030 16017
rect 3974 15943 4030 15952
rect 3884 15496 3936 15502
rect 3882 15464 3884 15473
rect 3936 15464 3938 15473
rect 3882 15399 3938 15408
rect 3988 15201 4016 15943
rect 3974 15192 4030 15201
rect 3516 15156 3568 15162
rect 3974 15127 4030 15136
rect 3516 15098 3568 15104
rect 3790 14648 3846 14657
rect 4080 14618 4108 17439
rect 4264 16794 4292 18391
rect 4434 17912 4490 17921
rect 4434 17847 4490 17856
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4356 16697 4384 17614
rect 4342 16688 4398 16697
rect 4342 16623 4344 16632
rect 4396 16623 4398 16632
rect 4344 16594 4396 16600
rect 4158 15600 4214 15609
rect 4158 15535 4214 15544
rect 3790 14583 3846 14592
rect 4068 14612 4120 14618
rect 3424 14000 3476 14006
rect 3476 13960 3556 13988
rect 3424 13942 3476 13948
rect 3330 12880 3386 12889
rect 3330 12815 3386 12824
rect 3238 12472 3294 12481
rect 3238 12407 3294 12416
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 2962 11727 3018 11736
rect 3056 11756 3108 11762
rect 2976 11626 3004 11727
rect 3056 11698 3108 11704
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 11082 2912 11494
rect 3068 11354 3096 11698
rect 3238 11656 3294 11665
rect 3238 11591 3294 11600
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2502 8871 2558 8880
rect 2688 8900 2740 8906
rect 1768 8230 1820 8236
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1398 7440 1454 7449
rect 1398 7375 1400 7384
rect 1452 7375 1454 7384
rect 1400 7346 1452 7352
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 5778 1440 6054
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 3058 1440 5714
rect 1492 5092 1544 5098
rect 1492 5034 1544 5040
rect 1504 4690 1532 5034
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1596 2553 1624 8230
rect 2148 8214 2268 8242
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1688 7585 1716 7890
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1688 7002 1716 7511
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 6322 2084 6598
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1950 6216 2006 6225
rect 1688 5914 1716 6190
rect 1950 6151 2006 6160
rect 1964 6118 1992 6151
rect 1952 6112 2004 6118
rect 1858 6080 1914 6089
rect 1952 6054 2004 6060
rect 1858 6015 1914 6024
rect 1872 5914 1900 6015
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1872 5370 1900 5850
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1964 5098 1992 5510
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1964 4978 1992 5034
rect 1872 4950 1992 4978
rect 1872 4486 1900 4950
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1688 3369 1716 3878
rect 1674 3360 1730 3369
rect 1674 3295 1730 3304
rect 1688 2582 1716 3295
rect 1872 2825 1900 4422
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2056 3602 2084 3878
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1858 2816 1914 2825
rect 1858 2751 1914 2760
rect 1676 2576 1728 2582
rect 1582 2544 1638 2553
rect 1676 2518 1728 2524
rect 1582 2479 1638 2488
rect 2148 2009 2176 8214
rect 2410 8120 2466 8129
rect 2410 8055 2466 8064
rect 2318 6896 2374 6905
rect 2318 6831 2374 6840
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2240 4146 2268 4626
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2240 2650 2268 4082
rect 2332 4078 2360 6831
rect 2424 6730 2452 8055
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2516 5001 2544 8871
rect 2688 8842 2740 8848
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 2608 7342 2636 8298
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2700 8072 2728 8230
rect 2780 8084 2832 8090
rect 2700 8044 2780 8072
rect 2780 8026 2832 8032
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2688 6860 2740 6866
rect 2884 6848 2912 11018
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2976 10266 3004 10406
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 3146 9752 3202 9761
rect 3146 9687 3202 9696
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3068 7342 3096 9046
rect 3056 7336 3108 7342
rect 2740 6820 2912 6848
rect 2976 7296 3056 7324
rect 2688 6802 2740 6808
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2502 4992 2558 5001
rect 2502 4927 2558 4936
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2332 3670 2360 4014
rect 2410 3768 2466 3777
rect 2410 3703 2412 3712
rect 2464 3703 2466 3712
rect 2412 3674 2464 3680
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2134 2000 2190 2009
rect 2134 1935 2190 1944
rect 1766 1728 1822 1737
rect 1766 1663 1822 1672
rect 1306 1456 1362 1465
rect 1306 1391 1362 1400
rect 1780 480 1808 1663
rect 2332 480 2360 3606
rect 2424 2854 2452 3674
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2516 2650 2544 3402
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2608 2378 2636 6054
rect 2700 5846 2728 6802
rect 2976 6798 3004 7296
rect 3056 7278 3108 7284
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2976 6458 3004 6734
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2792 5370 2820 6258
rect 3068 6118 3096 6802
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2792 4282 2820 5306
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 2976 4321 3004 5238
rect 2962 4312 3018 4321
rect 2780 4276 2832 4282
rect 2962 4247 3018 4256
rect 2780 4218 2832 4224
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2686 3904 2742 3913
rect 2686 3839 2742 3848
rect 2700 3670 2728 3839
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2700 2922 2728 3606
rect 2976 3534 3004 4082
rect 3068 4049 3096 6054
rect 3160 5302 3188 9687
rect 3252 8838 3280 11591
rect 3344 9897 3372 12815
rect 3528 12782 3556 13960
rect 3606 13832 3662 13841
rect 3606 13767 3662 13776
rect 3516 12776 3568 12782
rect 3436 12724 3516 12730
rect 3436 12718 3568 12724
rect 3436 12702 3556 12718
rect 3436 12442 3464 12702
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3422 12200 3478 12209
rect 3422 12135 3478 12144
rect 3330 9888 3386 9897
rect 3330 9823 3386 9832
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3160 4486 3188 4966
rect 3344 4593 3372 7754
rect 3436 7313 3464 12135
rect 3620 11665 3648 13767
rect 3804 12753 3832 14583
rect 4068 14554 4120 14560
rect 4066 14512 4122 14521
rect 4172 14482 4200 15535
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4264 15026 4292 15370
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4066 14447 4068 14456
rect 4120 14447 4122 14456
rect 4160 14476 4212 14482
rect 4068 14418 4120 14424
rect 4160 14418 4212 14424
rect 4448 14006 4476 17847
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4632 17338 4660 17614
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4540 15910 4568 16594
rect 4816 16153 4844 19110
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 5184 18086 5212 18838
rect 6196 18834 6224 20198
rect 6932 19378 6960 20266
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7010 19408 7066 19417
rect 6920 19372 6972 19378
rect 7010 19343 7066 19352
rect 6920 19314 6972 19320
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5184 17882 5212 18022
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 16998 5212 17682
rect 5828 17678 5856 18022
rect 6104 17814 6132 18566
rect 6196 18426 6224 18770
rect 6748 18630 6776 19110
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6932 18630 6960 18838
rect 6736 18624 6788 18630
rect 6920 18624 6972 18630
rect 6736 18566 6788 18572
rect 6840 18584 6920 18612
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5172 16992 5224 16998
rect 4986 16960 5042 16969
rect 4986 16895 5042 16904
rect 5170 16960 5172 16969
rect 5224 16960 5226 16969
rect 5170 16895 5226 16904
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4802 16144 4858 16153
rect 4802 16079 4858 16088
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4436 13728 4488 13734
rect 4540 13705 4568 15846
rect 4710 15600 4766 15609
rect 4710 15535 4766 15544
rect 4724 15502 4752 15535
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4632 14618 4660 14962
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4724 14414 4752 15438
rect 4816 15337 4844 15846
rect 4908 15473 4936 16662
rect 5000 16250 5028 16895
rect 5460 16794 5488 17478
rect 5552 17134 5580 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6104 17338 6132 17750
rect 6748 17542 6776 18566
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5184 15586 5212 16526
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5000 15570 5212 15586
rect 4988 15564 5212 15570
rect 5040 15558 5212 15564
rect 4988 15506 5040 15512
rect 4894 15464 4950 15473
rect 4894 15399 4950 15408
rect 4802 15328 4858 15337
rect 4802 15263 4858 15272
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 14793 4844 14826
rect 4802 14784 4858 14793
rect 4802 14719 4858 14728
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4436 13670 4488 13676
rect 4526 13696 4582 13705
rect 3882 13424 3938 13433
rect 3882 13359 3938 13368
rect 3790 12744 3846 12753
rect 3790 12679 3846 12688
rect 3790 12472 3846 12481
rect 3790 12407 3846 12416
rect 3606 11656 3662 11665
rect 3606 11591 3662 11600
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 8974 3556 10406
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3516 8968 3568 8974
rect 3514 8936 3516 8945
rect 3568 8936 3570 8945
rect 3514 8871 3570 8880
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3422 7304 3478 7313
rect 3422 7239 3478 7248
rect 3528 6769 3556 8774
rect 3620 8634 3648 9386
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3514 6760 3570 6769
rect 3514 6695 3570 6704
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6254 3464 6598
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3606 4856 3662 4865
rect 3606 4791 3662 4800
rect 3330 4584 3386 4593
rect 3330 4519 3386 4528
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 4078 3188 4422
rect 3148 4072 3200 4078
rect 3054 4040 3110 4049
rect 3148 4014 3200 4020
rect 3054 3975 3110 3984
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 3054 3496 3110 3505
rect 3054 3431 3110 3440
rect 3068 2922 3096 3431
rect 3160 2990 3188 4014
rect 3344 3584 3372 4519
rect 3620 4185 3648 4791
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3424 3596 3476 3602
rect 3344 3556 3424 3584
rect 3424 3538 3476 3544
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 2686 2816 2742 2825
rect 2686 2751 2742 2760
rect 2870 2816 2926 2825
rect 2870 2751 2926 2760
rect 2700 2446 2728 2751
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2884 480 2912 2751
rect 3068 2650 3096 2858
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3436 480 3464 3538
rect 3712 3233 3740 8463
rect 3804 8401 3832 12407
rect 3896 10169 3924 13359
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12345 4016 13126
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 3974 12336 4030 12345
rect 3974 12271 4030 12280
rect 3988 11393 4016 12271
rect 4080 11762 4108 12922
rect 4448 12628 4476 13670
rect 4526 13631 4582 13640
rect 4528 12640 4580 12646
rect 4448 12600 4528 12628
rect 4528 12582 4580 12588
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4172 11558 4200 12242
rect 4342 12200 4398 12209
rect 4342 12135 4344 12144
rect 4396 12135 4398 12144
rect 4344 12106 4396 12112
rect 4540 11626 4568 12582
rect 4802 12336 4858 12345
rect 4802 12271 4804 12280
rect 4856 12271 4858 12280
rect 4804 12242 4856 12248
rect 4528 11620 4580 11626
rect 4528 11562 4580 11568
rect 4160 11552 4212 11558
rect 4158 11520 4160 11529
rect 4212 11520 4214 11529
rect 4158 11455 4214 11464
rect 3974 11384 4030 11393
rect 4540 11354 4568 11562
rect 3974 11319 4030 11328
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4158 11248 4214 11257
rect 4158 11183 4160 11192
rect 4212 11183 4214 11192
rect 4160 11154 4212 11160
rect 4172 11098 4200 11154
rect 3988 11070 4200 11098
rect 3882 10160 3938 10169
rect 3988 10130 4016 11070
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 3882 10095 3938 10104
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3974 10024 4030 10033
rect 3974 9959 4030 9968
rect 3882 9480 3938 9489
rect 3882 9415 3938 9424
rect 3790 8392 3846 8401
rect 3790 8327 3846 8336
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3804 7002 3832 7958
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3804 5914 3832 6938
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3896 5681 3924 9415
rect 3988 9081 4016 9959
rect 4172 9194 4200 10066
rect 4264 9353 4292 10406
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4250 9344 4306 9353
rect 4250 9279 4306 9288
rect 4080 9178 4200 9194
rect 4068 9172 4200 9178
rect 4120 9166 4200 9172
rect 4068 9114 4120 9120
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3974 8392 4030 8401
rect 4264 8344 4292 9279
rect 4356 8838 4384 9998
rect 4540 9722 4568 10610
rect 4908 10305 4936 14894
rect 5000 14822 5028 15506
rect 5276 14822 5304 15846
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5368 15026 5396 15302
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5448 14952 5500 14958
rect 5446 14920 5448 14929
rect 5500 14920 5502 14929
rect 5446 14855 5502 14864
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5264 14816 5316 14822
rect 5552 14804 5580 17070
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5828 16833 5856 16934
rect 5814 16824 5870 16833
rect 5814 16759 5870 16768
rect 6104 16726 6132 17274
rect 6840 16794 6868 18584
rect 6920 18566 6972 18572
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6092 16720 6144 16726
rect 6932 16674 6960 18022
rect 6092 16662 6144 16668
rect 6564 16658 6960 16674
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6552 16652 6960 16658
rect 6604 16646 6960 16652
rect 6552 16594 6604 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16114 6040 16594
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5264 14758 5316 14764
rect 5368 14776 5580 14804
rect 5000 14618 5028 14758
rect 5276 14657 5304 14758
rect 5262 14648 5318 14657
rect 4988 14612 5040 14618
rect 5262 14583 5318 14592
rect 4988 14554 5040 14560
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4986 13968 5042 13977
rect 4986 13903 5042 13912
rect 5000 13802 5028 13903
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5092 12918 5120 14282
rect 5184 13394 5212 14350
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5276 13462 5304 13670
rect 5264 13456 5316 13462
rect 5262 13424 5264 13433
rect 5316 13424 5318 13433
rect 5172 13388 5224 13394
rect 5262 13359 5318 13368
rect 5172 13330 5224 13336
rect 5368 13326 5396 14776
rect 5736 14521 5764 14826
rect 5722 14512 5778 14521
rect 5540 14476 5592 14482
rect 5722 14447 5778 14456
rect 5540 14418 5592 14424
rect 5552 13988 5580 14418
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5552 13960 5672 13988
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5092 11558 5120 12174
rect 5368 11762 5396 12242
rect 5460 11898 5488 13806
rect 5644 13716 5672 13960
rect 5724 13728 5776 13734
rect 5644 13688 5724 13716
rect 5724 13670 5776 13676
rect 5736 13530 5764 13670
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 6012 13394 6040 16050
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5552 12306 5580 12922
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5828 12442 5856 12718
rect 6012 12714 6040 13330
rect 6104 12986 6132 16390
rect 6564 15910 6592 16594
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6826 16552 6882 16561
rect 6656 15978 6684 16526
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6552 15904 6604 15910
rect 6550 15872 6552 15881
rect 6604 15872 6606 15881
rect 6550 15807 6606 15816
rect 6748 15706 6776 16526
rect 6826 16487 6882 16496
rect 6840 16114 6868 16487
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6552 15088 6604 15094
rect 6550 15056 6552 15065
rect 6604 15056 6606 15065
rect 6550 14991 6606 15000
rect 6550 14240 6606 14249
rect 6550 14175 6606 14184
rect 6182 13968 6238 13977
rect 6182 13903 6238 13912
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5998 12608 6054 12617
rect 5998 12543 6054 12552
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 10577 5120 11494
rect 5368 11218 5396 11698
rect 5460 11268 5488 11834
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5540 11280 5592 11286
rect 5460 11240 5540 11268
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 10606 5304 10950
rect 5460 10810 5488 11240
rect 5540 11222 5592 11228
rect 5828 11121 5856 11290
rect 5814 11112 5870 11121
rect 5814 11047 5870 11056
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5264 10600 5316 10606
rect 5078 10568 5134 10577
rect 5264 10542 5316 10548
rect 5078 10503 5134 10512
rect 4894 10296 4950 10305
rect 5276 10266 5304 10542
rect 4894 10231 4950 10240
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4632 8838 4660 10134
rect 5644 10130 5672 10678
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5644 10010 5672 10066
rect 5552 9982 5672 10010
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 9042 4936 9454
rect 4986 9208 5042 9217
rect 4986 9143 4988 9152
rect 5040 9143 5042 9152
rect 4988 9114 5040 9120
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 3974 8327 4030 8336
rect 3882 5672 3938 5681
rect 3882 5607 3938 5616
rect 3988 3641 4016 8327
rect 4080 8316 4292 8344
rect 4080 8090 4108 8316
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4158 7576 4214 7585
rect 4356 7562 4384 8774
rect 4632 8129 4660 8774
rect 4908 8566 4936 8978
rect 5368 8634 5396 9590
rect 5552 9110 5580 9982
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5630 9616 5686 9625
rect 5630 9551 5632 9560
rect 5684 9551 5686 9560
rect 5632 9522 5684 9528
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5644 8922 5672 9318
rect 5552 8894 5672 8922
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4896 8560 4948 8566
rect 4816 8508 4896 8514
rect 5552 8537 5580 8894
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 4816 8502 4948 8508
rect 5538 8528 5594 8537
rect 4816 8486 4936 8502
rect 4988 8492 5040 8498
rect 4618 8120 4674 8129
rect 4816 8090 4844 8486
rect 5538 8463 5594 8472
rect 4988 8434 5040 8440
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4618 8055 4674 8064
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4908 7750 4936 8366
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4214 7534 4384 7562
rect 4158 7511 4160 7520
rect 4212 7511 4214 7520
rect 4160 7482 4212 7488
rect 4908 7002 4936 7686
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4620 6656 4672 6662
rect 4250 6624 4306 6633
rect 4620 6598 4672 6604
rect 4250 6559 4306 6568
rect 4264 6254 4292 6559
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4632 6304 4660 6598
rect 4712 6316 4764 6322
rect 4632 6276 4712 6304
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 5914 4292 6190
rect 4356 6118 4384 6258
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4068 5908 4120 5914
rect 4252 5908 4304 5914
rect 4120 5868 4200 5896
rect 4068 5850 4120 5856
rect 4172 4690 4200 5868
rect 4252 5850 4304 5856
rect 4356 4758 4384 6054
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4356 4570 4384 4694
rect 4172 4542 4384 4570
rect 3974 3632 4030 3641
rect 3974 3567 4030 3576
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3698 3224 3754 3233
rect 3988 3194 4016 3334
rect 3698 3159 3754 3168
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4172 2666 4200 4542
rect 4526 4040 4582 4049
rect 4526 3975 4582 3984
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4252 3392 4304 3398
rect 4250 3360 4252 3369
rect 4304 3360 4306 3369
rect 4250 3295 4306 3304
rect 4448 3194 4476 3470
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 3988 2638 4200 2666
rect 3988 480 4016 2638
rect 4356 2514 4384 2926
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4540 480 4568 3975
rect 4632 3942 4660 6276
rect 4712 6258 4764 6264
rect 5000 5234 5028 8434
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7954 5212 8230
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7546 5212 7890
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5184 5370 5212 7346
rect 5276 6905 5304 8298
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 7410 5396 7958
rect 5460 7818 5488 8230
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5448 7200 5500 7206
rect 5354 7168 5410 7177
rect 5448 7142 5500 7148
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5354 7103 5410 7112
rect 5262 6896 5318 6905
rect 5262 6831 5318 6840
rect 5368 6798 5396 7103
rect 5460 6934 5488 7142
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 5710 5304 6598
rect 5368 6458 5396 6734
rect 5460 6458 5488 6870
rect 5552 6798 5580 7142
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5078 5128 5134 5137
rect 5078 5063 5134 5072
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 2689 4660 3878
rect 5000 3777 5028 4966
rect 4986 3768 5042 3777
rect 4986 3703 5042 3712
rect 4618 2680 4674 2689
rect 4618 2615 4674 2624
rect 4632 2582 4660 2615
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 5092 480 5120 5063
rect 5276 4486 5304 5646
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5030 5396 5510
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 4146 5304 4422
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 3602 5304 4082
rect 5368 3913 5396 4966
rect 5460 4060 5488 6122
rect 5552 5778 5580 6734
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5234 6040 12543
rect 6090 11792 6146 11801
rect 6090 11727 6146 11736
rect 6104 10554 6132 11727
rect 6196 10674 6224 13903
rect 6564 13870 6592 14175
rect 6932 13870 6960 15302
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6288 11898 6316 12310
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6288 11354 6316 11834
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6380 11098 6408 13398
rect 6472 12782 6500 13670
rect 6564 12986 6592 13806
rect 6828 13728 6880 13734
rect 6826 13696 6828 13705
rect 6880 13696 6882 13705
rect 6826 13631 6882 13640
rect 7024 12986 7052 19343
rect 7116 19174 7144 19790
rect 7392 19174 7420 19858
rect 7104 19168 7156 19174
rect 7380 19168 7432 19174
rect 7104 19110 7156 19116
rect 7194 19136 7250 19145
rect 7380 19110 7432 19116
rect 7194 19071 7250 19080
rect 7208 18970 7236 19071
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7484 18426 7512 20198
rect 7576 20058 7604 20402
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8128 19514 8156 19994
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8312 19310 8340 19654
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7760 17882 7788 18702
rect 8312 18630 8340 19246
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8024 18080 8076 18086
rect 8022 18048 8024 18057
rect 8076 18048 8078 18057
rect 8022 17983 8078 17992
rect 8312 17898 8340 18566
rect 8680 18465 8708 19110
rect 8666 18456 8722 18465
rect 8666 18391 8668 18400
rect 8720 18391 8722 18400
rect 8668 18362 8720 18368
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 8220 17870 8340 17898
rect 7300 17134 7328 17818
rect 8220 17542 8248 17870
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7288 16992 7340 16998
rect 7392 16946 7420 17478
rect 7340 16940 7420 16946
rect 7288 16934 7420 16940
rect 7300 16918 7420 16934
rect 7300 16454 7328 16918
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7102 15056 7158 15065
rect 7102 14991 7104 15000
rect 7156 14991 7158 15000
rect 7104 14962 7156 14968
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6840 12424 6868 12650
rect 6920 12436 6972 12442
rect 6840 12396 6920 12424
rect 6920 12378 6972 12384
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11558 6592 12038
rect 6552 11552 6604 11558
rect 7104 11552 7156 11558
rect 6552 11494 6604 11500
rect 6918 11520 6974 11529
rect 6380 11070 6500 11098
rect 6366 10976 6422 10985
rect 6366 10911 6422 10920
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6104 10526 6224 10554
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6104 9450 6132 10066
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6104 7206 6132 7822
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5552 4690 5580 5170
rect 6196 4826 6224 10526
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6288 9586 6316 10202
rect 6380 10010 6408 10911
rect 6472 10130 6500 11070
rect 6564 10810 6592 11494
rect 7104 11494 7156 11500
rect 6918 11455 6974 11464
rect 6826 11384 6882 11393
rect 6826 11319 6882 11328
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6564 10554 6592 10746
rect 6564 10526 6776 10554
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6642 10432 6698 10441
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6380 9982 6500 10010
rect 6564 9994 6592 10406
rect 6642 10367 6698 10376
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 8634 6316 8978
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6472 6168 6500 9982
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6564 9722 6592 9930
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6550 8392 6606 8401
rect 6550 8327 6552 8336
rect 6604 8327 6606 8336
rect 6552 8298 6604 8304
rect 6656 7585 6684 10367
rect 6748 9586 6776 10526
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6840 8566 6868 11319
rect 6932 10674 6960 11455
rect 7116 11354 7144 11494
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 7102 10568 7158 10577
rect 7102 10503 7158 10512
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9518 6960 10066
rect 7116 9926 7144 10503
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9518 7144 9862
rect 6920 9512 6972 9518
rect 7104 9512 7156 9518
rect 6920 9454 6972 9460
rect 7102 9480 7104 9489
rect 7156 9480 7158 9489
rect 7102 9415 7158 9424
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7750 6960 8230
rect 6736 7744 6788 7750
rect 6920 7744 6972 7750
rect 6788 7704 6868 7732
rect 6736 7686 6788 7692
rect 6642 7576 6698 7585
rect 6642 7511 6698 7520
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6380 6140 6500 6168
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 5030 6316 5714
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4826 6316 4966
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 4214 5580 4626
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5540 4072 5592 4078
rect 5460 4032 5540 4060
rect 5540 4014 5592 4020
rect 5540 3936 5592 3942
rect 5354 3904 5410 3913
rect 5540 3878 5592 3884
rect 5354 3839 5410 3848
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5172 3120 5224 3126
rect 5170 3088 5172 3097
rect 5224 3088 5226 3097
rect 5170 3023 5226 3032
rect 5552 2990 5580 3878
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5736 2922 5764 2994
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 6012 2802 6040 4762
rect 6380 4706 6408 6140
rect 6458 6080 6514 6089
rect 6458 6015 6514 6024
rect 6472 5166 6500 6015
rect 6656 5370 6684 6802
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 6254 6776 6666
rect 6840 6440 6868 7704
rect 6920 7686 6972 7692
rect 6932 7449 6960 7686
rect 7024 7478 7052 8434
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7012 7472 7064 7478
rect 6918 7440 6974 7449
rect 7012 7414 7064 7420
rect 6918 7375 6974 7384
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 6866 6960 7278
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6840 6412 6960 6440
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6840 5914 6868 6258
rect 6932 6186 6960 6412
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 5736 2774 6040 2802
rect 6196 4678 6408 4706
rect 5736 2292 5764 2774
rect 5552 2264 5764 2292
rect 5552 1986 5580 2264
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5552 1958 5672 1986
rect 5644 480 5672 1958
rect 6196 480 6224 4678
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6288 2922 6316 3538
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 2990 6500 3402
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6288 2650 6316 2858
rect 6564 2854 6592 4014
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3398 6776 3878
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3058 6776 3334
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6656 1873 6684 2450
rect 6642 1864 6698 1873
rect 6642 1799 6698 1808
rect 6840 610 6868 5170
rect 7116 5137 7144 8298
rect 7208 8090 7236 15914
rect 7300 15609 7328 16390
rect 7576 16250 7604 16730
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7470 16144 7526 16153
rect 7470 16079 7526 16088
rect 7484 15706 7512 16079
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7286 15600 7342 15609
rect 7286 15535 7342 15544
rect 7300 15434 7328 15535
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7300 14006 7328 14418
rect 7380 14408 7432 14414
rect 7576 14396 7604 16186
rect 7944 15706 7972 16390
rect 8036 15910 8064 16526
rect 8116 16040 8168 16046
rect 8220 16028 8248 17478
rect 8168 16000 8248 16028
rect 8116 15982 8168 15988
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7668 15162 7696 15574
rect 7746 15464 7802 15473
rect 7746 15399 7802 15408
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7576 14368 7696 14396
rect 7380 14350 7432 14356
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7300 10606 7328 13942
rect 7392 13870 7420 14350
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 10198 7328 10406
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7206 7236 7822
rect 7392 7562 7420 13806
rect 7668 13462 7696 14368
rect 7760 14346 7788 15399
rect 7944 14618 7972 15642
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7852 13530 7880 14282
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12782 7512 13126
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 11082 7512 12718
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7576 11286 7604 12378
rect 7852 11762 7880 13194
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12345 7972 13126
rect 7930 12336 7986 12345
rect 7930 12271 7986 12280
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7576 10674 7604 11222
rect 7564 10668 7616 10674
rect 8036 10656 8064 15846
rect 8312 15722 8340 17614
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16726 8432 16934
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8220 15694 8340 15722
rect 8588 15706 8616 15982
rect 8576 15700 8628 15706
rect 8220 15638 8248 15694
rect 8576 15642 8628 15648
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8588 15502 8616 15642
rect 8116 15496 8168 15502
rect 8576 15496 8628 15502
rect 8116 15438 8168 15444
rect 8206 15464 8262 15473
rect 8128 15162 8156 15438
rect 8576 15438 8628 15444
rect 8206 15399 8208 15408
rect 8260 15399 8262 15408
rect 8208 15370 8260 15376
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8128 13938 8156 14894
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8772 13716 8800 21111
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 8942 17504 8998 17513
rect 8942 17439 8998 17448
rect 8850 16960 8906 16969
rect 8956 16946 8984 17439
rect 9048 16998 9076 17682
rect 8906 16918 8984 16946
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8850 16895 8906 16904
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 15366 8892 15846
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8864 14958 8892 15302
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8864 13870 8892 14554
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8772 13688 8892 13716
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8312 12918 8340 13330
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8128 11558 8156 12786
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 12186 8248 12582
rect 8312 12288 8340 12854
rect 8496 12442 8524 13262
rect 8588 12986 8616 13398
rect 8864 12986 8892 13688
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8758 12472 8814 12481
rect 8484 12436 8536 12442
rect 8758 12407 8814 12416
rect 8484 12378 8536 12384
rect 8312 12260 8524 12288
rect 8220 12158 8432 12186
rect 8404 12102 8432 12158
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11898 8432 12038
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8496 11778 8524 12260
rect 8404 11750 8524 11778
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8404 11354 8432 11750
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8036 10628 8156 10656
rect 7564 10610 7616 10616
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 8022 10568 8078 10577
rect 7760 10470 7788 10542
rect 8022 10503 8078 10512
rect 8036 10470 8064 10503
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7576 10130 7604 10406
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7760 10062 7788 10406
rect 7930 10296 7986 10305
rect 7930 10231 7986 10240
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7654 8936 7710 8945
rect 7654 8871 7656 8880
rect 7708 8871 7710 8880
rect 7656 8842 7708 8848
rect 7760 8838 7788 9998
rect 7944 9110 7972 10231
rect 8024 9648 8076 9654
rect 8022 9616 8024 9625
rect 8076 9616 8078 9625
rect 8022 9551 8078 9560
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7944 8362 7972 8910
rect 8036 8634 8064 9551
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 8128 8294 8156 10628
rect 8404 10266 8432 11290
rect 8496 11150 8524 11562
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10266 8616 10610
rect 8772 10538 8800 12407
rect 8864 10810 8892 12582
rect 8956 12481 8984 16918
rect 9048 15366 9076 16934
rect 9140 16794 9168 19110
rect 9232 18426 9260 23423
rect 10060 22658 10088 26318
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 21008 23866 21036 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 15290 23624 15346 23633
rect 15290 23559 15346 23568
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 9876 22630 10088 22658
rect 9678 21312 9734 21321
rect 9678 21247 9734 21256
rect 9692 21146 9720 21247
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9692 20602 9720 20946
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9508 19718 9536 20334
rect 9692 20058 9720 20538
rect 9772 20324 9824 20330
rect 9772 20266 9824 20272
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9784 19378 9812 20266
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9784 18970 9812 19314
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9692 18290 9720 18566
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9588 18080 9640 18086
rect 9640 18040 9720 18068
rect 9588 18022 9640 18028
rect 9692 17882 9720 18040
rect 9770 18048 9826 18057
rect 9770 17983 9826 17992
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9508 17202 9536 17478
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9126 16688 9182 16697
rect 9126 16623 9182 16632
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8942 12472 8998 12481
rect 8942 12407 8998 12416
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8220 8974 8248 9998
rect 9048 9926 9076 10474
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 9178 8340 9454
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8312 9058 8340 9114
rect 8312 9030 8524 9058
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7300 7534 7420 7562
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7102 5128 7158 5137
rect 7102 5063 7158 5072
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 2961 6960 4966
rect 6918 2952 6974 2961
rect 6918 2887 6974 2896
rect 7208 2446 7236 7142
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 6736 604 6788 610
rect 6736 546 6788 552
rect 6828 604 6880 610
rect 6828 546 6880 552
rect 6748 480 6776 546
rect 7300 480 7328 7534
rect 7484 6934 7512 7686
rect 7576 7002 7604 7890
rect 8128 7857 8156 7890
rect 8114 7848 8170 7857
rect 7656 7812 7708 7818
rect 8114 7783 8170 7792
rect 7656 7754 7708 7760
rect 7668 7342 7696 7754
rect 7748 7744 7800 7750
rect 7746 7712 7748 7721
rect 7800 7712 7802 7721
rect 7746 7647 7802 7656
rect 8128 7546 8156 7783
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 7392 8248 8774
rect 8312 8022 8340 8842
rect 8404 8022 8432 8910
rect 8496 8634 8524 9030
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8576 8560 8628 8566
rect 8574 8528 8576 8537
rect 8628 8528 8630 8537
rect 8574 8463 8630 8472
rect 8772 8362 8800 8774
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8128 7364 8248 7392
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7668 7002 7696 7278
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 6322 7420 6802
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7378 5672 7434 5681
rect 7378 5607 7434 5616
rect 7392 5370 7420 5607
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7576 4282 7604 6054
rect 7746 5264 7802 5273
rect 7746 5199 7802 5208
rect 7760 4758 7788 5199
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7470 2680 7526 2689
rect 7470 2615 7526 2624
rect 7484 2446 7512 2615
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7392 2281 7420 2382
rect 7378 2272 7434 2281
rect 7378 2207 7434 2216
rect 7576 2145 7604 2450
rect 7562 2136 7618 2145
rect 7562 2071 7618 2080
rect 7944 1873 7972 4966
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 3369 8064 4422
rect 8022 3360 8078 3369
rect 8022 3295 8078 3304
rect 7930 1864 7986 1873
rect 7930 1799 7986 1808
rect 8128 610 8156 7364
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8220 6304 8248 7210
rect 8300 6316 8352 6322
rect 8220 6276 8300 6304
rect 8352 6276 8432 6304
rect 8300 6258 8352 6264
rect 8404 5846 8432 6276
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8392 5840 8444 5846
rect 8588 5817 8616 6122
rect 8392 5782 8444 5788
rect 8574 5808 8630 5817
rect 8300 5772 8352 5778
rect 8574 5743 8630 5752
rect 8300 5714 8352 5720
rect 8312 5681 8340 5714
rect 8588 5710 8616 5743
rect 8392 5704 8444 5710
rect 8298 5672 8354 5681
rect 8392 5646 8444 5652
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8298 5607 8354 5616
rect 8208 5568 8260 5574
rect 8260 5516 8340 5522
rect 8208 5510 8340 5516
rect 8220 5494 8340 5510
rect 8312 5030 8340 5494
rect 8404 5166 8432 5646
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8482 5128 8538 5137
rect 8482 5063 8538 5072
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8220 3738 8248 4490
rect 8312 4049 8340 4966
rect 8496 4690 8524 5063
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4826 8616 4966
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4282 8432 4422
rect 8496 4282 8524 4626
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8298 4040 8354 4049
rect 8298 3975 8354 3984
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8404 2378 8432 3606
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8496 3194 8524 3470
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8680 2802 8708 8026
rect 8864 6866 8892 8366
rect 8956 8090 8984 8434
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8864 5914 8892 6802
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8772 4758 8800 5782
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 5030 8984 5170
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8772 3738 8800 4694
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8864 4593 8892 4626
rect 8850 4584 8906 4593
rect 8850 4519 8906 4528
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8772 2922 8800 3674
rect 8956 3505 8984 4966
rect 9048 3641 9076 9862
rect 9034 3632 9090 3641
rect 9034 3567 9090 3576
rect 8942 3496 8998 3505
rect 8942 3431 8998 3440
rect 8942 3088 8998 3097
rect 8942 3023 8998 3032
rect 8956 2990 8984 3023
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 9140 2854 9168 16623
rect 9496 16584 9548 16590
rect 9692 16538 9720 17274
rect 9496 16526 9548 16532
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9416 15910 9444 16390
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9508 15586 9536 16526
rect 9600 16510 9720 16538
rect 9600 16046 9628 16510
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9588 16040 9640 16046
rect 9692 16017 9720 16390
rect 9588 15982 9640 15988
rect 9678 16008 9734 16017
rect 9678 15943 9734 15952
rect 9508 15570 9720 15586
rect 9312 15564 9364 15570
rect 9508 15564 9732 15570
rect 9508 15558 9680 15564
rect 9312 15506 9364 15512
rect 9324 14278 9352 15506
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9312 14272 9364 14278
rect 9310 14240 9312 14249
rect 9364 14240 9366 14249
rect 9310 14175 9366 14184
rect 9416 13297 9444 15302
rect 9494 15192 9550 15201
rect 9494 15127 9496 15136
rect 9548 15127 9550 15136
rect 9496 15098 9548 15104
rect 9508 14618 9536 15098
rect 9600 14890 9628 15558
rect 9680 15506 9732 15512
rect 9784 15337 9812 17983
rect 9770 15328 9826 15337
rect 9770 15263 9826 15272
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9402 13288 9458 13297
rect 9402 13223 9458 13232
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12442 9260 12650
rect 9416 12646 9444 13126
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9508 12458 9536 13670
rect 9692 13530 9720 14214
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9416 12430 9536 12458
rect 9416 11762 9444 12430
rect 9588 12300 9640 12306
rect 9692 12288 9720 12786
rect 9640 12260 9720 12288
rect 9588 12242 9640 12248
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10470 9260 10950
rect 9508 10674 9536 11018
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9508 9450 9536 10066
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9178 9536 9386
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9600 9042 9628 11086
rect 9784 10606 9812 13126
rect 9876 11694 9904 22630
rect 9954 22536 10010 22545
rect 9954 22471 10010 22480
rect 9968 16708 9996 22471
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10046 22128 10102 22137
rect 10046 22063 10102 22072
rect 10060 17796 10088 22063
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11348 21049 11376 21082
rect 12348 21072 12400 21078
rect 11334 21040 11390 21049
rect 12348 21014 12400 21020
rect 11334 20975 11390 20984
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10152 20058 10180 20878
rect 10244 20398 10272 20878
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 11532 20398 11560 20810
rect 11992 20602 12020 20946
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 10232 20392 10284 20398
rect 11520 20392 11572 20398
rect 10232 20334 10284 20340
rect 11518 20360 11520 20369
rect 11572 20360 11574 20369
rect 11518 20295 11574 20304
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20198
rect 12176 20058 12204 20266
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 10152 19514 10180 19994
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10704 18766 10732 19790
rect 12176 19378 12204 19994
rect 12360 19514 12388 21014
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12452 20466 12480 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 13910 20496 13966 20505
rect 12440 20460 12492 20466
rect 13910 20431 13966 20440
rect 12440 20402 12492 20408
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12452 19496 12480 20402
rect 13818 20360 13874 20369
rect 13818 20295 13874 20304
rect 13832 20262 13860 20295
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 12532 19508 12584 19514
rect 12452 19468 12532 19496
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10060 17768 10640 17796
rect 10138 17096 10194 17105
rect 10138 17031 10194 17040
rect 10612 17048 10640 17768
rect 10704 17678 10732 18702
rect 10980 18086 11008 18770
rect 10968 18080 11020 18086
rect 11152 18080 11204 18086
rect 11020 18040 11100 18068
rect 10968 18022 11020 18028
rect 11072 17882 11100 18040
rect 11152 18022 11204 18028
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 11164 17542 11192 18022
rect 10784 17536 10836 17542
rect 10782 17504 10784 17513
rect 11152 17536 11204 17542
rect 10836 17504 10838 17513
rect 11152 17478 11204 17484
rect 10782 17439 10838 17448
rect 10784 17060 10836 17066
rect 10152 16794 10180 17031
rect 10612 17020 10732 17048
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16788 10192 16794
rect 10192 16748 10272 16776
rect 10140 16730 10192 16736
rect 9968 16680 10088 16708
rect 10060 16674 10088 16680
rect 10060 16646 10180 16674
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 15910 9996 16526
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 11354 9904 11494
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9784 9994 9812 10542
rect 9876 10538 9904 11290
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9716 9732 9722
rect 9784 9704 9812 9930
rect 9732 9676 9812 9704
rect 9680 9658 9732 9664
rect 9876 9518 9904 10134
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 4842 9260 8230
rect 9324 6866 9352 8978
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9416 7954 9444 8842
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9508 6458 9536 8026
rect 9600 7970 9628 8298
rect 9692 8090 9720 8570
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9600 7942 9720 7970
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9508 5370 9536 6394
rect 9692 5914 9720 7942
rect 9784 6633 9812 8774
rect 9876 7721 9904 8910
rect 9968 8480 9996 15846
rect 10152 15162 10180 16646
rect 10244 16182 10272 16748
rect 10704 16250 10732 17020
rect 10784 17002 10836 17008
rect 10796 16794 10824 17002
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10796 16114 10824 16730
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10980 15910 11008 16390
rect 10876 15904 10928 15910
rect 10968 15904 11020 15910
rect 10876 15846 10928 15852
rect 10966 15872 10968 15881
rect 11152 15904 11204 15910
rect 11020 15872 11022 15881
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10888 15706 10916 15846
rect 11152 15846 11204 15852
rect 10966 15807 11022 15816
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 11164 15638 11192 15846
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10152 14618 10180 14826
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10888 14414 10916 15506
rect 11164 15026 11192 15574
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11072 14550 11100 14758
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10876 14408 10928 14414
rect 10704 14368 10876 14396
rect 10704 14006 10732 14368
rect 10876 14350 10928 14356
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13326 10732 13942
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12646 10732 13262
rect 10796 12918 10824 13330
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12374 10732 12582
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11082 10088 12242
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10152 10198 10180 11630
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11354 10732 11698
rect 10888 11642 10916 13806
rect 10980 13802 11008 14418
rect 11072 14074 11100 14486
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11150 13288 11206 13297
rect 11150 13223 11206 13232
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10980 12424 11008 12854
rect 11164 12782 11192 13223
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11060 12436 11112 12442
rect 10980 12396 11060 12424
rect 11060 12378 11112 12384
rect 10888 11614 11008 11642
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10690 10432 10746 10441
rect 10289 10364 10585 10384
rect 10690 10367 10746 10376
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 10367
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10796 10062 10824 11154
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10324 10056 10376 10062
rect 10784 10056 10836 10062
rect 10324 9998 10376 10004
rect 10782 10024 10784 10033
rect 10836 10024 10838 10033
rect 10152 9382 10180 9998
rect 10336 9897 10364 9998
rect 10782 9959 10838 9968
rect 10322 9888 10378 9897
rect 10322 9823 10378 9832
rect 10690 9480 10746 9489
rect 10690 9415 10746 9424
rect 10704 9382 10732 9415
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10048 9036 10100 9042
rect 10152 9024 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10506 9072 10562 9081
rect 10152 8996 10272 9024
rect 10506 9007 10562 9016
rect 10048 8978 10100 8984
rect 10060 8634 10088 8978
rect 10138 8936 10194 8945
rect 10138 8871 10194 8880
rect 10152 8634 10180 8871
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10244 8566 10272 8996
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 9968 8452 10180 8480
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9862 7712 9918 7721
rect 9862 7647 9918 7656
rect 9876 6866 9904 7647
rect 9968 7274 9996 7822
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9968 6730 9996 7210
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9770 6624 9826 6633
rect 9770 6559 9826 6568
rect 9864 6112 9916 6118
rect 9862 6080 9864 6089
rect 9916 6080 9918 6089
rect 9862 6015 9918 6024
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9232 4814 9444 4842
rect 9128 2848 9180 2854
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8496 2258 8524 2790
rect 8680 2774 8984 2802
rect 9128 2790 9180 2796
rect 9218 2816 9274 2825
rect 8668 2440 8720 2446
rect 8666 2408 8668 2417
rect 8720 2408 8722 2417
rect 8666 2343 8722 2352
rect 8404 2230 8524 2258
rect 7840 604 7892 610
rect 7840 546 7892 552
rect 8116 604 8168 610
rect 8116 546 8168 552
rect 7852 480 7880 546
rect 8404 480 8432 2230
rect 8956 480 8984 2774
rect 9218 2751 9274 2760
rect 9232 2650 9260 2751
rect 9416 2666 9444 4814
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 4282 9536 4626
rect 9600 4593 9628 4966
rect 9680 4616 9732 4622
rect 9586 4584 9642 4593
rect 9680 4558 9732 4564
rect 9586 4519 9642 4528
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9588 3732 9640 3738
rect 9692 3720 9720 4558
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9876 4146 9904 4490
rect 10060 4214 10088 8230
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9640 3692 9720 3720
rect 9588 3674 9640 3680
rect 9220 2644 9272 2650
rect 9416 2638 9536 2666
rect 9220 2586 9272 2592
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9416 1737 9444 2246
rect 9402 1728 9458 1737
rect 9402 1663 9458 1672
rect 9508 480 9536 2638
rect 9600 2530 9628 3674
rect 9876 3670 9904 4082
rect 10152 4026 10180 8452
rect 10520 8430 10548 9007
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8910
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10704 7342 10732 8026
rect 10796 8022 10824 8298
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10888 7857 10916 11494
rect 10980 8401 11008 11614
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11072 11257 11100 11290
rect 11256 11286 11284 18022
rect 11348 13569 11376 19110
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 18086 11560 18226
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 17746 11560 18022
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11808 17105 11836 19110
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18465 12112 18566
rect 12070 18456 12126 18465
rect 12452 18426 12480 19468
rect 12532 19450 12584 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12636 18970 12664 19314
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12070 18391 12126 18400
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12452 17814 12480 18362
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12452 17202 12480 17750
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 11794 17096 11850 17105
rect 11794 17031 11850 17040
rect 12452 16726 12480 17138
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16794 12664 17002
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11900 16250 11928 16594
rect 12452 16250 12480 16662
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 11900 15706 11928 16186
rect 12438 15872 12494 15881
rect 12438 15807 12494 15816
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 12452 15162 12480 15807
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12622 15464 12678 15473
rect 12622 15399 12678 15408
rect 12530 15328 12586 15337
rect 12530 15263 12586 15272
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 11886 14920 11942 14929
rect 11886 14855 11888 14864
rect 11940 14855 11942 14864
rect 11888 14826 11940 14832
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11716 13938 11744 14418
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11716 13734 11744 13874
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11334 13560 11390 13569
rect 11716 13530 11744 13670
rect 11334 13495 11390 13504
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11440 12646 11468 13398
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12850 11928 13126
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11244 11280 11296 11286
rect 11058 11248 11114 11257
rect 11244 11222 11296 11228
rect 11058 11183 11114 11192
rect 11440 11150 11468 12582
rect 11900 12102 11928 12786
rect 12176 12356 12204 14758
rect 12452 14618 12480 14962
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12438 13424 12494 13433
rect 12438 13359 12494 13368
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12176 12328 12296 12356
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11808 11558 11836 11698
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11060 11008 11112 11014
rect 11808 10985 11836 11494
rect 11060 10950 11112 10956
rect 11794 10976 11850 10985
rect 11072 10810 11100 10950
rect 11794 10911 11850 10920
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11256 9722 11284 9930
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11256 9042 11284 9658
rect 11348 9178 11376 10066
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10966 8392 11022 8401
rect 10966 8327 11022 8336
rect 11060 8016 11112 8022
rect 10966 7984 11022 7993
rect 11060 7958 11112 7964
rect 10966 7919 11022 7928
rect 10874 7848 10930 7857
rect 10874 7783 10930 7792
rect 10692 7336 10744 7342
rect 10980 7290 11008 7919
rect 10692 7278 10744 7284
rect 10888 7262 11008 7290
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10888 6934 10916 7262
rect 11072 7206 11100 7958
rect 11060 7200 11112 7206
rect 10980 7148 11060 7154
rect 10980 7142 11112 7148
rect 10980 7126 11100 7142
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 6186 10456 6734
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 6361 10548 6598
rect 10612 6458 10640 6870
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10876 6724 10928 6730
rect 10980 6712 11008 7126
rect 10928 6684 11008 6712
rect 10876 6666 10928 6672
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10506 6352 10562 6361
rect 10506 6287 10562 6296
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10796 5710 10824 6666
rect 10888 5914 10916 6666
rect 11058 6216 11114 6225
rect 11058 6151 11114 6160
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10796 5098 10824 5646
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10796 4690 10824 5034
rect 11072 5001 11100 6151
rect 11164 5846 11192 8434
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 6934 11376 8298
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11440 6458 11468 10406
rect 11518 10160 11574 10169
rect 11518 10095 11574 10104
rect 11532 9382 11560 10095
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 11794 9752 11850 9761
rect 11794 9687 11850 9696
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11808 8634 11836 9687
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11808 8430 11836 8570
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11796 8424 11848 8430
rect 11702 8392 11758 8401
rect 11796 8366 11848 8372
rect 11702 8327 11758 8336
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11624 7002 11652 7890
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11518 6760 11574 6769
rect 11518 6695 11574 6704
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11334 6216 11390 6225
rect 11334 6151 11336 6160
rect 11388 6151 11390 6160
rect 11336 6122 11388 6128
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11164 5370 11192 5782
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11058 4992 11114 5001
rect 11058 4927 11114 4936
rect 10874 4856 10930 4865
rect 10874 4791 10930 4800
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10888 4282 10916 4791
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10060 3998 10180 4026
rect 10692 4072 10744 4078
rect 10980 4060 11008 4558
rect 10980 4032 11100 4060
rect 10692 4014 10744 4020
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9770 3496 9826 3505
rect 9770 3431 9826 3440
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 2650 9720 3334
rect 9784 3126 9812 3431
rect 9876 3194 9904 3606
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9678 2544 9734 2553
rect 9600 2502 9678 2530
rect 9678 2479 9734 2488
rect 9968 2310 9996 2586
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 10060 480 10088 3998
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3505 10180 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10138 3496 10194 3505
rect 10138 3431 10194 3440
rect 10152 2582 10180 3431
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2650 10732 4014
rect 11072 3942 11100 4032
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 3398 11100 3878
rect 11150 3632 11206 3641
rect 11150 3567 11206 3576
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 3097 11100 3334
rect 11058 3088 11114 3097
rect 11058 3023 11060 3032
rect 11112 3023 11114 3032
rect 11060 2994 11112 3000
rect 11072 2963 11100 2994
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10598 1048 10654 1057
rect 10598 983 10654 992
rect 10612 480 10640 983
rect 11164 480 11192 3567
rect 11256 3194 11284 5607
rect 11532 5409 11560 6695
rect 11518 5400 11574 5409
rect 11518 5335 11574 5344
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11336 3936 11388 3942
rect 11334 3904 11336 3913
rect 11388 3904 11390 3913
rect 11334 3839 11390 3848
rect 11624 3602 11652 4558
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11624 3466 11652 3538
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11256 2990 11284 3130
rect 11428 3120 11480 3126
rect 11426 3088 11428 3097
rect 11480 3088 11482 3097
rect 11426 3023 11482 3032
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11334 2680 11390 2689
rect 11334 2615 11336 2624
rect 11388 2615 11390 2624
rect 11336 2586 11388 2592
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1465 11652 2246
rect 11610 1456 11666 1465
rect 11610 1391 11666 1400
rect 11716 480 11744 8327
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 4690 11928 5510
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 3942 11928 4626
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3641 11928 3878
rect 11886 3632 11942 3641
rect 11886 3567 11942 3576
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11808 3369 11836 3470
rect 11794 3360 11850 3369
rect 11794 3295 11850 3304
rect 11808 3194 11836 3295
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11992 2038 12020 8502
rect 12084 2530 12112 9522
rect 12176 9518 12204 9862
rect 12268 9654 12296 12328
rect 12360 12238 12388 12582
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11937 12388 12038
rect 12346 11928 12402 11937
rect 12346 11863 12402 11872
rect 12452 11830 12480 13359
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12360 9659 12388 10746
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12346 9650 12402 9659
rect 12346 9585 12402 9594
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 7818 12388 9454
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12176 6866 12204 7346
rect 12452 6934 12480 7686
rect 12544 7478 12572 15263
rect 12636 12986 12664 15399
rect 13004 15026 13032 15642
rect 13818 15056 13874 15065
rect 12992 15020 13044 15026
rect 13818 14991 13820 15000
rect 12992 14962 13044 14968
rect 13872 14991 13874 15000
rect 13820 14962 13872 14968
rect 13924 14822 13952 20431
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14002 16008 14058 16017
rect 14002 15943 14058 15952
rect 14016 15706 14044 15943
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14016 15314 14044 15642
rect 14016 15286 14136 15314
rect 14002 15192 14058 15201
rect 14002 15127 14058 15136
rect 14016 15094 14044 15127
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13464 14006 13492 14758
rect 14016 14618 14044 15030
rect 14108 14890 14136 15286
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 14094 13560 14150 13569
rect 14094 13495 14150 13504
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12714 12336 12770 12345
rect 12714 12271 12716 12280
rect 12768 12271 12770 12280
rect 12716 12242 12768 12248
rect 12622 12200 12678 12209
rect 12622 12135 12678 12144
rect 12636 11354 12664 12135
rect 12728 11898 12756 12242
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13818 11928 13874 11937
rect 12716 11892 12768 11898
rect 13818 11863 13820 11872
rect 12716 11834 12768 11840
rect 13872 11863 13874 11872
rect 13820 11834 13872 11840
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12728 10470 12756 11086
rect 12820 10810 12848 11086
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12808 10600 12860 10606
rect 12806 10568 12808 10577
rect 12860 10568 12862 10577
rect 12806 10503 12862 10512
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12716 10464 12768 10470
rect 12912 10441 12940 10474
rect 12716 10406 12768 10412
rect 12898 10432 12954 10441
rect 12898 10367 12954 10376
rect 12808 9920 12860 9926
rect 12806 9888 12808 9897
rect 12860 9888 12862 9897
rect 12806 9823 12862 9832
rect 13004 9489 13032 10610
rect 12990 9480 13046 9489
rect 12716 9444 12768 9450
rect 12990 9415 13046 9424
rect 12716 9386 12768 9392
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12440 6928 12492 6934
rect 12360 6888 12440 6916
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12360 6390 12388 6888
rect 12440 6870 12492 6876
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 12452 6458 12480 6695
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12728 5234 12756 9386
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12820 8906 12848 9114
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7546 12940 7822
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13004 7410 13032 8230
rect 13096 8090 13124 8434
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12898 6352 12954 6361
rect 12898 6287 12900 6296
rect 12952 6287 12954 6296
rect 12992 6316 13044 6322
rect 12900 6258 12952 6264
rect 12992 6258 13044 6264
rect 13004 5914 13032 6258
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12728 5098 12756 5170
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12360 4706 12388 5034
rect 13188 4842 13216 11222
rect 13280 11150 13308 11698
rect 13268 11144 13320 11150
rect 13266 11112 13268 11121
rect 13320 11112 13322 11121
rect 13266 11047 13322 11056
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13372 10266 13400 10406
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13924 9602 13952 12038
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13832 9574 13952 9602
rect 13556 9382 13584 9522
rect 13544 9376 13596 9382
rect 13542 9344 13544 9353
rect 13596 9344 13598 9353
rect 13542 9279 13598 9288
rect 13556 9110 13584 9279
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13726 9072 13782 9081
rect 13452 9036 13504 9042
rect 13726 9007 13782 9016
rect 13452 8978 13504 8984
rect 13464 8838 13492 8978
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8294 13492 8774
rect 13740 8537 13768 9007
rect 13832 8650 13860 9574
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13924 9178 13952 9386
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13832 8622 13952 8650
rect 13820 8560 13872 8566
rect 13726 8528 13782 8537
rect 13820 8502 13872 8508
rect 13726 8463 13782 8472
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13832 8090 13860 8502
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13280 7546 13308 7890
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 12820 4814 13216 4842
rect 12360 4678 12480 4706
rect 12162 4040 12218 4049
rect 12162 3975 12218 3984
rect 12176 3738 12204 3975
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12084 2502 12204 2530
rect 12452 2514 12480 4678
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12544 3194 12572 3538
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12728 3194 12756 3470
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12544 2961 12572 3130
rect 12530 2952 12586 2961
rect 12530 2887 12586 2896
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12636 2553 12664 2586
rect 12622 2544 12678 2553
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12084 2281 12112 2382
rect 12070 2272 12126 2281
rect 12070 2207 12126 2216
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 12176 610 12204 2502
rect 12440 2508 12492 2514
rect 12622 2479 12678 2488
rect 12440 2450 12492 2456
rect 12452 2378 12480 2450
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12452 2145 12480 2314
rect 12438 2136 12494 2145
rect 12438 2071 12494 2080
rect 12164 604 12216 610
rect 12164 546 12216 552
rect 12256 604 12308 610
rect 12256 546 12308 552
rect 12268 480 12296 546
rect 12820 480 12848 4814
rect 12990 4584 13046 4593
rect 12990 4519 12992 4528
rect 13044 4519 13046 4528
rect 12992 4490 13044 4496
rect 13004 4078 13032 4490
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13280 3466 13308 3946
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13280 2990 13308 3402
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13096 2009 13124 2382
rect 13082 2000 13138 2009
rect 13082 1935 13138 1944
rect 13372 480 13400 7414
rect 13464 7342 13492 7686
rect 13648 7449 13676 7686
rect 13634 7440 13690 7449
rect 13634 7375 13690 7384
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 7002 13492 7278
rect 13832 7002 13860 8026
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13464 5914 13492 6938
rect 13634 6080 13690 6089
rect 13634 6015 13690 6024
rect 13648 5914 13676 6015
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13464 5234 13492 5850
rect 13740 5794 13768 5850
rect 13648 5766 13768 5794
rect 13648 5370 13676 5766
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13740 5012 13768 5238
rect 13832 5012 13860 5646
rect 13740 4984 13860 5012
rect 13740 4826 13768 4984
rect 13924 4865 13952 8622
rect 14016 8537 14044 9318
rect 14002 8528 14058 8537
rect 14002 8463 14058 8472
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 6730 14044 7142
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6322 14044 6666
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14002 5944 14058 5953
rect 14002 5879 14004 5888
rect 14056 5879 14058 5888
rect 14004 5850 14056 5856
rect 13910 4856 13966 4865
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13832 4814 13910 4842
rect 13832 4706 13860 4814
rect 13910 4791 13966 4800
rect 14108 4740 14136 13495
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 11898 14228 12582
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 9042 14320 9862
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14200 8294 14228 8366
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 8090 14228 8230
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14292 5710 14320 6122
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14292 5370 14320 5646
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13740 4678 13860 4706
rect 13924 4712 14136 4740
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 2990 13584 3878
rect 13544 2984 13596 2990
rect 13542 2952 13544 2961
rect 13596 2952 13598 2961
rect 13542 2887 13598 2896
rect 13740 2650 13768 4678
rect 13924 3720 13952 4712
rect 14200 4554 14228 5102
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 13832 3692 13952 3720
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13740 2446 13768 2586
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13832 610 13860 3692
rect 14292 3641 14320 4422
rect 14278 3632 14334 3641
rect 13912 3596 13964 3602
rect 14278 3567 14334 3576
rect 13912 3538 13964 3544
rect 13924 3233 13952 3538
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13910 3224 13966 3233
rect 13910 3159 13966 3168
rect 14108 2689 14136 3470
rect 14094 2680 14150 2689
rect 14094 2615 14150 2624
rect 14186 2544 14242 2553
rect 14186 2479 14188 2488
rect 14240 2479 14242 2488
rect 14188 2450 14240 2456
rect 13820 604 13872 610
rect 13820 546 13872 552
rect 13912 604 13964 610
rect 13912 546 13964 552
rect 13924 480 13952 546
rect 14384 480 14412 19110
rect 15304 18737 15332 23559
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 23478 23352 23534 23361
rect 23478 23287 23534 23296
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 23492 20369 23520 23287
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 23478 20360 23534 20369
rect 23478 20295 23534 20304
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 15290 18728 15346 18737
rect 15290 18663 15346 18672
rect 26238 18728 26294 18737
rect 26238 18663 26294 18672
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 23662 16144 23718 16153
rect 23662 16079 23718 16088
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 14830 15600 14886 15609
rect 14830 15535 14886 15544
rect 14844 14521 14872 15535
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 14830 14512 14886 14521
rect 14830 14447 14886 14456
rect 23386 14512 23442 14521
rect 23386 14447 23388 14456
rect 23440 14447 23442 14456
rect 23388 14418 23440 14424
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 23400 14074 23428 14418
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23570 13968 23626 13977
rect 23570 13903 23626 13912
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 22388 12782 22416 13330
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 22376 12776 22428 12782
rect 22374 12744 22376 12753
rect 22428 12744 22430 12753
rect 22374 12679 22430 12688
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 21836 11694 21864 12242
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21824 11688 21876 11694
rect 21822 11656 21824 11665
rect 21876 11656 21878 11665
rect 21822 11591 21878 11600
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 22020 11121 22048 12038
rect 22006 11112 22062 11121
rect 22006 11047 22062 11056
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15750 10704 15806 10713
rect 15750 10639 15806 10648
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14568 9586 14596 9930
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 9178 14504 9454
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14568 8906 14596 9522
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15580 8566 15608 8978
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 14462 8392 14518 8401
rect 14462 8327 14464 8336
rect 14516 8327 14518 8336
rect 14464 8298 14516 8304
rect 15212 7886 15240 8502
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 6866 14688 7754
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14660 5914 14688 6802
rect 14752 6254 14780 7142
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 6769 15424 6802
rect 15660 6792 15712 6798
rect 15382 6760 15438 6769
rect 15660 6734 15712 6740
rect 15382 6695 15438 6704
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15396 6458 15424 6695
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15290 6352 15346 6361
rect 15290 6287 15346 6296
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 15304 5778 15332 6287
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5817 15516 6054
rect 15474 5808 15530 5817
rect 15292 5772 15344 5778
rect 15474 5743 15530 5752
rect 15292 5714 15344 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14738 5400 14794 5409
rect 14956 5392 15252 5412
rect 14738 5335 14740 5344
rect 14792 5335 14794 5344
rect 14740 5306 14792 5312
rect 15304 5114 15332 5714
rect 15476 5704 15528 5710
rect 15474 5672 15476 5681
rect 15528 5672 15530 5681
rect 15474 5607 15530 5616
rect 14464 5092 14516 5098
rect 15304 5086 15424 5114
rect 14464 5034 14516 5040
rect 14476 4690 14504 5034
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15198 4992 15254 5001
rect 15028 4758 15056 4966
rect 15198 4927 15254 4936
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 15212 4690 15240 4927
rect 15396 4826 15424 5086
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14476 4282 14504 4626
rect 15212 4570 15240 4626
rect 15212 4542 15332 4570
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 15304 4214 15332 4542
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15488 4146 15516 4694
rect 15672 4321 15700 6734
rect 15658 4312 15714 4321
rect 15658 4247 15714 4256
rect 15476 4140 15528 4146
rect 15396 4100 15476 4128
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14752 3194 14780 3538
rect 15292 3528 15344 3534
rect 15396 3516 15424 4100
rect 15476 4082 15528 4088
rect 15344 3488 15424 3516
rect 15292 3470 15344 3476
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 15396 2582 15424 3488
rect 15566 3496 15622 3505
rect 15566 3431 15622 3440
rect 15580 3194 15608 3431
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15764 3126 15792 10639
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19338 10024 19394 10033
rect 19338 9959 19340 9968
rect 19392 9959 19394 9968
rect 19340 9930 19392 9936
rect 16670 9344 16726 9353
rect 16670 9279 16726 9288
rect 16684 9178 16712 9279
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 19982 9072 20038 9081
rect 19982 9007 20038 9016
rect 18234 8936 18290 8945
rect 18234 8871 18290 8880
rect 18142 8392 18198 8401
rect 16672 8356 16724 8362
rect 18142 8327 18198 8336
rect 16672 8298 16724 8304
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15856 7954 15884 8026
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15856 7546 15884 7890
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 16210 7304 16266 7313
rect 16210 7239 16212 7248
rect 16264 7239 16266 7248
rect 16212 7210 16264 7216
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16396 6112 16448 6118
rect 16394 6080 16396 6089
rect 16448 6080 16450 6089
rect 16394 6015 16450 6024
rect 16592 5914 16620 7142
rect 16684 5953 16712 8298
rect 18156 8090 18184 8327
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 7410 16988 7686
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 6934 16804 7142
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16960 6866 16988 7346
rect 17328 7206 17356 7890
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16670 5944 16726 5953
rect 16580 5908 16632 5914
rect 16670 5879 16726 5888
rect 16580 5850 16632 5856
rect 16776 5642 16804 6190
rect 16868 6100 16896 6734
rect 16960 6458 16988 6802
rect 17328 6610 17356 7142
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17500 6656 17552 6662
rect 17328 6604 17500 6610
rect 17328 6598 17552 6604
rect 17328 6582 17540 6598
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16948 6112 17000 6118
rect 16868 6072 16948 6100
rect 16948 6054 17000 6060
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 4690 16896 5102
rect 17236 4826 17264 5850
rect 17328 5710 17356 6582
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17328 5370 17356 5646
rect 17420 5642 17448 6394
rect 17880 6322 17908 6870
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 18050 6216 18106 6225
rect 17592 6180 17644 6186
rect 18050 6151 18106 6160
rect 17592 6122 17644 6128
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17420 5370 17448 5578
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15764 2650 15792 2790
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15212 2417 15240 2450
rect 16040 2446 16068 3946
rect 16224 2514 16252 4558
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16684 3738 16712 3946
rect 16868 3942 16896 4626
rect 17512 4060 17540 4966
rect 17604 4690 17632 6122
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17972 5658 18000 5714
rect 17880 5630 18000 5658
rect 17880 5386 17908 5630
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17788 5358 17908 5386
rect 17788 5166 17816 5358
rect 17776 5160 17828 5166
rect 17774 5128 17776 5137
rect 17828 5128 17830 5137
rect 17972 5098 18000 5510
rect 17774 5063 17830 5072
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17972 4486 18000 5034
rect 17960 4480 18012 4486
rect 17880 4428 17960 4434
rect 17880 4422 18012 4428
rect 17880 4406 18000 4422
rect 17880 4146 17908 4406
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17592 4072 17644 4078
rect 17512 4032 17592 4060
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3738 16896 3878
rect 17406 3768 17462 3777
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16856 3732 16908 3738
rect 17406 3703 17408 3712
rect 16856 3674 16908 3680
rect 17460 3703 17462 3712
rect 17408 3674 17460 3680
rect 17130 3632 17186 3641
rect 16396 3596 16448 3602
rect 17130 3567 17186 3576
rect 16396 3538 16448 3544
rect 16408 3058 16436 3538
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16028 2440 16080 2446
rect 15198 2408 15254 2417
rect 15198 2343 15254 2352
rect 15474 2408 15530 2417
rect 16028 2382 16080 2388
rect 15474 2343 15476 2352
rect 15528 2343 15530 2352
rect 16120 2372 16172 2378
rect 15476 2314 15528 2320
rect 16120 2314 16172 2320
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14924 2032 14976 2038
rect 14924 1974 14976 1980
rect 14936 480 14964 1974
rect 15396 1170 15424 2246
rect 16132 1170 16160 2314
rect 16578 1456 16634 1465
rect 16578 1391 16634 1400
rect 15396 1142 15516 1170
rect 15488 480 15516 1142
rect 16040 1142 16160 1170
rect 16040 480 16068 1142
rect 16592 480 16620 1391
rect 17144 480 17172 3567
rect 17420 3194 17448 3674
rect 17512 3670 17540 4032
rect 18064 4026 18092 6151
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5166 18184 6054
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18156 4826 18184 5102
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17592 4014 17644 4020
rect 17972 3998 18092 4026
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17682 3088 17738 3097
rect 17682 3023 17738 3032
rect 17696 480 17724 3023
rect 17972 2990 18000 3998
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18142 3904 18198 3913
rect 18064 3369 18092 3878
rect 18142 3839 18198 3848
rect 18156 3602 18184 3839
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18050 3360 18106 3369
rect 18050 3295 18106 3304
rect 18156 3194 18184 3538
rect 18248 3534 18276 8871
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19062 7848 19118 7857
rect 19062 7783 19118 7792
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18892 4486 18920 5782
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18418 4040 18474 4049
rect 18418 3975 18420 3984
rect 18472 3975 18474 3984
rect 18420 3946 18472 3952
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 3346 18276 3470
rect 18248 3318 18368 3346
rect 18234 3224 18290 3233
rect 18144 3188 18196 3194
rect 18340 3194 18368 3318
rect 18234 3159 18290 3168
rect 18328 3188 18380 3194
rect 18144 3130 18196 3136
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17972 2650 18000 2926
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18248 480 18276 3159
rect 18328 3130 18380 3136
rect 18524 3058 18552 3674
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18708 2961 18736 2994
rect 18694 2952 18750 2961
rect 18694 2887 18750 2896
rect 18510 2544 18566 2553
rect 18328 2508 18380 2514
rect 18510 2479 18566 2488
rect 18328 2450 18380 2456
rect 18340 1873 18368 2450
rect 18524 2446 18552 2479
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18326 1864 18382 1873
rect 18326 1799 18382 1808
rect 18800 480 18828 4082
rect 18892 2961 18920 4422
rect 19076 4078 19104 7783
rect 19706 7440 19762 7449
rect 19706 7375 19762 7384
rect 19720 7342 19748 7375
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19522 6896 19578 6905
rect 19522 6831 19578 6840
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19352 5370 19380 5578
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5166 19472 6122
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19352 3754 19380 4626
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4214 19472 4422
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19536 4146 19564 6831
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19890 4584 19946 4593
rect 19890 4519 19946 4528
rect 19904 4486 19932 4519
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19904 4214 19932 4422
rect 19892 4208 19944 4214
rect 19892 4150 19944 4156
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19352 3726 19472 3754
rect 19536 3738 19564 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19444 3670 19472 3726
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 18878 2952 18934 2961
rect 18878 2887 18934 2896
rect 18892 2009 18920 2887
rect 19352 2514 19380 3062
rect 19444 2650 19472 3402
rect 19628 3097 19656 3470
rect 19614 3088 19670 3097
rect 19614 3023 19670 3032
rect 19996 2990 20024 9007
rect 20258 8528 20314 8537
rect 20258 8463 20314 8472
rect 20272 8430 20300 8463
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20364 3505 20392 8298
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20732 6866 20760 7210
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20732 6458 20760 6802
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20902 4312 20958 4321
rect 20902 4247 20958 4256
rect 20720 4072 20772 4078
rect 20548 4032 20720 4060
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20350 3496 20406 3505
rect 20350 3431 20406 3440
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 18878 2000 18934 2009
rect 18878 1935 18934 1944
rect 19338 1456 19394 1465
rect 19338 1391 19394 1400
rect 19352 480 19380 1391
rect 20180 898 20208 2790
rect 19904 870 20208 898
rect 19904 480 19932 870
rect 20456 480 20484 3946
rect 20548 2582 20576 4032
rect 20720 4014 20772 4020
rect 20916 3602 20944 4247
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20810 3360 20866 3369
rect 20732 3233 20760 3334
rect 20810 3295 20866 3304
rect 20718 3224 20774 3233
rect 20824 3194 20852 3295
rect 20916 3194 20944 3538
rect 20718 3159 20774 3168
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20824 2990 20852 3130
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20536 2576 20588 2582
rect 20640 2553 20668 2858
rect 20536 2518 20588 2524
rect 20626 2544 20682 2553
rect 20626 2479 20682 2488
rect 21008 480 21036 4422
rect 21100 3942 21128 4626
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 2582 21128 3878
rect 21548 3392 21600 3398
rect 21652 3369 21680 6598
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 21548 3334 21600 3340
rect 21638 3360 21694 3369
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21192 2417 21220 2450
rect 21178 2408 21234 2417
rect 21178 2343 21234 2352
rect 21560 480 21588 3334
rect 21638 3295 21694 3304
rect 22020 3194 22048 3538
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22112 480 22140 4966
rect 22282 4040 22338 4049
rect 22282 3975 22284 3984
rect 22336 3975 22338 3984
rect 22284 3946 22336 3952
rect 22558 3360 22614 3369
rect 22558 3295 22614 3304
rect 22190 3088 22246 3097
rect 22190 3023 22246 3032
rect 22204 2990 22232 3023
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22466 2544 22522 2553
rect 22466 2479 22468 2488
rect 22520 2479 22522 2488
rect 22468 2450 22520 2456
rect 22572 1306 22600 3295
rect 23204 3120 23256 3126
rect 23204 3062 23256 3068
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22664 1465 22692 2246
rect 22650 1456 22706 1465
rect 22650 1391 22706 1400
rect 22572 1278 22692 1306
rect 22664 480 22692 1278
rect 23216 480 23244 3062
rect 23492 2038 23520 13126
rect 23584 12345 23612 13903
rect 23676 13870 23704 16079
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 23570 12336 23626 12345
rect 23570 12271 23626 12280
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 23662 11112 23718 11121
rect 23662 11047 23718 11056
rect 23570 3496 23626 3505
rect 23570 3431 23626 3440
rect 23584 3194 23612 3431
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23584 2990 23612 3130
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23480 2032 23532 2038
rect 23480 1974 23532 1980
rect 23676 626 23704 11047
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24124 9988 24176 9994
rect 24124 9930 24176 9936
rect 24136 4729 24164 9930
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24122 4720 24178 4729
rect 24122 4655 24178 4664
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24030 4176 24086 4185
rect 24030 4111 24086 4120
rect 24044 3602 24072 4111
rect 24032 3596 24084 3602
rect 24032 3538 24084 3544
rect 24044 3194 24072 3538
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24228 3097 24256 3334
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24214 3088 24270 3097
rect 24214 3023 24270 3032
rect 24766 2816 24822 2825
rect 24766 2751 24822 2760
rect 24780 2650 24808 2751
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24308 2032 24360 2038
rect 24308 1974 24360 1980
rect 23676 598 23796 626
rect 23768 480 23796 598
rect 24320 480 24348 1974
rect 24872 480 24900 13942
rect 24964 610 24992 14214
rect 25962 3088 26018 3097
rect 25962 3023 26018 3032
rect 24952 604 25004 610
rect 24952 546 25004 552
rect 25412 604 25464 610
rect 25412 546 25464 552
rect 25424 480 25452 546
rect 25976 480 26004 3023
rect 26252 610 26280 18663
rect 26514 2952 26570 2961
rect 26514 2887 26570 2896
rect 26240 604 26292 610
rect 26240 546 26292 552
rect 26528 480 26556 2887
rect 27618 2816 27674 2825
rect 27618 2751 27674 2760
rect 27068 604 27120 610
rect 27068 546 27120 552
rect 27080 480 27108 546
rect 27632 480 27660 2751
rect 1122 368 1178 377
rect 1122 303 1178 312
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3974 0 4030 480
rect 4526 0 4582 480
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6734 0 6790 480
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 8942 0 8998 480
rect 9494 0 9550 480
rect 10046 0 10102 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14370 0 14426 480
rect 14922 0 14978 480
rect 15474 0 15530 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17682 0 17738 480
rect 18234 0 18290 480
rect 18786 0 18842 480
rect 19338 0 19394 480
rect 19890 0 19946 480
rect 20442 0 20498 480
rect 20994 0 21050 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3238 27648 3294 27704
rect 1582 26560 1638 26616
rect 4158 27104 4214 27160
rect 3146 26016 3202 26072
rect 2686 25336 2742 25392
rect 1582 24792 1638 24848
rect 1582 24248 1638 24304
rect 1674 23432 1730 23488
rect 2410 22500 2466 22536
rect 2410 22480 2412 22500
rect 2412 22480 2464 22500
rect 2464 22480 2466 22500
rect 3054 23704 3110 23760
rect 3606 23296 3662 23352
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 7470 23588 7526 23624
rect 7470 23568 7472 23588
rect 7472 23568 7524 23588
rect 7524 23568 7526 23588
rect 9218 23432 9274 23488
rect 6274 23296 6330 23352
rect 4250 23160 4306 23216
rect 2778 22072 2834 22128
rect 2594 21800 2650 21856
rect 1950 21412 2006 21448
rect 1950 21392 1952 21412
rect 1952 21392 2004 21412
rect 2004 21392 2006 21412
rect 3514 21936 3570 21992
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 4434 22344 4490 22400
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 4250 21428 4252 21448
rect 4252 21428 4304 21448
rect 4304 21428 4306 21448
rect 4250 21392 4306 21428
rect 3790 21120 3846 21176
rect 5538 21256 5594 21312
rect 2962 20984 3018 21040
rect 2502 20440 2558 20496
rect 3054 20304 3110 20360
rect 4250 20848 4306 20904
rect 2318 19352 2374 19408
rect 2226 18400 2282 18456
rect 1582 17992 1638 18048
rect 1490 16224 1546 16280
rect 1674 17040 1730 17096
rect 1398 15272 1454 15328
rect 1766 16632 1822 16688
rect 1858 15544 1914 15600
rect 1674 15000 1730 15056
rect 1858 14728 1914 14784
rect 2226 14864 2282 14920
rect 2134 12588 2136 12608
rect 2136 12588 2188 12608
rect 2188 12588 2190 12608
rect 2134 12552 2190 12588
rect 1950 12416 2006 12472
rect 1766 12300 1822 12336
rect 1766 12280 1768 12300
rect 1768 12280 1820 12300
rect 1820 12280 1822 12300
rect 662 1808 718 1864
rect 1858 9324 1860 9344
rect 1860 9324 1912 9344
rect 1912 9324 1914 9344
rect 1858 9288 1914 9324
rect 2962 19660 2964 19680
rect 2964 19660 3016 19680
rect 3016 19660 3018 19680
rect 2962 19624 3018 19660
rect 2962 19080 3018 19136
rect 2870 18536 2926 18592
rect 2686 17856 2742 17912
rect 8114 21972 8116 21992
rect 8116 21972 8168 21992
rect 8168 21972 8170 21992
rect 8114 21936 8170 21972
rect 8022 21292 8024 21312
rect 8024 21292 8076 21312
rect 8076 21292 8078 21312
rect 8022 21256 8078 21292
rect 8758 21120 8814 21176
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 4434 19116 4436 19136
rect 4436 19116 4488 19136
rect 4488 19116 4490 19136
rect 4434 19080 4490 19116
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4250 18400 4306 18456
rect 2502 16904 2558 16960
rect 4066 17448 4122 17504
rect 3238 17040 3294 17096
rect 2778 16496 2834 16552
rect 2502 15952 2558 16008
rect 2410 15852 2412 15872
rect 2412 15852 2464 15872
rect 2464 15852 2466 15872
rect 2410 15816 2466 15852
rect 2778 15816 2834 15872
rect 2410 13912 2466 13968
rect 2870 14068 2926 14104
rect 2870 14048 2872 14068
rect 2872 14048 2924 14068
rect 2924 14048 2926 14068
rect 2962 12436 3018 12472
rect 2962 12416 2964 12436
rect 2964 12416 3016 12436
rect 3016 12416 3018 12436
rect 1030 856 1086 912
rect 2594 9152 2650 9208
rect 2502 8880 2558 8936
rect 2962 11736 3018 11792
rect 3790 16668 3792 16688
rect 3792 16668 3844 16688
rect 3844 16668 3846 16688
rect 3790 16632 3846 16668
rect 3974 15952 4030 16008
rect 3882 15444 3884 15464
rect 3884 15444 3936 15464
rect 3936 15444 3938 15464
rect 3882 15408 3938 15444
rect 3974 15136 4030 15192
rect 3790 14592 3846 14648
rect 4434 17856 4490 17912
rect 4342 16652 4398 16688
rect 4342 16632 4344 16652
rect 4344 16632 4396 16652
rect 4396 16632 4398 16652
rect 4158 15544 4214 15600
rect 3330 12824 3386 12880
rect 3238 12416 3294 12472
rect 3238 11600 3294 11656
rect 1398 7404 1454 7440
rect 1398 7384 1400 7404
rect 1400 7384 1452 7404
rect 1452 7384 1454 7404
rect 1674 7520 1730 7576
rect 1950 6160 2006 6216
rect 1858 6024 1914 6080
rect 1674 3304 1730 3360
rect 1858 2760 1914 2816
rect 1582 2488 1638 2544
rect 2410 8064 2466 8120
rect 2318 6840 2374 6896
rect 3146 9696 3202 9752
rect 2502 4936 2558 4992
rect 2410 3732 2466 3768
rect 2410 3712 2412 3732
rect 2412 3712 2464 3732
rect 2464 3712 2466 3732
rect 2134 1944 2190 2000
rect 1766 1672 1822 1728
rect 1306 1400 1362 1456
rect 2962 4256 3018 4312
rect 2686 3848 2742 3904
rect 3606 13776 3662 13832
rect 3422 12144 3478 12200
rect 3330 9832 3386 9888
rect 4066 14476 4122 14512
rect 4066 14456 4068 14476
rect 4068 14456 4120 14476
rect 4120 14456 4122 14476
rect 7010 19352 7066 19408
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 4986 16904 5042 16960
rect 5170 16940 5172 16960
rect 5172 16940 5224 16960
rect 5224 16940 5226 16960
rect 5170 16904 5226 16940
rect 4802 16088 4858 16144
rect 4710 15544 4766 15600
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 4894 15408 4950 15464
rect 4802 15272 4858 15328
rect 4802 14728 4858 14784
rect 3882 13368 3938 13424
rect 3790 12688 3846 12744
rect 3790 12416 3846 12472
rect 3606 11600 3662 11656
rect 3514 8916 3516 8936
rect 3516 8916 3568 8936
rect 3568 8916 3570 8936
rect 3514 8880 3570 8916
rect 3422 7248 3478 7304
rect 3698 8472 3754 8528
rect 3514 6704 3570 6760
rect 3606 4800 3662 4856
rect 3330 4528 3386 4584
rect 3054 3984 3110 4040
rect 3054 3440 3110 3496
rect 3606 4120 3662 4176
rect 2686 2760 2742 2816
rect 2870 2760 2926 2816
rect 3974 12280 4030 12336
rect 4526 13640 4582 13696
rect 4342 12164 4398 12200
rect 4342 12144 4344 12164
rect 4344 12144 4396 12164
rect 4396 12144 4398 12164
rect 4802 12300 4858 12336
rect 4802 12280 4804 12300
rect 4804 12280 4856 12300
rect 4856 12280 4858 12300
rect 4158 11500 4160 11520
rect 4160 11500 4212 11520
rect 4212 11500 4214 11520
rect 4158 11464 4214 11500
rect 3974 11328 4030 11384
rect 4158 11212 4214 11248
rect 4158 11192 4160 11212
rect 4160 11192 4212 11212
rect 4212 11192 4214 11212
rect 3882 10104 3938 10160
rect 3974 9968 4030 10024
rect 3882 9424 3938 9480
rect 3790 8336 3846 8392
rect 4250 9288 4306 9344
rect 3974 9016 4030 9072
rect 3974 8336 4030 8392
rect 5446 14900 5448 14920
rect 5448 14900 5500 14920
rect 5500 14900 5502 14920
rect 5446 14864 5502 14900
rect 5814 16768 5870 16824
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5262 14592 5318 14648
rect 4986 13912 5042 13968
rect 5262 13404 5264 13424
rect 5264 13404 5316 13424
rect 5316 13404 5318 13424
rect 5262 13368 5318 13404
rect 5722 14456 5778 14512
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6550 15852 6552 15872
rect 6552 15852 6604 15872
rect 6604 15852 6606 15872
rect 6550 15816 6606 15852
rect 6826 16496 6882 16552
rect 6550 15036 6552 15056
rect 6552 15036 6604 15056
rect 6604 15036 6606 15056
rect 6550 15000 6606 15036
rect 6550 14184 6606 14240
rect 6182 13912 6238 13968
rect 5998 12552 6054 12608
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5814 11056 5870 11112
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5078 10512 5134 10568
rect 4894 10240 4950 10296
rect 4986 9172 5042 9208
rect 4986 9152 4988 9172
rect 4988 9152 5040 9172
rect 5040 9152 5042 9172
rect 3882 5616 3938 5672
rect 4158 7540 4214 7576
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5630 9580 5686 9616
rect 5630 9560 5632 9580
rect 5632 9560 5684 9580
rect 5684 9560 5686 9580
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 4618 8064 4674 8120
rect 5538 8472 5594 8528
rect 4158 7520 4160 7540
rect 4160 7520 4212 7540
rect 4212 7520 4214 7540
rect 4250 6568 4306 6624
rect 3974 3576 4030 3632
rect 3698 3168 3754 3224
rect 4526 3984 4582 4040
rect 4250 3340 4252 3360
rect 4252 3340 4304 3360
rect 4304 3340 4306 3360
rect 4250 3304 4306 3340
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5354 7112 5410 7168
rect 5262 6840 5318 6896
rect 5078 5072 5134 5128
rect 4986 3712 5042 3768
rect 4618 2624 4674 2680
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6090 11736 6146 11792
rect 6826 13676 6828 13696
rect 6828 13676 6880 13696
rect 6880 13676 6882 13696
rect 6826 13640 6882 13676
rect 7194 19080 7250 19136
rect 8022 18028 8024 18048
rect 8024 18028 8076 18048
rect 8076 18028 8078 18048
rect 8022 17992 8078 18028
rect 8666 18420 8722 18456
rect 8666 18400 8668 18420
rect 8668 18400 8720 18420
rect 8720 18400 8722 18420
rect 7102 15020 7158 15056
rect 7102 15000 7104 15020
rect 7104 15000 7156 15020
rect 7156 15000 7158 15020
rect 6366 10920 6422 10976
rect 6918 11464 6974 11520
rect 6826 11328 6882 11384
rect 6642 10376 6698 10432
rect 6550 8356 6606 8392
rect 6550 8336 6552 8356
rect 6552 8336 6604 8356
rect 6604 8336 6606 8356
rect 7102 10512 7158 10568
rect 7102 9460 7104 9480
rect 7104 9460 7156 9480
rect 7156 9460 7158 9480
rect 7102 9424 7158 9460
rect 6642 7520 6698 7576
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5354 3848 5410 3904
rect 5170 3068 5172 3088
rect 5172 3068 5224 3088
rect 5224 3068 5226 3088
rect 5170 3032 5226 3068
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6458 6024 6514 6080
rect 6918 7384 6974 7440
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6642 1808 6698 1864
rect 7470 16088 7526 16144
rect 7286 15544 7342 15600
rect 7746 15408 7802 15464
rect 7930 12280 7986 12336
rect 8206 15428 8262 15464
rect 8206 15408 8208 15428
rect 8208 15408 8260 15428
rect 8260 15408 8262 15428
rect 8942 17448 8998 17504
rect 8850 16904 8906 16960
rect 8758 12416 8814 12472
rect 8022 10512 8078 10568
rect 7930 10240 7986 10296
rect 7654 8900 7710 8936
rect 7654 8880 7656 8900
rect 7656 8880 7708 8900
rect 7708 8880 7710 8900
rect 8022 9596 8024 9616
rect 8024 9596 8076 9616
rect 8076 9596 8078 9616
rect 8022 9560 8078 9596
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 15290 23568 15346 23624
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 9678 21256 9734 21312
rect 9770 17992 9826 18048
rect 9126 16632 9182 16688
rect 8942 12416 8998 12472
rect 7102 5072 7158 5128
rect 6918 2896 6974 2952
rect 8114 7792 8170 7848
rect 7746 7692 7748 7712
rect 7748 7692 7800 7712
rect 7800 7692 7802 7712
rect 7746 7656 7802 7692
rect 8574 8508 8576 8528
rect 8576 8508 8628 8528
rect 8628 8508 8630 8528
rect 8574 8472 8630 8508
rect 7378 5616 7434 5672
rect 7746 5208 7802 5264
rect 7470 2624 7526 2680
rect 7378 2216 7434 2272
rect 7562 2080 7618 2136
rect 8022 3304 8078 3360
rect 7930 1808 7986 1864
rect 8574 5752 8630 5808
rect 8298 5616 8354 5672
rect 8482 5072 8538 5128
rect 8298 3984 8354 4040
rect 8850 4528 8906 4584
rect 9034 3576 9090 3632
rect 8942 3440 8998 3496
rect 8942 3032 8998 3088
rect 9678 15952 9734 16008
rect 9310 14220 9312 14240
rect 9312 14220 9364 14240
rect 9364 14220 9366 14240
rect 9310 14184 9366 14220
rect 9494 15156 9550 15192
rect 9494 15136 9496 15156
rect 9496 15136 9548 15156
rect 9548 15136 9550 15156
rect 9770 15272 9826 15328
rect 9402 13232 9458 13288
rect 9954 22480 10010 22536
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10046 22072 10102 22128
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 11334 20984 11390 21040
rect 11518 20340 11520 20360
rect 11520 20340 11572 20360
rect 11572 20340 11574 20360
rect 11518 20304 11574 20340
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 13910 20440 13966 20496
rect 13818 20304 13874 20360
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 17040 10194 17096
rect 10782 17484 10784 17504
rect 10784 17484 10836 17504
rect 10836 17484 10838 17504
rect 10782 17448 10838 17484
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10966 15852 10968 15872
rect 10968 15852 11020 15872
rect 11020 15852 11022 15872
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10966 15816 11022 15852
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 11150 13232 11206 13288
rect 10690 10376 10746 10432
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10782 10004 10784 10024
rect 10784 10004 10836 10024
rect 10836 10004 10838 10024
rect 10782 9968 10838 10004
rect 10322 9832 10378 9888
rect 10690 9424 10746 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10506 9016 10562 9072
rect 10138 8880 10194 8936
rect 9862 7656 9918 7712
rect 9770 6568 9826 6624
rect 9862 6060 9864 6080
rect 9864 6060 9916 6080
rect 9916 6060 9918 6080
rect 9862 6024 9918 6060
rect 8666 2388 8668 2408
rect 8668 2388 8720 2408
rect 8720 2388 8722 2408
rect 8666 2352 8722 2388
rect 9218 2760 9274 2816
rect 9586 4528 9642 4584
rect 9402 1672 9458 1728
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 12070 18400 12126 18456
rect 11794 17040 11850 17096
rect 12438 15816 12494 15872
rect 12622 15408 12678 15464
rect 12530 15272 12586 15328
rect 11886 14884 11942 14920
rect 11886 14864 11888 14884
rect 11888 14864 11940 14884
rect 11940 14864 11942 14884
rect 11334 13504 11390 13560
rect 11058 11192 11114 11248
rect 12438 13368 12494 13424
rect 11794 10920 11850 10976
rect 10966 8336 11022 8392
rect 10966 7928 11022 7984
rect 10874 7792 10930 7848
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10506 6296 10562 6352
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11058 6160 11114 6216
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11518 10104 11574 10160
rect 11794 9696 11850 9752
rect 11702 8336 11758 8392
rect 11518 6704 11574 6760
rect 11334 6180 11390 6216
rect 11334 6160 11336 6180
rect 11336 6160 11388 6180
rect 11388 6160 11390 6180
rect 11242 5616 11298 5672
rect 11058 4936 11114 4992
rect 10874 4800 10930 4856
rect 9770 3440 9826 3496
rect 9678 2488 9734 2544
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3440 10194 3496
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11150 3576 11206 3632
rect 11058 3052 11114 3088
rect 11058 3032 11060 3052
rect 11060 3032 11112 3052
rect 11112 3032 11114 3052
rect 10598 992 10654 1048
rect 11518 5344 11574 5400
rect 11334 3884 11336 3904
rect 11336 3884 11388 3904
rect 11388 3884 11390 3904
rect 11334 3848 11390 3884
rect 11426 3068 11428 3088
rect 11428 3068 11480 3088
rect 11480 3068 11482 3088
rect 11426 3032 11482 3068
rect 11334 2644 11390 2680
rect 11334 2624 11336 2644
rect 11336 2624 11388 2644
rect 11388 2624 11390 2644
rect 11610 1400 11666 1456
rect 11886 3576 11942 3632
rect 11794 3304 11850 3360
rect 12346 11872 12402 11928
rect 12346 9594 12402 9650
rect 13818 15020 13874 15056
rect 13818 15000 13820 15020
rect 13820 15000 13872 15020
rect 13872 15000 13874 15020
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14002 15952 14058 16008
rect 14002 15136 14058 15192
rect 14094 13504 14150 13560
rect 12714 12300 12770 12336
rect 12714 12280 12716 12300
rect 12716 12280 12768 12300
rect 12768 12280 12770 12300
rect 12622 12144 12678 12200
rect 13818 11892 13874 11928
rect 13818 11872 13820 11892
rect 13820 11872 13872 11892
rect 13872 11872 13874 11892
rect 12806 10548 12808 10568
rect 12808 10548 12860 10568
rect 12860 10548 12862 10568
rect 12806 10512 12862 10548
rect 12898 10376 12954 10432
rect 12806 9868 12808 9888
rect 12808 9868 12860 9888
rect 12860 9868 12862 9888
rect 12806 9832 12862 9868
rect 12990 9424 13046 9480
rect 12438 6704 12494 6760
rect 12898 6316 12954 6352
rect 12898 6296 12900 6316
rect 12900 6296 12952 6316
rect 12952 6296 12954 6316
rect 13266 11092 13268 11112
rect 13268 11092 13320 11112
rect 13320 11092 13322 11112
rect 13266 11056 13322 11092
rect 13542 9324 13544 9344
rect 13544 9324 13596 9344
rect 13596 9324 13598 9344
rect 13542 9288 13598 9324
rect 13726 9016 13782 9072
rect 13726 8472 13782 8528
rect 12162 3984 12218 4040
rect 12530 2896 12586 2952
rect 12070 2216 12126 2272
rect 12622 2488 12678 2544
rect 12438 2080 12494 2136
rect 12990 4548 13046 4584
rect 12990 4528 12992 4548
rect 12992 4528 13044 4548
rect 13044 4528 13046 4548
rect 13082 1944 13138 2000
rect 13634 7384 13690 7440
rect 13634 6024 13690 6080
rect 14002 8472 14058 8528
rect 14002 5908 14058 5944
rect 14002 5888 14004 5908
rect 14004 5888 14056 5908
rect 14056 5888 14058 5908
rect 13910 4800 13966 4856
rect 13542 2932 13544 2952
rect 13544 2932 13596 2952
rect 13596 2932 13598 2952
rect 13542 2896 13598 2932
rect 14278 3576 14334 3632
rect 13910 3168 13966 3224
rect 14094 2624 14150 2680
rect 14186 2508 14242 2544
rect 14186 2488 14188 2508
rect 14188 2488 14240 2508
rect 14240 2488 14242 2508
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 23478 23296 23534 23352
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 23478 20304 23534 20360
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 15290 18672 15346 18728
rect 26238 18672 26294 18728
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 23662 16088 23718 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14830 15544 14886 15600
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 14830 14456 14886 14512
rect 23386 14476 23442 14512
rect 23386 14456 23388 14476
rect 23388 14456 23440 14476
rect 23440 14456 23442 14476
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 23570 13912 23626 13968
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 22374 12724 22376 12744
rect 22376 12724 22428 12744
rect 22428 12724 22430 12744
rect 22374 12688 22430 12724
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 21822 11636 21824 11656
rect 21824 11636 21876 11656
rect 21876 11636 21878 11656
rect 21822 11600 21878 11636
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 22006 11056 22062 11112
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15750 10648 15806 10704
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14462 8356 14518 8392
rect 14462 8336 14464 8356
rect 14464 8336 14516 8356
rect 14516 8336 14518 8356
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15382 6704 15438 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15290 6296 15346 6352
rect 15474 5752 15530 5808
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14738 5364 14794 5400
rect 14738 5344 14740 5364
rect 14740 5344 14792 5364
rect 14792 5344 14794 5364
rect 15474 5652 15476 5672
rect 15476 5652 15528 5672
rect 15528 5652 15530 5672
rect 15474 5616 15530 5652
rect 15198 4936 15254 4992
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15658 4256 15714 4312
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15566 3440 15622 3496
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19338 9988 19394 10024
rect 19338 9968 19340 9988
rect 19340 9968 19392 9988
rect 19392 9968 19394 9988
rect 16670 9288 16726 9344
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19982 9016 20038 9072
rect 18234 8880 18290 8936
rect 18142 8336 18198 8392
rect 16210 7268 16266 7304
rect 16210 7248 16212 7268
rect 16212 7248 16264 7268
rect 16264 7248 16266 7268
rect 16394 6060 16396 6080
rect 16396 6060 16448 6080
rect 16448 6060 16450 6080
rect 16394 6024 16450 6060
rect 16670 5888 16726 5944
rect 18050 6160 18106 6216
rect 17774 5108 17776 5128
rect 17776 5108 17828 5128
rect 17828 5108 17830 5128
rect 17774 5072 17830 5108
rect 17406 3732 17462 3768
rect 17406 3712 17408 3732
rect 17408 3712 17460 3732
rect 17460 3712 17462 3732
rect 17130 3576 17186 3632
rect 15198 2352 15254 2408
rect 15474 2372 15530 2408
rect 15474 2352 15476 2372
rect 15476 2352 15528 2372
rect 15528 2352 15530 2372
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16578 1400 16634 1456
rect 17682 3032 17738 3088
rect 18142 3848 18198 3904
rect 18050 3304 18106 3360
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19062 7792 19118 7848
rect 18418 4004 18474 4040
rect 18418 3984 18420 4004
rect 18420 3984 18472 4004
rect 18472 3984 18474 4004
rect 18234 3168 18290 3224
rect 18694 2896 18750 2952
rect 18510 2488 18566 2544
rect 18326 1808 18382 1864
rect 19706 7384 19762 7440
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19522 6840 19578 6896
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19890 4528 19946 4584
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 18878 2896 18934 2952
rect 19614 3032 19670 3088
rect 20258 8472 20314 8528
rect 20902 4256 20958 4312
rect 20350 3440 20406 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 18878 1944 18934 2000
rect 19338 1400 19394 1456
rect 20810 3304 20866 3360
rect 20718 3168 20774 3224
rect 20626 2488 20682 2544
rect 21178 2352 21234 2408
rect 21638 3304 21694 3360
rect 22282 4004 22338 4040
rect 22282 3984 22284 4004
rect 22284 3984 22336 4004
rect 22336 3984 22338 4004
rect 22558 3304 22614 3360
rect 22190 3032 22246 3088
rect 22466 2508 22522 2544
rect 22466 2488 22468 2508
rect 22468 2488 22520 2508
rect 22520 2488 22522 2508
rect 22650 1400 22706 1456
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 23570 12280 23626 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23662 11056 23718 11112
rect 23570 3440 23626 3496
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24122 4664 24178 4720
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24030 4120 24086 4176
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24214 3032 24270 3088
rect 24766 2760 24822 2816
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25962 3032 26018 3088
rect 26514 2896 26570 2952
rect 27618 2760 27674 2816
rect 1122 312 1178 368
<< metal3 >>
rect 0 27706 480 27736
rect 3233 27706 3299 27709
rect 0 27704 3299 27706
rect 0 27648 3238 27704
rect 3294 27648 3299 27704
rect 0 27646 3299 27648
rect 0 27616 480 27646
rect 3233 27643 3299 27646
rect 0 27162 480 27192
rect 4153 27162 4219 27165
rect 0 27160 4219 27162
rect 0 27104 4158 27160
rect 4214 27104 4219 27160
rect 0 27102 4219 27104
rect 0 27072 480 27102
rect 4153 27099 4219 27102
rect 0 26618 480 26648
rect 1577 26618 1643 26621
rect 0 26616 1643 26618
rect 0 26560 1582 26616
rect 1638 26560 1643 26616
rect 0 26558 1643 26560
rect 0 26528 480 26558
rect 1577 26555 1643 26558
rect 0 26074 480 26104
rect 3141 26074 3207 26077
rect 0 26072 3207 26074
rect 0 26016 3146 26072
rect 3202 26016 3207 26072
rect 0 26014 3207 26016
rect 0 25984 480 26014
rect 3141 26011 3207 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 2681 25394 2747 25397
rect 0 25392 2747 25394
rect 0 25336 2686 25392
rect 2742 25336 2747 25392
rect 0 25334 2747 25336
rect 0 25304 480 25334
rect 2681 25331 2747 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 1577 24850 1643 24853
rect 0 24848 1643 24850
rect 0 24792 1582 24848
rect 1638 24792 1643 24848
rect 0 24790 1643 24792
rect 0 24760 480 24790
rect 1577 24787 1643 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24306 480 24336
rect 1577 24306 1643 24309
rect 0 24304 1643 24306
rect 0 24248 1582 24304
rect 1638 24248 1643 24304
rect 0 24246 1643 24248
rect 0 24216 480 24246
rect 1577 24243 1643 24246
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 0 23762 480 23792
rect 3049 23762 3115 23765
rect 0 23760 3115 23762
rect 0 23704 3054 23760
rect 3110 23704 3115 23760
rect 0 23702 3115 23704
rect 0 23672 480 23702
rect 3049 23699 3115 23702
rect 7465 23626 7531 23629
rect 15285 23626 15351 23629
rect 7465 23624 15351 23626
rect 7465 23568 7470 23624
rect 7526 23568 15290 23624
rect 15346 23568 15351 23624
rect 7465 23566 15351 23568
rect 7465 23563 7531 23566
rect 15285 23563 15351 23566
rect 1669 23490 1735 23493
rect 9213 23490 9279 23493
rect 1669 23488 9279 23490
rect 1669 23432 1674 23488
rect 1730 23432 9218 23488
rect 9274 23432 9279 23488
rect 1669 23430 9279 23432
rect 1669 23427 1735 23430
rect 9213 23427 9279 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 3601 23354 3667 23357
rect 6269 23354 6335 23357
rect 3601 23352 6335 23354
rect 3601 23296 3606 23352
rect 3662 23296 6274 23352
rect 6330 23296 6335 23352
rect 3601 23294 6335 23296
rect 3601 23291 3667 23294
rect 6269 23291 6335 23294
rect 23473 23354 23539 23357
rect 27520 23354 28000 23384
rect 23473 23352 28000 23354
rect 23473 23296 23478 23352
rect 23534 23296 28000 23352
rect 23473 23294 28000 23296
rect 23473 23291 23539 23294
rect 27520 23264 28000 23294
rect 0 23218 480 23248
rect 4245 23218 4311 23221
rect 0 23216 4311 23218
rect 0 23160 4250 23216
rect 4306 23160 4311 23216
rect 0 23158 4311 23160
rect 0 23128 480 23158
rect 4245 23155 4311 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22538 480 22568
rect 2405 22538 2471 22541
rect 9949 22538 10015 22541
rect 0 22478 2330 22538
rect 0 22448 480 22478
rect 2270 22402 2330 22478
rect 2405 22536 10015 22538
rect 2405 22480 2410 22536
rect 2466 22480 9954 22536
rect 10010 22480 10015 22536
rect 2405 22478 10015 22480
rect 2405 22475 2471 22478
rect 9949 22475 10015 22478
rect 4429 22402 4495 22405
rect 2270 22400 4495 22402
rect 2270 22344 4434 22400
rect 4490 22344 4495 22400
rect 2270 22342 4495 22344
rect 4429 22339 4495 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 2773 22130 2839 22133
rect 10041 22130 10107 22133
rect 2773 22128 10107 22130
rect 2773 22072 2778 22128
rect 2834 22072 10046 22128
rect 10102 22072 10107 22128
rect 2773 22070 10107 22072
rect 2773 22067 2839 22070
rect 10041 22067 10107 22070
rect 0 21994 480 22024
rect 3509 21994 3575 21997
rect 8109 21994 8175 21997
rect 0 21992 3575 21994
rect 0 21936 3514 21992
rect 3570 21936 3575 21992
rect 0 21934 3575 21936
rect 0 21904 480 21934
rect 3509 21931 3575 21934
rect 5398 21992 8175 21994
rect 5398 21936 8114 21992
rect 8170 21936 8175 21992
rect 5398 21934 8175 21936
rect 2589 21858 2655 21861
rect 5398 21858 5458 21934
rect 8109 21931 8175 21934
rect 2589 21856 5458 21858
rect 2589 21800 2594 21856
rect 2650 21800 5458 21856
rect 2589 21798 5458 21800
rect 2589 21795 2655 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21450 480 21480
rect 1945 21450 2011 21453
rect 4245 21450 4311 21453
rect 0 21390 1410 21450
rect 0 21360 480 21390
rect 1350 21314 1410 21390
rect 1945 21448 4311 21450
rect 1945 21392 1950 21448
rect 2006 21392 4250 21448
rect 4306 21392 4311 21448
rect 1945 21390 4311 21392
rect 1945 21387 2011 21390
rect 4245 21387 4311 21390
rect 5533 21314 5599 21317
rect 1350 21312 5599 21314
rect 1350 21256 5538 21312
rect 5594 21256 5599 21312
rect 1350 21254 5599 21256
rect 5533 21251 5599 21254
rect 8017 21314 8083 21317
rect 9673 21314 9739 21317
rect 8017 21312 9739 21314
rect 8017 21256 8022 21312
rect 8078 21256 9678 21312
rect 9734 21256 9739 21312
rect 8017 21254 9739 21256
rect 8017 21251 8083 21254
rect 9673 21251 9739 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 3785 21178 3851 21181
rect 8753 21178 8819 21181
rect 3785 21176 8819 21178
rect 3785 21120 3790 21176
rect 3846 21120 8758 21176
rect 8814 21120 8819 21176
rect 3785 21118 8819 21120
rect 3785 21115 3851 21118
rect 8753 21115 8819 21118
rect 2957 21042 3023 21045
rect 11329 21042 11395 21045
rect 2957 21040 11395 21042
rect 2957 20984 2962 21040
rect 3018 20984 11334 21040
rect 11390 20984 11395 21040
rect 2957 20982 11395 20984
rect 2957 20979 3023 20982
rect 11329 20979 11395 20982
rect 0 20906 480 20936
rect 4245 20906 4311 20909
rect 0 20904 4311 20906
rect 0 20848 4250 20904
rect 4306 20848 4311 20904
rect 0 20846 4311 20848
rect 0 20816 480 20846
rect 4245 20843 4311 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 2497 20498 2563 20501
rect 13905 20498 13971 20501
rect 2497 20496 13971 20498
rect 2497 20440 2502 20496
rect 2558 20440 13910 20496
rect 13966 20440 13971 20496
rect 2497 20438 13971 20440
rect 2497 20435 2563 20438
rect 13905 20435 13971 20438
rect 0 20362 480 20392
rect 3049 20362 3115 20365
rect 0 20360 3115 20362
rect 0 20304 3054 20360
rect 3110 20304 3115 20360
rect 0 20302 3115 20304
rect 0 20272 480 20302
rect 3049 20299 3115 20302
rect 11513 20362 11579 20365
rect 13813 20362 13879 20365
rect 23473 20362 23539 20365
rect 11513 20360 23539 20362
rect 11513 20304 11518 20360
rect 11574 20304 13818 20360
rect 13874 20304 23478 20360
rect 23534 20304 23539 20360
rect 11513 20302 23539 20304
rect 11513 20299 11579 20302
rect 13813 20299 13879 20302
rect 23473 20299 23539 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19682 480 19712
rect 2957 19682 3023 19685
rect 0 19680 3023 19682
rect 0 19624 2962 19680
rect 3018 19624 3023 19680
rect 0 19622 3023 19624
rect 0 19592 480 19622
rect 2957 19619 3023 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 2313 19410 2379 19413
rect 7005 19410 7071 19413
rect 2313 19408 7071 19410
rect 2313 19352 2318 19408
rect 2374 19352 7010 19408
rect 7066 19352 7071 19408
rect 2313 19350 7071 19352
rect 2313 19347 2379 19350
rect 7005 19347 7071 19350
rect 0 19138 480 19168
rect 2957 19138 3023 19141
rect 0 19136 3023 19138
rect 0 19080 2962 19136
rect 3018 19080 3023 19136
rect 0 19078 3023 19080
rect 0 19048 480 19078
rect 2957 19075 3023 19078
rect 4429 19138 4495 19141
rect 7189 19138 7255 19141
rect 4429 19136 7255 19138
rect 4429 19080 4434 19136
rect 4490 19080 7194 19136
rect 7250 19080 7255 19136
rect 4429 19078 7255 19080
rect 4429 19075 4495 19078
rect 7189 19075 7255 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 15285 18730 15351 18733
rect 26233 18730 26299 18733
rect 15285 18728 26299 18730
rect 15285 18672 15290 18728
rect 15346 18672 26238 18728
rect 26294 18672 26299 18728
rect 15285 18670 26299 18672
rect 15285 18667 15351 18670
rect 26233 18667 26299 18670
rect 0 18594 480 18624
rect 2865 18594 2931 18597
rect 0 18592 2931 18594
rect 0 18536 2870 18592
rect 2926 18536 2931 18592
rect 0 18534 2931 18536
rect 0 18504 480 18534
rect 2865 18531 2931 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 2221 18458 2287 18461
rect 4245 18458 4311 18461
rect 2221 18456 4311 18458
rect 2221 18400 2226 18456
rect 2282 18400 4250 18456
rect 4306 18400 4311 18456
rect 2221 18398 4311 18400
rect 2221 18395 2287 18398
rect 4245 18395 4311 18398
rect 8661 18458 8727 18461
rect 12065 18458 12131 18461
rect 8661 18456 12131 18458
rect 8661 18400 8666 18456
rect 8722 18400 12070 18456
rect 12126 18400 12131 18456
rect 8661 18398 12131 18400
rect 8661 18395 8727 18398
rect 12065 18395 12131 18398
rect 0 18050 480 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 480 17990
rect 1577 17987 1643 17990
rect 8017 18050 8083 18053
rect 9765 18050 9831 18053
rect 8017 18048 9831 18050
rect 8017 17992 8022 18048
rect 8078 17992 9770 18048
rect 9826 17992 9831 18048
rect 8017 17990 9831 17992
rect 8017 17987 8083 17990
rect 9765 17987 9831 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 2681 17914 2747 17917
rect 4429 17914 4495 17917
rect 2681 17912 4495 17914
rect 2681 17856 2686 17912
rect 2742 17856 4434 17912
rect 4490 17856 4495 17912
rect 2681 17854 4495 17856
rect 2681 17851 2747 17854
rect 4429 17851 4495 17854
rect 0 17506 480 17536
rect 4061 17506 4127 17509
rect 0 17504 4127 17506
rect 0 17448 4066 17504
rect 4122 17448 4127 17504
rect 0 17446 4127 17448
rect 0 17416 480 17446
rect 4061 17443 4127 17446
rect 8937 17506 9003 17509
rect 10777 17506 10843 17509
rect 8937 17504 10843 17506
rect 8937 17448 8942 17504
rect 8998 17448 10782 17504
rect 10838 17448 10843 17504
rect 8937 17446 10843 17448
rect 8937 17443 9003 17446
rect 10777 17443 10843 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 1669 17098 1735 17101
rect 3233 17098 3299 17101
rect 10133 17098 10199 17101
rect 11789 17098 11855 17101
rect 1669 17096 11855 17098
rect 1669 17040 1674 17096
rect 1730 17040 3238 17096
rect 3294 17040 10138 17096
rect 10194 17040 11794 17096
rect 11850 17040 11855 17096
rect 1669 17038 11855 17040
rect 1669 17035 1735 17038
rect 3233 17035 3299 17038
rect 10133 17035 10199 17038
rect 11789 17035 11855 17038
rect 2497 16962 2563 16965
rect 4981 16962 5047 16965
rect 2497 16960 5047 16962
rect 2497 16904 2502 16960
rect 2558 16904 4986 16960
rect 5042 16904 5047 16960
rect 2497 16902 5047 16904
rect 2497 16899 2563 16902
rect 4981 16899 5047 16902
rect 5165 16962 5231 16965
rect 8845 16962 8911 16965
rect 5165 16960 8911 16962
rect 5165 16904 5170 16960
rect 5226 16904 8850 16960
rect 8906 16904 8911 16960
rect 5165 16902 8911 16904
rect 5165 16899 5231 16902
rect 8845 16899 8911 16902
rect 10277 16896 10597 16897
rect 0 16826 480 16856
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5809 16826 5875 16829
rect 0 16824 5875 16826
rect 0 16768 5814 16824
rect 5870 16768 5875 16824
rect 0 16766 5875 16768
rect 0 16736 480 16766
rect 5809 16763 5875 16766
rect 1761 16690 1827 16693
rect 3785 16690 3851 16693
rect 1761 16688 3851 16690
rect 1761 16632 1766 16688
rect 1822 16632 3790 16688
rect 3846 16632 3851 16688
rect 1761 16630 3851 16632
rect 1761 16627 1827 16630
rect 3785 16627 3851 16630
rect 4337 16690 4403 16693
rect 9121 16690 9187 16693
rect 4337 16688 9187 16690
rect 4337 16632 4342 16688
rect 4398 16632 9126 16688
rect 9182 16632 9187 16688
rect 4337 16630 9187 16632
rect 4337 16627 4403 16630
rect 9121 16627 9187 16630
rect 2773 16554 2839 16557
rect 6821 16554 6887 16557
rect 2773 16552 6887 16554
rect 2773 16496 2778 16552
rect 2834 16496 6826 16552
rect 6882 16496 6887 16552
rect 2773 16494 6887 16496
rect 2773 16491 2839 16494
rect 6821 16491 6887 16494
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 1485 16282 1551 16285
rect 0 16280 1551 16282
rect 0 16224 1490 16280
rect 1546 16224 1551 16280
rect 0 16222 1551 16224
rect 0 16192 480 16222
rect 1485 16219 1551 16222
rect 4797 16146 4863 16149
rect 7465 16146 7531 16149
rect 23657 16146 23723 16149
rect 4797 16144 7531 16146
rect 4797 16088 4802 16144
rect 4858 16088 7470 16144
rect 7526 16088 7531 16144
rect 4797 16086 7531 16088
rect 4797 16083 4863 16086
rect 7465 16083 7531 16086
rect 7606 16144 23723 16146
rect 7606 16088 23662 16144
rect 23718 16088 23723 16144
rect 7606 16086 23723 16088
rect 2497 16010 2563 16013
rect 3969 16010 4035 16013
rect 7606 16010 7666 16086
rect 23657 16083 23723 16086
rect 2497 16008 3802 16010
rect 2497 15952 2502 16008
rect 2558 15952 3802 16008
rect 2497 15950 3802 15952
rect 2497 15947 2563 15950
rect 2405 15874 2471 15877
rect 2773 15874 2839 15877
rect 2405 15872 2839 15874
rect 2405 15816 2410 15872
rect 2466 15816 2778 15872
rect 2834 15816 2839 15872
rect 2405 15814 2839 15816
rect 3742 15874 3802 15950
rect 3969 16008 7666 16010
rect 3969 15952 3974 16008
rect 4030 15952 7666 16008
rect 3969 15950 7666 15952
rect 9673 16010 9739 16013
rect 13997 16010 14063 16013
rect 9673 16008 14063 16010
rect 9673 15952 9678 16008
rect 9734 15952 14002 16008
rect 14058 15952 14063 16008
rect 9673 15950 14063 15952
rect 3969 15947 4035 15950
rect 9673 15947 9739 15950
rect 13997 15947 14063 15950
rect 6545 15874 6611 15877
rect 3742 15872 6611 15874
rect 3742 15816 6550 15872
rect 6606 15816 6611 15872
rect 3742 15814 6611 15816
rect 2405 15811 2471 15814
rect 2773 15811 2839 15814
rect 6545 15811 6611 15814
rect 10961 15874 11027 15877
rect 12433 15874 12499 15877
rect 10961 15872 12499 15874
rect 10961 15816 10966 15872
rect 11022 15816 12438 15872
rect 12494 15816 12499 15872
rect 10961 15814 12499 15816
rect 10961 15811 11027 15814
rect 12433 15811 12499 15814
rect 10277 15808 10597 15809
rect 0 15738 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 0 15678 7666 15738
rect 0 15648 480 15678
rect 1853 15602 1919 15605
rect 4153 15602 4219 15605
rect 1853 15600 4219 15602
rect 1853 15544 1858 15600
rect 1914 15544 4158 15600
rect 4214 15544 4219 15600
rect 1853 15542 4219 15544
rect 1853 15539 1919 15542
rect 4153 15539 4219 15542
rect 4705 15602 4771 15605
rect 7281 15602 7347 15605
rect 4705 15600 7347 15602
rect 4705 15544 4710 15600
rect 4766 15544 7286 15600
rect 7342 15544 7347 15600
rect 4705 15542 7347 15544
rect 7606 15602 7666 15678
rect 14825 15602 14891 15605
rect 7606 15600 14891 15602
rect 7606 15544 14830 15600
rect 14886 15544 14891 15600
rect 7606 15542 14891 15544
rect 4705 15539 4771 15542
rect 7281 15539 7347 15542
rect 14825 15539 14891 15542
rect 3877 15466 3943 15469
rect 4889 15466 4955 15469
rect 7741 15466 7807 15469
rect 3877 15464 7807 15466
rect 3877 15408 3882 15464
rect 3938 15408 4894 15464
rect 4950 15408 7746 15464
rect 7802 15408 7807 15464
rect 3877 15406 7807 15408
rect 3877 15403 3943 15406
rect 4889 15403 4955 15406
rect 7741 15403 7807 15406
rect 8201 15466 8267 15469
rect 12617 15466 12683 15469
rect 8201 15464 12683 15466
rect 8201 15408 8206 15464
rect 8262 15408 12622 15464
rect 12678 15408 12683 15464
rect 8201 15406 12683 15408
rect 8201 15403 8267 15406
rect 12617 15403 12683 15406
rect 1393 15330 1459 15333
rect 4797 15330 4863 15333
rect 1393 15328 4863 15330
rect 1393 15272 1398 15328
rect 1454 15272 4802 15328
rect 4858 15272 4863 15328
rect 1393 15270 4863 15272
rect 1393 15267 1459 15270
rect 4797 15267 4863 15270
rect 9765 15330 9831 15333
rect 12525 15330 12591 15333
rect 9765 15328 12591 15330
rect 9765 15272 9770 15328
rect 9826 15272 12530 15328
rect 12586 15272 12591 15328
rect 9765 15270 12591 15272
rect 9765 15267 9831 15270
rect 12525 15267 12591 15270
rect 5610 15264 5930 15265
rect 0 15194 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3969 15194 4035 15197
rect 0 15192 4035 15194
rect 0 15136 3974 15192
rect 4030 15136 4035 15192
rect 0 15134 4035 15136
rect 0 15104 480 15134
rect 3969 15131 4035 15134
rect 9489 15194 9555 15197
rect 13997 15194 14063 15197
rect 9489 15192 14063 15194
rect 9489 15136 9494 15192
rect 9550 15136 14002 15192
rect 14058 15136 14063 15192
rect 9489 15134 14063 15136
rect 9489 15131 9555 15134
rect 13997 15131 14063 15134
rect 1669 15058 1735 15061
rect 6545 15058 6611 15061
rect 1669 15056 6611 15058
rect 1669 15000 1674 15056
rect 1730 15000 6550 15056
rect 6606 15000 6611 15056
rect 1669 14998 6611 15000
rect 1669 14995 1735 14998
rect 6545 14995 6611 14998
rect 7097 15058 7163 15061
rect 13813 15058 13879 15061
rect 7097 15056 13879 15058
rect 7097 15000 7102 15056
rect 7158 15000 13818 15056
rect 13874 15000 13879 15056
rect 7097 14998 13879 15000
rect 7097 14995 7163 14998
rect 13813 14995 13879 14998
rect 2221 14922 2287 14925
rect 5441 14922 5507 14925
rect 11881 14922 11947 14925
rect 2221 14920 5507 14922
rect 2221 14864 2226 14920
rect 2282 14864 5446 14920
rect 5502 14864 5507 14920
rect 2221 14862 5507 14864
rect 2221 14859 2287 14862
rect 5441 14859 5507 14862
rect 5582 14920 11947 14922
rect 5582 14864 11886 14920
rect 11942 14864 11947 14920
rect 5582 14862 11947 14864
rect 1853 14786 1919 14789
rect 4797 14786 4863 14789
rect 5582 14786 5642 14862
rect 11881 14859 11947 14862
rect 1853 14784 4170 14786
rect 1853 14728 1858 14784
rect 1914 14728 4170 14784
rect 1853 14726 4170 14728
rect 1853 14723 1919 14726
rect 0 14650 480 14680
rect 3785 14650 3851 14653
rect 0 14648 3851 14650
rect 0 14592 3790 14648
rect 3846 14592 3851 14648
rect 0 14590 3851 14592
rect 4110 14650 4170 14726
rect 4797 14784 5642 14786
rect 4797 14728 4802 14784
rect 4858 14728 5642 14784
rect 4797 14726 5642 14728
rect 4797 14723 4863 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 5257 14650 5323 14653
rect 4110 14648 5323 14650
rect 4110 14592 5262 14648
rect 5318 14592 5323 14648
rect 4110 14590 5323 14592
rect 0 14560 480 14590
rect 3785 14587 3851 14590
rect 5257 14587 5323 14590
rect 4061 14514 4127 14517
rect 5717 14514 5783 14517
rect 4061 14512 5783 14514
rect 4061 14456 4066 14512
rect 4122 14456 5722 14512
rect 5778 14456 5783 14512
rect 4061 14454 5783 14456
rect 4061 14451 4127 14454
rect 5717 14451 5783 14454
rect 14825 14514 14891 14517
rect 23381 14514 23447 14517
rect 14825 14512 23447 14514
rect 14825 14456 14830 14512
rect 14886 14456 23386 14512
rect 23442 14456 23447 14512
rect 14825 14454 23447 14456
rect 14825 14451 14891 14454
rect 23381 14451 23447 14454
rect 6545 14242 6611 14245
rect 9305 14242 9371 14245
rect 6545 14240 9371 14242
rect 6545 14184 6550 14240
rect 6606 14184 9310 14240
rect 9366 14184 9371 14240
rect 6545 14182 9371 14184
rect 6545 14179 6611 14182
rect 9305 14179 9371 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 2865 14106 2931 14109
rect 2865 14104 5274 14106
rect 2865 14048 2870 14104
rect 2926 14048 5274 14104
rect 2865 14046 5274 14048
rect 2865 14043 2931 14046
rect 0 13970 480 14000
rect 2405 13970 2471 13973
rect 4981 13970 5047 13973
rect 0 13910 1410 13970
rect 0 13880 480 13910
rect 1350 13834 1410 13910
rect 2405 13968 5047 13970
rect 2405 13912 2410 13968
rect 2466 13912 4986 13968
rect 5042 13912 5047 13968
rect 2405 13910 5047 13912
rect 5214 13970 5274 14046
rect 6177 13970 6243 13973
rect 5214 13968 6243 13970
rect 5214 13912 6182 13968
rect 6238 13912 6243 13968
rect 5214 13910 6243 13912
rect 2405 13907 2471 13910
rect 4981 13907 5047 13910
rect 6177 13907 6243 13910
rect 23565 13970 23631 13973
rect 27520 13970 28000 14000
rect 23565 13968 28000 13970
rect 23565 13912 23570 13968
rect 23626 13912 28000 13968
rect 23565 13910 28000 13912
rect 23565 13907 23631 13910
rect 27520 13880 28000 13910
rect 3601 13834 3667 13837
rect 1350 13832 3667 13834
rect 1350 13776 3606 13832
rect 3662 13776 3667 13832
rect 1350 13774 3667 13776
rect 3601 13771 3667 13774
rect 4521 13698 4587 13701
rect 6821 13698 6887 13701
rect 4521 13696 6887 13698
rect 4521 13640 4526 13696
rect 4582 13640 6826 13696
rect 6882 13640 6887 13696
rect 4521 13638 6887 13640
rect 4521 13635 4587 13638
rect 6821 13635 6887 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 11329 13562 11395 13565
rect 14089 13562 14155 13565
rect 11329 13560 14155 13562
rect 11329 13504 11334 13560
rect 11390 13504 14094 13560
rect 14150 13504 14155 13560
rect 11329 13502 14155 13504
rect 11329 13499 11395 13502
rect 14089 13499 14155 13502
rect 0 13426 480 13456
rect 3877 13426 3943 13429
rect 0 13424 3943 13426
rect 0 13368 3882 13424
rect 3938 13368 3943 13424
rect 0 13366 3943 13368
rect 0 13336 480 13366
rect 3877 13363 3943 13366
rect 5257 13426 5323 13429
rect 12433 13426 12499 13429
rect 5257 13424 12499 13426
rect 5257 13368 5262 13424
rect 5318 13368 12438 13424
rect 12494 13368 12499 13424
rect 5257 13366 12499 13368
rect 5257 13363 5323 13366
rect 12433 13363 12499 13366
rect 9397 13290 9463 13293
rect 11145 13290 11211 13293
rect 9397 13288 11211 13290
rect 9397 13232 9402 13288
rect 9458 13232 11150 13288
rect 11206 13232 11211 13288
rect 9397 13230 11211 13232
rect 9397 13227 9463 13230
rect 11145 13227 11211 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12882 480 12912
rect 3325 12882 3391 12885
rect 0 12880 3391 12882
rect 0 12824 3330 12880
rect 3386 12824 3391 12880
rect 0 12822 3391 12824
rect 0 12792 480 12822
rect 3325 12819 3391 12822
rect 3785 12746 3851 12749
rect 22369 12746 22435 12749
rect 3785 12744 22435 12746
rect 3785 12688 3790 12744
rect 3846 12688 22374 12744
rect 22430 12688 22435 12744
rect 3785 12686 22435 12688
rect 3785 12683 3851 12686
rect 22369 12683 22435 12686
rect 2129 12610 2195 12613
rect 5993 12610 6059 12613
rect 2129 12608 6059 12610
rect 2129 12552 2134 12608
rect 2190 12552 5998 12608
rect 6054 12552 6059 12608
rect 2129 12550 6059 12552
rect 2129 12547 2195 12550
rect 5993 12547 6059 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 1945 12474 2011 12477
rect 2957 12474 3023 12477
rect 1945 12472 3023 12474
rect 1945 12416 1950 12472
rect 2006 12416 2962 12472
rect 3018 12416 3023 12472
rect 1945 12414 3023 12416
rect 1945 12411 2011 12414
rect 2957 12411 3023 12414
rect 3233 12474 3299 12477
rect 3785 12474 3851 12477
rect 3233 12472 3851 12474
rect 3233 12416 3238 12472
rect 3294 12416 3790 12472
rect 3846 12416 3851 12472
rect 3233 12414 3851 12416
rect 3233 12411 3299 12414
rect 3785 12411 3851 12414
rect 8753 12474 8819 12477
rect 8937 12474 9003 12477
rect 8753 12472 9003 12474
rect 8753 12416 8758 12472
rect 8814 12416 8942 12472
rect 8998 12416 9003 12472
rect 8753 12414 9003 12416
rect 8753 12411 8819 12414
rect 8937 12411 9003 12414
rect 0 12338 480 12368
rect 1761 12338 1827 12341
rect 3969 12338 4035 12341
rect 0 12278 1410 12338
rect 0 12248 480 12278
rect 1350 12202 1410 12278
rect 1761 12336 4035 12338
rect 1761 12280 1766 12336
rect 1822 12280 3974 12336
rect 4030 12280 4035 12336
rect 1761 12278 4035 12280
rect 1761 12275 1827 12278
rect 3969 12275 4035 12278
rect 4797 12338 4863 12341
rect 7925 12338 7991 12341
rect 4797 12336 7991 12338
rect 4797 12280 4802 12336
rect 4858 12280 7930 12336
rect 7986 12280 7991 12336
rect 4797 12278 7991 12280
rect 4797 12275 4863 12278
rect 7925 12275 7991 12278
rect 12709 12338 12775 12341
rect 23565 12338 23631 12341
rect 12709 12336 23631 12338
rect 12709 12280 12714 12336
rect 12770 12280 23570 12336
rect 23626 12280 23631 12336
rect 12709 12278 23631 12280
rect 12709 12275 12775 12278
rect 23565 12275 23631 12278
rect 3417 12202 3483 12205
rect 1350 12200 3483 12202
rect 1350 12144 3422 12200
rect 3478 12144 3483 12200
rect 1350 12142 3483 12144
rect 3417 12139 3483 12142
rect 4337 12202 4403 12205
rect 12617 12202 12683 12205
rect 4337 12200 12683 12202
rect 4337 12144 4342 12200
rect 4398 12144 12622 12200
rect 12678 12144 12683 12200
rect 4337 12142 12683 12144
rect 4337 12139 4403 12142
rect 12617 12139 12683 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 12341 11930 12407 11933
rect 13813 11930 13879 11933
rect 12341 11928 13879 11930
rect 12341 11872 12346 11928
rect 12402 11872 13818 11928
rect 13874 11872 13879 11928
rect 12341 11870 13879 11872
rect 12341 11867 12407 11870
rect 13813 11867 13879 11870
rect 0 11794 480 11824
rect 2957 11794 3023 11797
rect 6085 11794 6151 11797
rect 0 11734 2744 11794
rect 0 11704 480 11734
rect 2684 11692 2744 11734
rect 2957 11792 6151 11794
rect 2957 11736 2962 11792
rect 3018 11736 6090 11792
rect 6146 11736 6151 11792
rect 2957 11734 6151 11736
rect 2957 11731 3023 11734
rect 6085 11731 6151 11734
rect 2684 11658 2836 11692
rect 3233 11658 3299 11661
rect 2684 11656 3299 11658
rect 2684 11632 3238 11656
rect 2776 11600 3238 11632
rect 3294 11600 3299 11656
rect 2776 11598 3299 11600
rect 3233 11595 3299 11598
rect 3601 11658 3667 11661
rect 21817 11658 21883 11661
rect 3601 11656 21883 11658
rect 3601 11600 3606 11656
rect 3662 11600 21822 11656
rect 21878 11600 21883 11656
rect 3601 11598 21883 11600
rect 3601 11595 3667 11598
rect 21817 11595 21883 11598
rect 4153 11522 4219 11525
rect 6913 11522 6979 11525
rect 4153 11520 6979 11522
rect 4153 11464 4158 11520
rect 4214 11464 6918 11520
rect 6974 11464 6979 11520
rect 4153 11462 6979 11464
rect 4153 11459 4219 11462
rect 6913 11459 6979 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3969 11386 4035 11389
rect 6821 11386 6887 11389
rect 3969 11384 6887 11386
rect 3969 11328 3974 11384
rect 4030 11328 6826 11384
rect 6882 11328 6887 11384
rect 3969 11326 6887 11328
rect 3969 11323 4035 11326
rect 6821 11323 6887 11326
rect 4153 11250 4219 11253
rect 11053 11250 11119 11253
rect 4153 11248 11119 11250
rect 4153 11192 4158 11248
rect 4214 11192 11058 11248
rect 11114 11192 11119 11248
rect 4153 11190 11119 11192
rect 4153 11187 4219 11190
rect 11053 11187 11119 11190
rect 0 11114 480 11144
rect 5809 11114 5875 11117
rect 13261 11114 13327 11117
rect 0 11054 5458 11114
rect 0 11024 480 11054
rect 5398 10706 5458 11054
rect 5809 11112 13327 11114
rect 5809 11056 5814 11112
rect 5870 11056 13266 11112
rect 13322 11056 13327 11112
rect 5809 11054 13327 11056
rect 5809 11051 5875 11054
rect 13261 11051 13327 11054
rect 22001 11114 22067 11117
rect 23657 11114 23723 11117
rect 22001 11112 23723 11114
rect 22001 11056 22006 11112
rect 22062 11056 23662 11112
rect 23718 11056 23723 11112
rect 22001 11054 23723 11056
rect 22001 11051 22067 11054
rect 23657 11051 23723 11054
rect 6361 10978 6427 10981
rect 11789 10978 11855 10981
rect 6361 10976 11855 10978
rect 6361 10920 6366 10976
rect 6422 10920 11794 10976
rect 11850 10920 11855 10976
rect 6361 10918 11855 10920
rect 6361 10915 6427 10918
rect 11789 10915 11855 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 15745 10706 15811 10709
rect 5398 10704 15811 10706
rect 5398 10648 15750 10704
rect 15806 10648 15811 10704
rect 5398 10646 15811 10648
rect 15745 10643 15811 10646
rect 0 10570 480 10600
rect 5073 10570 5139 10573
rect 7097 10570 7163 10573
rect 0 10510 2744 10570
rect 0 10480 480 10510
rect 2684 10468 2744 10510
rect 5073 10568 7163 10570
rect 5073 10512 5078 10568
rect 5134 10512 7102 10568
rect 7158 10512 7163 10568
rect 5073 10510 7163 10512
rect 5073 10507 5139 10510
rect 7097 10507 7163 10510
rect 8017 10570 8083 10573
rect 12801 10570 12867 10573
rect 8017 10568 12867 10570
rect 8017 10512 8022 10568
rect 8078 10512 12806 10568
rect 12862 10512 12867 10568
rect 8017 10510 12867 10512
rect 8017 10507 8083 10510
rect 12801 10507 12867 10510
rect 2684 10434 2836 10468
rect 6637 10434 6703 10437
rect 2684 10432 6703 10434
rect 2684 10408 6642 10432
rect 2776 10376 6642 10408
rect 6698 10376 6703 10432
rect 2776 10374 6703 10376
rect 6637 10371 6703 10374
rect 10685 10434 10751 10437
rect 12893 10434 12959 10437
rect 10685 10432 12959 10434
rect 10685 10376 10690 10432
rect 10746 10376 12898 10432
rect 12954 10376 12959 10432
rect 10685 10374 12959 10376
rect 10685 10371 10751 10374
rect 12893 10371 12959 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 4889 10298 4955 10301
rect 7925 10298 7991 10301
rect 4889 10296 7991 10298
rect 4889 10240 4894 10296
rect 4950 10240 7930 10296
rect 7986 10240 7991 10296
rect 4889 10238 7991 10240
rect 4889 10235 4955 10238
rect 7925 10235 7991 10238
rect 3877 10162 3943 10165
rect 11513 10162 11579 10165
rect 3877 10160 11579 10162
rect 3877 10104 3882 10160
rect 3938 10104 11518 10160
rect 11574 10104 11579 10160
rect 3877 10102 11579 10104
rect 3877 10099 3943 10102
rect 11513 10099 11579 10102
rect 0 10026 480 10056
rect 3969 10026 4035 10029
rect 10777 10026 10843 10029
rect 19333 10026 19399 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 480 9966
rect 3969 9963 4035 9966
rect 5398 9966 10242 10026
rect 3325 9890 3391 9893
rect 5398 9890 5458 9966
rect 3325 9888 5458 9890
rect 3325 9832 3330 9888
rect 3386 9832 5458 9888
rect 3325 9830 5458 9832
rect 3325 9827 3391 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 3141 9754 3207 9757
rect 10182 9754 10242 9966
rect 10777 10024 19399 10026
rect 10777 9968 10782 10024
rect 10838 9968 19338 10024
rect 19394 9968 19399 10024
rect 10777 9966 19399 9968
rect 10777 9963 10843 9966
rect 19333 9963 19399 9966
rect 10317 9890 10383 9893
rect 12801 9890 12867 9893
rect 10317 9888 12867 9890
rect 10317 9832 10322 9888
rect 10378 9832 12806 9888
rect 12862 9832 12867 9888
rect 10317 9830 12867 9832
rect 10317 9827 10383 9830
rect 12801 9827 12867 9830
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 11789 9754 11855 9757
rect 3141 9752 5458 9754
rect 3141 9696 3146 9752
rect 3202 9696 5458 9752
rect 3141 9694 5458 9696
rect 10182 9752 11855 9754
rect 10182 9696 11794 9752
rect 11850 9696 11855 9752
rect 10182 9694 11855 9696
rect 3141 9691 3207 9694
rect 5398 9618 5458 9694
rect 11789 9691 11855 9694
rect 12341 9652 12407 9655
rect 12206 9650 12407 9652
rect 5625 9618 5691 9621
rect 5398 9616 5691 9618
rect 5398 9560 5630 9616
rect 5686 9560 5691 9616
rect 5398 9558 5691 9560
rect 5625 9555 5691 9558
rect 8017 9618 8083 9621
rect 12206 9618 12346 9650
rect 8017 9616 12346 9618
rect 8017 9560 8022 9616
rect 8078 9594 12346 9616
rect 12402 9594 12407 9650
rect 8078 9592 12407 9594
rect 8078 9560 12266 9592
rect 12341 9589 12407 9592
rect 8017 9558 12266 9560
rect 8017 9555 8083 9558
rect 0 9482 480 9512
rect 3877 9482 3943 9485
rect 0 9480 3943 9482
rect 0 9424 3882 9480
rect 3938 9424 3943 9480
rect 0 9422 3943 9424
rect 0 9392 480 9422
rect 3877 9419 3943 9422
rect 7097 9482 7163 9485
rect 10685 9482 10751 9485
rect 12985 9482 13051 9485
rect 7097 9480 13051 9482
rect 7097 9424 7102 9480
rect 7158 9424 10690 9480
rect 10746 9424 12990 9480
rect 13046 9424 13051 9480
rect 7097 9422 13051 9424
rect 7097 9419 7163 9422
rect 10685 9419 10751 9422
rect 12985 9419 13051 9422
rect 1853 9346 1919 9349
rect 4245 9346 4311 9349
rect 1853 9344 4311 9346
rect 1853 9288 1858 9344
rect 1914 9288 4250 9344
rect 4306 9288 4311 9344
rect 1853 9286 4311 9288
rect 1853 9283 1919 9286
rect 4245 9283 4311 9286
rect 13537 9346 13603 9349
rect 16665 9346 16731 9349
rect 13537 9344 16731 9346
rect 13537 9288 13542 9344
rect 13598 9288 16670 9344
rect 16726 9288 16731 9344
rect 13537 9286 16731 9288
rect 13537 9283 13603 9286
rect 16665 9283 16731 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2589 9210 2655 9213
rect 4981 9210 5047 9213
rect 2589 9208 5047 9210
rect 2589 9152 2594 9208
rect 2650 9152 4986 9208
rect 5042 9152 5047 9208
rect 2589 9150 5047 9152
rect 2589 9147 2655 9150
rect 4981 9147 5047 9150
rect 3969 9074 4035 9077
rect 10501 9074 10567 9077
rect 3969 9072 10567 9074
rect 3969 9016 3974 9072
rect 4030 9016 10506 9072
rect 10562 9016 10567 9072
rect 3969 9014 10567 9016
rect 3969 9011 4035 9014
rect 10501 9011 10567 9014
rect 13721 9074 13787 9077
rect 19977 9074 20043 9077
rect 13721 9072 20043 9074
rect 13721 9016 13726 9072
rect 13782 9016 19982 9072
rect 20038 9016 20043 9072
rect 13721 9014 20043 9016
rect 13721 9011 13787 9014
rect 19977 9011 20043 9014
rect 0 8938 480 8968
rect 2497 8938 2563 8941
rect 0 8936 2563 8938
rect 0 8880 2502 8936
rect 2558 8880 2563 8936
rect 0 8878 2563 8880
rect 0 8848 480 8878
rect 2497 8875 2563 8878
rect 3509 8938 3575 8941
rect 7649 8938 7715 8941
rect 3509 8936 7715 8938
rect 3509 8880 3514 8936
rect 3570 8880 7654 8936
rect 7710 8880 7715 8936
rect 3509 8878 7715 8880
rect 3509 8875 3575 8878
rect 7649 8875 7715 8878
rect 10133 8938 10199 8941
rect 18229 8938 18295 8941
rect 10133 8936 18295 8938
rect 10133 8880 10138 8936
rect 10194 8880 18234 8936
rect 18290 8880 18295 8936
rect 10133 8878 18295 8880
rect 10133 8875 10199 8878
rect 18229 8875 18295 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 3693 8530 3759 8533
rect 5533 8530 5599 8533
rect 3693 8528 5599 8530
rect 3693 8472 3698 8528
rect 3754 8472 5538 8528
rect 5594 8472 5599 8528
rect 3693 8470 5599 8472
rect 3693 8467 3759 8470
rect 5533 8467 5599 8470
rect 8569 8530 8635 8533
rect 13721 8530 13787 8533
rect 8569 8528 13787 8530
rect 8569 8472 8574 8528
rect 8630 8472 13726 8528
rect 13782 8472 13787 8528
rect 8569 8470 13787 8472
rect 8569 8467 8635 8470
rect 13721 8467 13787 8470
rect 13997 8530 14063 8533
rect 20253 8530 20319 8533
rect 13997 8528 20319 8530
rect 13997 8472 14002 8528
rect 14058 8472 20258 8528
rect 20314 8472 20319 8528
rect 13997 8470 20319 8472
rect 13997 8467 14063 8470
rect 20253 8467 20319 8470
rect 3785 8394 3851 8397
rect 3969 8394 4035 8397
rect 6545 8394 6611 8397
rect 3785 8392 6611 8394
rect 3785 8336 3790 8392
rect 3846 8336 3974 8392
rect 4030 8336 6550 8392
rect 6606 8336 6611 8392
rect 3785 8334 6611 8336
rect 3785 8331 3851 8334
rect 3969 8331 4035 8334
rect 6545 8331 6611 8334
rect 10961 8394 11027 8397
rect 11697 8394 11763 8397
rect 10961 8392 11763 8394
rect 10961 8336 10966 8392
rect 11022 8336 11702 8392
rect 11758 8336 11763 8392
rect 10961 8334 11763 8336
rect 10961 8331 11027 8334
rect 11697 8331 11763 8334
rect 14457 8394 14523 8397
rect 18137 8394 18203 8397
rect 14457 8392 18203 8394
rect 14457 8336 14462 8392
rect 14518 8336 18142 8392
rect 18198 8336 18203 8392
rect 14457 8334 18203 8336
rect 14457 8331 14523 8334
rect 18137 8331 18203 8334
rect 0 8258 480 8288
rect 0 8198 10058 8258
rect 0 8168 480 8198
rect 2405 8122 2471 8125
rect 4613 8122 4679 8125
rect 2405 8120 4679 8122
rect 2405 8064 2410 8120
rect 2466 8064 4618 8120
rect 4674 8064 4679 8120
rect 2405 8062 4679 8064
rect 2405 8059 2471 8062
rect 4613 8059 4679 8062
rect 9998 7986 10058 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 10961 7986 11027 7989
rect 9998 7984 11027 7986
rect 9998 7928 10966 7984
rect 11022 7928 11027 7984
rect 9998 7926 11027 7928
rect 10961 7923 11027 7926
rect 8109 7850 8175 7853
rect 5398 7848 8175 7850
rect 5398 7792 8114 7848
rect 8170 7792 8175 7848
rect 5398 7790 8175 7792
rect 0 7714 480 7744
rect 5398 7714 5458 7790
rect 8109 7787 8175 7790
rect 10726 7788 10732 7852
rect 10796 7850 10802 7852
rect 10869 7850 10935 7853
rect 19057 7850 19123 7853
rect 10796 7848 10935 7850
rect 10796 7792 10874 7848
rect 10930 7792 10935 7848
rect 10796 7790 10935 7792
rect 10796 7788 10802 7790
rect 10869 7787 10935 7790
rect 14782 7848 19123 7850
rect 14782 7792 19062 7848
rect 19118 7792 19123 7848
rect 14782 7790 19123 7792
rect 0 7654 5458 7714
rect 7741 7714 7807 7717
rect 9857 7714 9923 7717
rect 7741 7712 9923 7714
rect 7741 7656 7746 7712
rect 7802 7656 9862 7712
rect 9918 7656 9923 7712
rect 7741 7654 9923 7656
rect 0 7624 480 7654
rect 7741 7651 7807 7654
rect 9857 7651 9923 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 1669 7578 1735 7581
rect 4153 7578 4219 7581
rect 1669 7576 4219 7578
rect 1669 7520 1674 7576
rect 1730 7520 4158 7576
rect 4214 7520 4219 7576
rect 1669 7518 4219 7520
rect 1669 7515 1735 7518
rect 4153 7515 4219 7518
rect 6637 7578 6703 7581
rect 14782 7578 14842 7790
rect 19057 7787 19123 7790
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 6637 7576 14842 7578
rect 6637 7520 6642 7576
rect 6698 7520 14842 7576
rect 6637 7518 14842 7520
rect 6637 7515 6703 7518
rect 1393 7442 1459 7445
rect 6913 7442 6979 7445
rect 1393 7440 6979 7442
rect 1393 7384 1398 7440
rect 1454 7384 6918 7440
rect 6974 7384 6979 7440
rect 1393 7382 6979 7384
rect 1393 7379 1459 7382
rect 6913 7379 6979 7382
rect 13629 7442 13695 7445
rect 19701 7442 19767 7445
rect 13629 7440 19767 7442
rect 13629 7384 13634 7440
rect 13690 7384 19706 7440
rect 19762 7384 19767 7440
rect 13629 7382 19767 7384
rect 13629 7379 13695 7382
rect 19701 7379 19767 7382
rect 3417 7306 3483 7309
rect 16205 7306 16271 7309
rect 3417 7304 16271 7306
rect 3417 7248 3422 7304
rect 3478 7248 16210 7304
rect 16266 7248 16271 7304
rect 3417 7246 16271 7248
rect 3417 7243 3483 7246
rect 16205 7243 16271 7246
rect 0 7170 480 7200
rect 5349 7170 5415 7173
rect 0 7168 5415 7170
rect 0 7112 5354 7168
rect 5410 7112 5415 7168
rect 0 7110 5415 7112
rect 0 7080 480 7110
rect 5349 7107 5415 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2313 6898 2379 6901
rect 5257 6898 5323 6901
rect 19517 6898 19583 6901
rect 2313 6896 19583 6898
rect 2313 6840 2318 6896
rect 2374 6840 5262 6896
rect 5318 6840 19522 6896
rect 19578 6840 19583 6896
rect 2313 6838 19583 6840
rect 2313 6835 2379 6838
rect 5257 6835 5323 6838
rect 19517 6835 19583 6838
rect 3509 6762 3575 6765
rect 11513 6762 11579 6765
rect 3509 6760 11579 6762
rect 3509 6704 3514 6760
rect 3570 6704 11518 6760
rect 11574 6704 11579 6760
rect 3509 6702 11579 6704
rect 3509 6699 3575 6702
rect 11513 6699 11579 6702
rect 12433 6762 12499 6765
rect 15377 6762 15443 6765
rect 12433 6760 15443 6762
rect 12433 6704 12438 6760
rect 12494 6704 15382 6760
rect 15438 6704 15443 6760
rect 12433 6702 15443 6704
rect 12433 6699 12499 6702
rect 15377 6699 15443 6702
rect 0 6626 480 6656
rect 4245 6626 4311 6629
rect 0 6624 4311 6626
rect 0 6568 4250 6624
rect 4306 6568 4311 6624
rect 0 6566 4311 6568
rect 0 6536 480 6566
rect 4245 6563 4311 6566
rect 9765 6626 9831 6629
rect 9765 6624 14842 6626
rect 9765 6568 9770 6624
rect 9826 6568 14842 6624
rect 9765 6566 14842 6568
rect 9765 6563 9831 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 10501 6354 10567 6357
rect 12893 6354 12959 6357
rect 10501 6352 12959 6354
rect 10501 6296 10506 6352
rect 10562 6296 12898 6352
rect 12954 6296 12959 6352
rect 10501 6294 12959 6296
rect 14782 6354 14842 6566
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 15285 6354 15351 6357
rect 14782 6352 15351 6354
rect 14782 6296 15290 6352
rect 15346 6296 15351 6352
rect 14782 6294 15351 6296
rect 10501 6291 10567 6294
rect 12893 6291 12959 6294
rect 15285 6291 15351 6294
rect 1945 6218 2011 6221
rect 11053 6218 11119 6221
rect 1945 6216 11119 6218
rect 1945 6160 1950 6216
rect 2006 6160 11058 6216
rect 11114 6160 11119 6216
rect 1945 6158 11119 6160
rect 1945 6155 2011 6158
rect 11053 6155 11119 6158
rect 11329 6218 11395 6221
rect 18045 6218 18111 6221
rect 11329 6216 18111 6218
rect 11329 6160 11334 6216
rect 11390 6160 18050 6216
rect 18106 6160 18111 6216
rect 11329 6158 18111 6160
rect 11329 6155 11395 6158
rect 18045 6155 18111 6158
rect 0 6082 480 6112
rect 1853 6082 1919 6085
rect 0 6080 1919 6082
rect 0 6024 1858 6080
rect 1914 6024 1919 6080
rect 0 6022 1919 6024
rect 0 5992 480 6022
rect 1853 6019 1919 6022
rect 6453 6082 6519 6085
rect 9857 6082 9923 6085
rect 6453 6080 9923 6082
rect 6453 6024 6458 6080
rect 6514 6024 9862 6080
rect 9918 6024 9923 6080
rect 6453 6022 9923 6024
rect 6453 6019 6519 6022
rect 9857 6019 9923 6022
rect 13629 6082 13695 6085
rect 16389 6082 16455 6085
rect 13629 6080 16455 6082
rect 13629 6024 13634 6080
rect 13690 6024 16394 6080
rect 16450 6024 16455 6080
rect 13629 6022 16455 6024
rect 13629 6019 13695 6022
rect 16389 6019 16455 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 13997 5946 14063 5949
rect 16665 5946 16731 5949
rect 13997 5944 16731 5946
rect 13997 5888 14002 5944
rect 14058 5888 16670 5944
rect 16726 5888 16731 5944
rect 13997 5886 16731 5888
rect 13997 5883 14063 5886
rect 16665 5883 16731 5886
rect 8569 5810 8635 5813
rect 15469 5810 15535 5813
rect 8569 5808 15535 5810
rect 8569 5752 8574 5808
rect 8630 5752 15474 5808
rect 15530 5752 15535 5808
rect 8569 5750 15535 5752
rect 8569 5747 8635 5750
rect 15469 5747 15535 5750
rect 3877 5674 3943 5677
rect 7373 5674 7439 5677
rect 8293 5674 8359 5677
rect 3877 5672 8359 5674
rect 3877 5616 3882 5672
rect 3938 5616 7378 5672
rect 7434 5616 8298 5672
rect 8354 5616 8359 5672
rect 3877 5614 8359 5616
rect 3877 5611 3943 5614
rect 7373 5611 7439 5614
rect 8293 5611 8359 5614
rect 11237 5674 11303 5677
rect 15469 5674 15535 5677
rect 11237 5672 15535 5674
rect 11237 5616 11242 5672
rect 11298 5616 15474 5672
rect 15530 5616 15535 5672
rect 11237 5614 15535 5616
rect 11237 5611 11303 5614
rect 15469 5611 15535 5614
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 11513 5402 11579 5405
rect 14733 5402 14799 5405
rect 0 5342 5458 5402
rect 0 5312 480 5342
rect 5398 5266 5458 5342
rect 11513 5400 14799 5402
rect 11513 5344 11518 5400
rect 11574 5344 14738 5400
rect 14794 5344 14799 5400
rect 11513 5342 14799 5344
rect 11513 5339 11579 5342
rect 14733 5339 14799 5342
rect 7741 5266 7807 5269
rect 5398 5264 7807 5266
rect 5398 5208 7746 5264
rect 7802 5208 7807 5264
rect 5398 5206 7807 5208
rect 7741 5203 7807 5206
rect 5073 5130 5139 5133
rect 7097 5130 7163 5133
rect 5073 5128 7163 5130
rect 5073 5072 5078 5128
rect 5134 5072 7102 5128
rect 7158 5072 7163 5128
rect 5073 5070 7163 5072
rect 5073 5067 5139 5070
rect 7097 5067 7163 5070
rect 8477 5130 8543 5133
rect 17769 5130 17835 5133
rect 8477 5128 17835 5130
rect 8477 5072 8482 5128
rect 8538 5072 17774 5128
rect 17830 5072 17835 5128
rect 8477 5070 17835 5072
rect 8477 5067 8543 5070
rect 17769 5067 17835 5070
rect 2497 4994 2563 4997
rect 8150 4994 8156 4996
rect 2497 4992 8156 4994
rect 2497 4936 2502 4992
rect 2558 4936 8156 4992
rect 2497 4934 8156 4936
rect 2497 4931 2563 4934
rect 8150 4932 8156 4934
rect 8220 4932 8226 4996
rect 11053 4994 11119 4997
rect 15193 4994 15259 4997
rect 11053 4992 15259 4994
rect 11053 4936 11058 4992
rect 11114 4936 15198 4992
rect 15254 4936 15259 4992
rect 11053 4934 15259 4936
rect 11053 4931 11119 4934
rect 15193 4931 15259 4934
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3601 4858 3667 4861
rect 0 4856 3667 4858
rect 0 4800 3606 4856
rect 3662 4800 3667 4856
rect 0 4798 3667 4800
rect 0 4768 480 4798
rect 3601 4795 3667 4798
rect 10869 4858 10935 4861
rect 13905 4858 13971 4861
rect 10869 4856 13971 4858
rect 10869 4800 10874 4856
rect 10930 4800 13910 4856
rect 13966 4800 13971 4856
rect 10869 4798 13971 4800
rect 10869 4795 10935 4798
rect 13905 4795 13971 4798
rect 8150 4660 8156 4724
rect 8220 4722 8226 4724
rect 24117 4722 24183 4725
rect 27520 4722 28000 4752
rect 8220 4662 9506 4722
rect 8220 4660 8226 4662
rect 3325 4586 3391 4589
rect 8845 4586 8911 4589
rect 3325 4584 7850 4586
rect 3325 4528 3330 4584
rect 3386 4552 7850 4584
rect 7974 4584 8911 4586
rect 7974 4552 8850 4584
rect 3386 4528 8850 4552
rect 8906 4528 8911 4584
rect 3325 4526 8911 4528
rect 9446 4586 9506 4662
rect 24117 4720 28000 4722
rect 24117 4664 24122 4720
rect 24178 4664 28000 4720
rect 24117 4662 28000 4664
rect 24117 4659 24183 4662
rect 27520 4632 28000 4662
rect 9581 4586 9647 4589
rect 9446 4584 9647 4586
rect 9446 4528 9586 4584
rect 9642 4528 9647 4584
rect 9446 4526 9647 4528
rect 3325 4523 3391 4526
rect 7790 4492 8034 4526
rect 8845 4523 8911 4526
rect 9581 4523 9647 4526
rect 12985 4586 13051 4589
rect 19885 4586 19951 4589
rect 12985 4584 19951 4586
rect 12985 4528 12990 4584
rect 13046 4528 19890 4584
rect 19946 4528 19951 4584
rect 12985 4526 19951 4528
rect 12985 4523 13051 4526
rect 19885 4523 19951 4526
rect 5610 4384 5930 4385
rect 0 4314 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 2957 4314 3023 4317
rect 0 4312 3023 4314
rect 0 4256 2962 4312
rect 3018 4256 3023 4312
rect 0 4254 3023 4256
rect 0 4224 480 4254
rect 2957 4251 3023 4254
rect 15653 4314 15719 4317
rect 20897 4314 20963 4317
rect 15653 4312 20963 4314
rect 15653 4256 15658 4312
rect 15714 4256 20902 4312
rect 20958 4256 20963 4312
rect 15653 4254 20963 4256
rect 15653 4251 15719 4254
rect 20897 4251 20963 4254
rect 3601 4178 3667 4181
rect 24025 4178 24091 4181
rect 3601 4176 24091 4178
rect 3601 4120 3606 4176
rect 3662 4120 24030 4176
rect 24086 4120 24091 4176
rect 3601 4118 24091 4120
rect 3601 4115 3667 4118
rect 24025 4115 24091 4118
rect 3049 4042 3115 4045
rect 4521 4042 4587 4045
rect 3049 4040 4587 4042
rect 3049 3984 3054 4040
rect 3110 3984 4526 4040
rect 4582 3984 4587 4040
rect 3049 3982 4587 3984
rect 3049 3979 3115 3982
rect 4521 3979 4587 3982
rect 8293 4042 8359 4045
rect 12157 4042 12223 4045
rect 8293 4040 12223 4042
rect 8293 3984 8298 4040
rect 8354 3984 12162 4040
rect 12218 3984 12223 4040
rect 8293 3982 12223 3984
rect 8293 3979 8359 3982
rect 12157 3979 12223 3982
rect 18413 4042 18479 4045
rect 22277 4042 22343 4045
rect 18413 4040 22343 4042
rect 18413 3984 18418 4040
rect 18474 3984 22282 4040
rect 22338 3984 22343 4040
rect 18413 3982 22343 3984
rect 18413 3979 18479 3982
rect 22277 3979 22343 3982
rect 2681 3906 2747 3909
rect 5349 3906 5415 3909
rect 2681 3904 5415 3906
rect 2681 3848 2686 3904
rect 2742 3848 5354 3904
rect 5410 3848 5415 3904
rect 2681 3846 5415 3848
rect 2681 3843 2747 3846
rect 5349 3843 5415 3846
rect 11329 3906 11395 3909
rect 18137 3906 18203 3909
rect 11329 3904 18203 3906
rect 11329 3848 11334 3904
rect 11390 3848 18142 3904
rect 18198 3848 18203 3904
rect 11329 3846 18203 3848
rect 11329 3843 11395 3846
rect 18137 3843 18203 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2405 3770 2471 3773
rect 4981 3770 5047 3773
rect 17401 3770 17467 3773
rect 0 3710 1410 3770
rect 0 3680 480 3710
rect 1350 3634 1410 3710
rect 2405 3768 5047 3770
rect 2405 3712 2410 3768
rect 2466 3712 4986 3768
rect 5042 3712 5047 3768
rect 2405 3710 5047 3712
rect 2405 3707 2471 3710
rect 4981 3707 5047 3710
rect 14092 3768 17467 3770
rect 14092 3712 17406 3768
rect 17462 3712 17467 3768
rect 14092 3710 17467 3712
rect 3969 3634 4035 3637
rect 1350 3632 4035 3634
rect 1350 3576 3974 3632
rect 4030 3576 4035 3632
rect 1350 3574 4035 3576
rect 3969 3571 4035 3574
rect 9029 3634 9095 3637
rect 11145 3634 11211 3637
rect 9029 3632 11211 3634
rect 9029 3576 9034 3632
rect 9090 3576 11150 3632
rect 11206 3576 11211 3632
rect 9029 3574 11211 3576
rect 9029 3571 9095 3574
rect 11145 3571 11211 3574
rect 11881 3634 11947 3637
rect 14092 3634 14152 3710
rect 17401 3707 17467 3710
rect 11881 3632 14152 3634
rect 11881 3576 11886 3632
rect 11942 3576 14152 3632
rect 11881 3574 14152 3576
rect 14273 3634 14339 3637
rect 17125 3634 17191 3637
rect 14273 3632 17191 3634
rect 14273 3576 14278 3632
rect 14334 3576 17130 3632
rect 17186 3576 17191 3632
rect 14273 3574 17191 3576
rect 11881 3571 11947 3574
rect 14273 3571 14339 3574
rect 17125 3571 17191 3574
rect 3049 3498 3115 3501
rect 8937 3498 9003 3501
rect 9765 3498 9831 3501
rect 3049 3496 9831 3498
rect 3049 3440 3054 3496
rect 3110 3440 8942 3496
rect 8998 3440 9770 3496
rect 9826 3440 9831 3496
rect 3049 3438 9831 3440
rect 3049 3435 3115 3438
rect 8937 3435 9003 3438
rect 9765 3435 9831 3438
rect 10133 3498 10199 3501
rect 15561 3498 15627 3501
rect 10133 3496 15627 3498
rect 10133 3440 10138 3496
rect 10194 3440 15566 3496
rect 15622 3440 15627 3496
rect 10133 3438 15627 3440
rect 10133 3435 10199 3438
rect 15561 3435 15627 3438
rect 20345 3498 20411 3501
rect 23565 3498 23631 3501
rect 20345 3496 23631 3498
rect 20345 3440 20350 3496
rect 20406 3440 23570 3496
rect 23626 3440 23631 3496
rect 20345 3438 23631 3440
rect 20345 3435 20411 3438
rect 23565 3435 23631 3438
rect 1669 3362 1735 3365
rect 4245 3362 4311 3365
rect 1669 3360 4311 3362
rect 1669 3304 1674 3360
rect 1730 3304 4250 3360
rect 4306 3304 4311 3360
rect 1669 3302 4311 3304
rect 1669 3299 1735 3302
rect 4245 3299 4311 3302
rect 8017 3362 8083 3365
rect 11789 3362 11855 3365
rect 8017 3360 11855 3362
rect 8017 3304 8022 3360
rect 8078 3304 11794 3360
rect 11850 3304 11855 3360
rect 8017 3302 11855 3304
rect 8017 3299 8083 3302
rect 11789 3299 11855 3302
rect 18045 3362 18111 3365
rect 20805 3362 20871 3365
rect 18045 3360 20871 3362
rect 18045 3304 18050 3360
rect 18106 3304 20810 3360
rect 20866 3304 20871 3360
rect 18045 3302 20871 3304
rect 18045 3299 18111 3302
rect 20805 3299 20871 3302
rect 21633 3362 21699 3365
rect 22553 3362 22619 3365
rect 21633 3360 22619 3362
rect 21633 3304 21638 3360
rect 21694 3304 22558 3360
rect 22614 3304 22619 3360
rect 21633 3302 22619 3304
rect 21633 3299 21699 3302
rect 22553 3299 22619 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 3693 3226 3759 3229
rect 13905 3226 13971 3229
rect 0 3224 3759 3226
rect 0 3168 3698 3224
rect 3754 3168 3759 3224
rect 0 3166 3759 3168
rect 0 3136 480 3166
rect 3693 3163 3759 3166
rect 8756 3224 13971 3226
rect 8756 3168 13910 3224
rect 13966 3168 13971 3224
rect 8756 3166 13971 3168
rect 5165 3090 5231 3093
rect 8756 3090 8816 3166
rect 13905 3163 13971 3166
rect 18229 3226 18295 3229
rect 20713 3226 20779 3229
rect 18229 3224 20779 3226
rect 18229 3168 18234 3224
rect 18290 3168 20718 3224
rect 20774 3168 20779 3224
rect 18229 3166 20779 3168
rect 18229 3163 18295 3166
rect 20713 3163 20779 3166
rect 5165 3088 8816 3090
rect 5165 3032 5170 3088
rect 5226 3032 8816 3088
rect 5165 3030 8816 3032
rect 8937 3090 9003 3093
rect 11053 3090 11119 3093
rect 8937 3088 11119 3090
rect 8937 3032 8942 3088
rect 8998 3032 11058 3088
rect 11114 3032 11119 3088
rect 8937 3030 11119 3032
rect 5165 3027 5231 3030
rect 8937 3027 9003 3030
rect 11053 3027 11119 3030
rect 11421 3090 11487 3093
rect 17677 3090 17743 3093
rect 11421 3088 17743 3090
rect 11421 3032 11426 3088
rect 11482 3032 17682 3088
rect 17738 3032 17743 3088
rect 11421 3030 17743 3032
rect 11421 3027 11487 3030
rect 17677 3027 17743 3030
rect 19609 3090 19675 3093
rect 22185 3090 22251 3093
rect 19609 3088 22251 3090
rect 19609 3032 19614 3088
rect 19670 3032 22190 3088
rect 22246 3032 22251 3088
rect 19609 3030 22251 3032
rect 19609 3027 19675 3030
rect 22185 3027 22251 3030
rect 24209 3090 24275 3093
rect 25957 3090 26023 3093
rect 24209 3088 26023 3090
rect 24209 3032 24214 3088
rect 24270 3032 25962 3088
rect 26018 3032 26023 3088
rect 24209 3030 26023 3032
rect 24209 3027 24275 3030
rect 25957 3027 26023 3030
rect 6913 2954 6979 2957
rect 12525 2954 12591 2957
rect 6913 2952 12591 2954
rect 6913 2896 6918 2952
rect 6974 2896 12530 2952
rect 12586 2896 12591 2952
rect 6913 2894 12591 2896
rect 6913 2891 6979 2894
rect 12525 2891 12591 2894
rect 13537 2954 13603 2957
rect 18689 2954 18755 2957
rect 13537 2952 18755 2954
rect 13537 2896 13542 2952
rect 13598 2896 18694 2952
rect 18750 2896 18755 2952
rect 13537 2894 18755 2896
rect 13537 2891 13603 2894
rect 18689 2891 18755 2894
rect 18873 2954 18939 2957
rect 26509 2954 26575 2957
rect 18873 2952 26575 2954
rect 18873 2896 18878 2952
rect 18934 2896 26514 2952
rect 26570 2896 26575 2952
rect 18873 2894 26575 2896
rect 18873 2891 18939 2894
rect 26509 2891 26575 2894
rect 1853 2818 1919 2821
rect 2681 2818 2747 2821
rect 1853 2816 2747 2818
rect 1853 2760 1858 2816
rect 1914 2760 2686 2816
rect 2742 2760 2747 2816
rect 1853 2758 2747 2760
rect 1853 2755 1919 2758
rect 2681 2755 2747 2758
rect 2865 2818 2931 2821
rect 9213 2818 9279 2821
rect 2865 2816 9279 2818
rect 2865 2760 2870 2816
rect 2926 2760 9218 2816
rect 9274 2760 9279 2816
rect 2865 2758 9279 2760
rect 2865 2755 2931 2758
rect 9213 2755 9279 2758
rect 24761 2818 24827 2821
rect 27613 2818 27679 2821
rect 24761 2816 27679 2818
rect 24761 2760 24766 2816
rect 24822 2760 27618 2816
rect 27674 2760 27679 2816
rect 24761 2758 27679 2760
rect 24761 2755 24827 2758
rect 27613 2755 27679 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 4613 2682 4679 2685
rect 7465 2682 7531 2685
rect 4613 2680 7531 2682
rect 4613 2624 4618 2680
rect 4674 2624 7470 2680
rect 7526 2624 7531 2680
rect 4613 2622 7531 2624
rect 4613 2619 4679 2622
rect 7465 2619 7531 2622
rect 11329 2682 11395 2685
rect 14089 2682 14155 2685
rect 11329 2680 14155 2682
rect 11329 2624 11334 2680
rect 11390 2624 14094 2680
rect 14150 2624 14155 2680
rect 11329 2622 14155 2624
rect 11329 2619 11395 2622
rect 14089 2619 14155 2622
rect 0 2546 480 2576
rect 1577 2546 1643 2549
rect 0 2544 1643 2546
rect 0 2488 1582 2544
rect 1638 2488 1643 2544
rect 0 2486 1643 2488
rect 0 2456 480 2486
rect 1577 2483 1643 2486
rect 9673 2546 9739 2549
rect 12617 2546 12683 2549
rect 9673 2544 12683 2546
rect 9673 2488 9678 2544
rect 9734 2488 12622 2544
rect 12678 2488 12683 2544
rect 9673 2486 12683 2488
rect 9673 2483 9739 2486
rect 12617 2483 12683 2486
rect 14181 2546 14247 2549
rect 18505 2546 18571 2549
rect 14181 2544 18571 2546
rect 14181 2488 14186 2544
rect 14242 2488 18510 2544
rect 18566 2488 18571 2544
rect 14181 2486 18571 2488
rect 14181 2483 14247 2486
rect 18505 2483 18571 2486
rect 20621 2546 20687 2549
rect 22461 2546 22527 2549
rect 20621 2544 22527 2546
rect 20621 2488 20626 2544
rect 20682 2488 22466 2544
rect 22522 2488 22527 2544
rect 20621 2486 22527 2488
rect 20621 2483 20687 2486
rect 22461 2483 22527 2486
rect 8661 2410 8727 2413
rect 15193 2410 15259 2413
rect 8661 2408 15259 2410
rect 8661 2352 8666 2408
rect 8722 2352 15198 2408
rect 15254 2352 15259 2408
rect 8661 2350 15259 2352
rect 8661 2347 8727 2350
rect 15193 2347 15259 2350
rect 15469 2410 15535 2413
rect 21173 2410 21239 2413
rect 15469 2408 21239 2410
rect 15469 2352 15474 2408
rect 15530 2352 21178 2408
rect 21234 2352 21239 2408
rect 15469 2350 21239 2352
rect 15469 2347 15535 2350
rect 21173 2347 21239 2350
rect 7373 2274 7439 2277
rect 12065 2274 12131 2277
rect 7373 2272 12131 2274
rect 7373 2216 7378 2272
rect 7434 2216 12070 2272
rect 12126 2216 12131 2272
rect 7373 2214 12131 2216
rect 7373 2211 7439 2214
rect 12065 2211 12131 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 7557 2138 7623 2141
rect 12433 2138 12499 2141
rect 7557 2136 12499 2138
rect 7557 2080 7562 2136
rect 7618 2080 12438 2136
rect 12494 2080 12499 2136
rect 7557 2078 12499 2080
rect 7557 2075 7623 2078
rect 12433 2075 12499 2078
rect 0 2002 480 2032
rect 2129 2002 2195 2005
rect 0 2000 2195 2002
rect 0 1944 2134 2000
rect 2190 1944 2195 2000
rect 0 1942 2195 1944
rect 0 1912 480 1942
rect 2129 1939 2195 1942
rect 13077 2002 13143 2005
rect 18873 2002 18939 2005
rect 13077 2000 18939 2002
rect 13077 1944 13082 2000
rect 13138 1944 18878 2000
rect 18934 1944 18939 2000
rect 13077 1942 18939 1944
rect 13077 1939 13143 1942
rect 18873 1939 18939 1942
rect 657 1866 723 1869
rect 6637 1866 6703 1869
rect 657 1864 6703 1866
rect 657 1808 662 1864
rect 718 1808 6642 1864
rect 6698 1808 6703 1864
rect 657 1806 6703 1808
rect 657 1803 723 1806
rect 6637 1803 6703 1806
rect 7925 1866 7991 1869
rect 18321 1866 18387 1869
rect 7925 1864 18387 1866
rect 7925 1808 7930 1864
rect 7986 1808 18326 1864
rect 18382 1808 18387 1864
rect 7925 1806 18387 1808
rect 7925 1803 7991 1806
rect 18321 1803 18387 1806
rect 1761 1730 1827 1733
rect 9397 1730 9463 1733
rect 1761 1728 9463 1730
rect 1761 1672 1766 1728
rect 1822 1672 9402 1728
rect 9458 1672 9463 1728
rect 1761 1670 9463 1672
rect 1761 1667 1827 1670
rect 9397 1667 9463 1670
rect 0 1458 480 1488
rect 1301 1458 1367 1461
rect 0 1456 1367 1458
rect 0 1400 1306 1456
rect 1362 1400 1367 1456
rect 0 1398 1367 1400
rect 0 1368 480 1398
rect 1301 1395 1367 1398
rect 11605 1458 11671 1461
rect 16573 1458 16639 1461
rect 11605 1456 16639 1458
rect 11605 1400 11610 1456
rect 11666 1400 16578 1456
rect 16634 1400 16639 1456
rect 11605 1398 16639 1400
rect 11605 1395 11671 1398
rect 16573 1395 16639 1398
rect 19333 1458 19399 1461
rect 22645 1458 22711 1461
rect 19333 1456 22711 1458
rect 19333 1400 19338 1456
rect 19394 1400 22650 1456
rect 22706 1400 22711 1456
rect 19333 1398 22711 1400
rect 19333 1395 19399 1398
rect 22645 1395 22711 1398
rect 10593 1050 10659 1053
rect 10726 1050 10732 1052
rect 10593 1048 10732 1050
rect 10593 992 10598 1048
rect 10654 992 10732 1048
rect 10593 990 10732 992
rect 10593 987 10659 990
rect 10726 988 10732 990
rect 10796 988 10802 1052
rect 0 914 480 944
rect 1025 914 1091 917
rect 0 912 1091 914
rect 0 856 1030 912
rect 1086 856 1091 912
rect 0 854 1091 856
rect 0 824 480 854
rect 1025 851 1091 854
rect 0 370 480 400
rect 1117 370 1183 373
rect 0 368 1183 370
rect 0 312 1122 368
rect 1178 312 1183 368
rect 0 310 1183 312
rect 0 280 480 310
rect 1117 307 1183 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 10732 7788 10796 7852
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 8156 4932 8220 4996
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 8156 4660 8220 4724
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 10732 988 10796 1052
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 10731 7852 10797 7853
rect 10731 7788 10732 7852
rect 10796 7788 10797 7852
rect 10731 7787 10797 7788
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 8155 4996 8221 4997
rect 8155 4932 8156 4996
rect 8220 4932 8221 4996
rect 8155 4931 8221 4932
rect 8158 4725 8218 4931
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 8155 4724 8221 4725
rect 8155 4660 8156 4724
rect 8220 4660 8221 4724
rect 8155 4659 8221 4660
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 10734 1053 10794 7787
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 10731 1052 10797 1053
rect 10731 988 10732 1052
rect 10796 988 10797 1052
rect 10731 987 10797 988
use sky130_fd_sc_hd__decap_3  FILLER_1_6 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _068_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1604681595
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_71
timestamp 1604681595
transform 1 0 7636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1604681595
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8648 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1604681595
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp 1604681595
transform 1 0 10764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107
timestamp 1604681595
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_127
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1604681595
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1604681595
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_146
timestamp 1604681595
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_176
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_168
timestamp 1604681595
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1604681595
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1604681595
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1604681595
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1604681595
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_224
timestamp 1604681595
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1604681595
transform 1 0 22908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_233
timestamp 1604681595
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_236
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_241
timestamp 1604681595
transform 1 0 23276 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1604681595
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_259 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2300 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_8
timestamp 1604681595
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_12
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1604681595
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1604681595
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1604681595
transform 1 0 3496 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1604681595
transform 1 0 4692 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5428 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_43
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1604681595
transform 1 0 5336 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7912 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1604681595
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1604681595
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_83
timestamp 1604681595
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_87
timestamp 1604681595
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12144 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1604681595
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1604681595
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_133
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_137
timestamp 1604681595
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1604681595
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1604681595
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_194
timestamp 1604681595
transform 1 0 18952 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1604681595
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_208
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 24012 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_231
timestamp 1604681595
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_243
timestamp 1604681595
transform 1 0 23460 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1604681595
transform 1 0 24380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_265
timestamp 1604681595
transform 1 0 25484 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_273
timestamp 1604681595
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1604681595
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_85
timestamp 1604681595
transform 1 0 8924 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1604681595
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_103
timestamp 1604681595
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_107
timestamp 1604681595
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_142
timestamp 1604681595
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_146
timestamp 1604681595
transform 1 0 14536 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_152
timestamp 1604681595
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 21160 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_210
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_214
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1604681595
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_226
timestamp 1604681595
transform 1 0 21896 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 22264 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_233
timestamp 1604681595
transform 1 0 22540 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_241
timestamp 1604681595
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_40
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5244 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_64
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11592 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_108
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp 1604681595
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_138
timestamp 1604681595
transform 1 0 13800 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_160
timestamp 1604681595
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1604681595
transform 1 0 16192 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 19228 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_189
timestamp 1604681595
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1604681595
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1604681595
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_205
timestamp 1604681595
transform 1 0 19964 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604681595
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_231
timestamp 1604681595
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_243
timestamp 1604681595
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_255
timestamp 1604681595
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp 1604681595
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_31
timestamp 1604681595
transform 1 0 3956 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1604681595
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1604681595
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1604681595
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_83
timestamp 1604681595
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9476 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1604681595
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1604681595
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_173
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_203
timestamp 1604681595
transform 1 0 19780 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_219
timestamp 1604681595
transform 1 0 21252 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_231
timestamp 1604681595
transform 1 0 22356 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1604681595
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1604681595
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_16
timestamp 1604681595
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_20
timestamp 1604681595
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_26
timestamp 1604681595
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1604681595
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1604681595
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1604681595
transform 1 0 3312 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_47
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1604681595
transform 1 0 5336 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_42
timestamp 1604681595
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5428 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_70
timestamp 1604681595
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1604681595
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_83
timestamp 1604681595
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7912 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 1604681595
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_96
timestamp 1604681595
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_100
timestamp 1604681595
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_104
timestamp 1604681595
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_108
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10856 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_136
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14076 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_160
timestamp 1604681595
transform 1 0 15824 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_164
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_174
timestamp 1604681595
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1604681595
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1604681595
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_186
timestamp 1604681595
transform 1 0 18216 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_183
timestamp 1604681595
transform 1 0 17940 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_179
timestamp 1604681595
transform 1 0 17572 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_187
timestamp 1604681595
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1604681595
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_195
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_202
timestamp 1604681595
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_206
timestamp 1604681595
transform 1 0 20056 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_214
timestamp 1604681595
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_217
timestamp 1604681595
transform 1 0 21068 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_241
timestamp 1604681595
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4968 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_51
timestamp 1604681595
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 1604681595
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604681595
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1604681595
transform 1 0 8924 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1604681595
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_111
timestamp 1604681595
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1604681595
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1604681595
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_142
timestamp 1604681595
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 14536 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_161
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_165
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16836 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp 1604681595
transform 1 0 16560 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_219
timestamp 1604681595
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_231
timestamp 1604681595
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_243
timestamp 1604681595
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_255
timestamp 1604681595
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_267
timestamp 1604681595
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2760 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1604681595
transform 1 0 1656 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_16
timestamp 1604681595
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1604681595
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_41
timestamp 1604681595
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 5244 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1604681595
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_52
timestamp 1604681595
transform 1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1604681595
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_152
timestamp 1604681595
transform 1 0 15088 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1604681595
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19688 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_212
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_224
timestamp 1604681595
transform 1 0 21712 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1604681595
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1604681595
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1604681595
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_38
timestamp 1604681595
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_46
timestamp 1604681595
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_57
timestamp 1604681595
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1604681595
transform 1 0 6716 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_64
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_81
timestamp 1604681595
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1604681595
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1604681595
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1604681595
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 1604681595
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11040 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1604681595
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1604681595
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_165
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16744 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_168
timestamp 1604681595
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_189
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1604681595
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2208 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_8
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1604681595
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_37
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_90
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_94
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_111
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_107
timestamp 1604681595
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14168 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_138
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1604681595
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_165
timestamp 1604681595
transform 1 0 16284 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_172
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1604681595
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_214
timestamp 1604681595
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_218
timestamp 1604681595
transform 1 0 21160 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_230
timestamp 1604681595
transform 1 0 22264 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_11
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_36
timestamp 1604681595
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_63
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11408 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1604681595
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1604681595
transform 1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_131
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_135
timestamp 1604681595
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1604681595
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_173
timestamp 1604681595
transform 1 0 17020 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_185
timestamp 1604681595
transform 1 0 18124 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1604681595
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1604681595
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1472 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_13
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_17
timestamp 1604681595
transform 1 0 2668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3128 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_41
timestamp 1604681595
transform 1 0 4876 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_26
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1604681595
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1604681595
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_55
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_112
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11408 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604681595
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_161
timestamp 1604681595
transform 1 0 15916 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_146
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_173
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604681595
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_8
timestamp 1604681595
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_25
timestamp 1604681595
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_29
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_46
timestamp 1604681595
transform 1 0 5336 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_49
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 6900 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_144
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_168
timestamp 1604681595
transform 1 0 16560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 1472 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4140 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_39
timestamp 1604681595
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5428 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_83
timestamp 1604681595
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1604681595
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1604681595
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1604681595
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1604681595
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_138
timestamp 1604681595
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1604681595
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_24
timestamp 1604681595
transform 1 0 3312 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8096 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_68
timestamp 1604681595
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_72
timestamp 1604681595
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_168
timestamp 1604681595
transform 1 0 16560 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_224
timestamp 1604681595
transform 1 0 21712 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_227
timestamp 1604681595
transform 1 0 21988 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1604681595
transform 1 0 23092 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1604681595
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_12
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_17
timestamp 1604681595
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4324 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_71
timestamp 1604681595
transform 1 0 7636 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_76
timestamp 1604681595
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9936 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1604681595
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_119
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_142
timestamp 1604681595
transform 1 0 14168 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1604681595
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 21804 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_223
timestamp 1604681595
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_229
timestamp 1604681595
transform 1 0 22172 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_241
timestamp 1604681595
transform 1 0 23276 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1604681595
transform 1 0 24380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1604681595
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1604681595
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1604681595
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_38
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_46
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1604681595
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_49
timestamp 1604681595
transform 1 0 5612 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_44
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 5888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1604681595
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_55
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5428 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1604681595
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1604681595
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_67
timestamp 1604681595
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_83
timestamp 1604681595
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_87
timestamp 1604681595
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_106
timestamp 1604681595
transform 1 0 10856 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_135
timestamp 1604681595
transform 1 0 13524 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_147
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_228
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 22356 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_233
timestamp 1604681595
transform 1 0 22540 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_241
timestamp 1604681595
transform 1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_235
timestamp 1604681595
transform 1 0 22724 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2116 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1604681595
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8096 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_65
timestamp 1604681595
transform 1 0 7084 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1604681595
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1604681595
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1604681595
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_163
timestamp 1604681595
transform 1 0 16100 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_249
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1604681595
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1604681595
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5244 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_71
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_81
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1604681595
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1604681595
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_100
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_127
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_142
timestamp 1604681595
transform 1 0 14168 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1604681595
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 23368 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_246
timestamp 1604681595
transform 1 0 23736 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1604681595
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604681595
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3864 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_23
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1604681595
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5428 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1604681595
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 7084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8096 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1604681595
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_72
timestamp 1604681595
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_95
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_112
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1604681595
transform 1 0 14812 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_161
timestamp 1604681595
transform 1 0 15916 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_173
timestamp 1604681595
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_14
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4692 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1604681595
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_26
timestamp 1604681595
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_36
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_62
timestamp 1604681595
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 7176 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1604681595
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 9936 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_99
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_104
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1604681595
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1604681595
transform 1 0 13064 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1604681595
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_65
timestamp 1604681595
transform 1 0 7084 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_94
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_111
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1604681595
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1604681595
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1604681595
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_163
timestamp 1604681595
transform 1 0 16100 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_6
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1564 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_10
timestamp 1604681595
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_41
timestamp 1604681595
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1604681595
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_45
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 1604681595
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1604681595
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 5612 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6164 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6992 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7912 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_83
timestamp 1604681595
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_87
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_87
timestamp 1604681595
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_106
timestamp 1604681595
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_142
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_166
timestamp 1604681595
transform 1 0 16376 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1604681595
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1604681595
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_21
timestamp 1604681595
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_25
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5796 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_70
timestamp 1604681595
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_81
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 9936 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1604681595
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_99
timestamp 1604681595
transform 1 0 10212 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_103
timestamp 1604681595
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_126
timestamp 1604681595
transform 1 0 12696 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_138
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1604681595
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 1604681595
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3772 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_21
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_25
timestamp 1604681595
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_48
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_52
timestamp 1604681595
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_56
timestamp 1604681595
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7544 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_66
timestamp 1604681595
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_83
timestamp 1604681595
transform 1 0 8740 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 2760 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_14
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1604681595
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1604681595
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1604681595
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4692 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_62
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_75
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1604681595
transform 1 0 10028 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_101
timestamp 1604681595
transform 1 0 10396 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_123
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_127
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_17
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_20
timestamp 1604681595
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3312 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4876 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp 1604681595
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1604681595
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 6992 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8280 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp 1604681595
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_75
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1604681595
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_136
timestamp 1604681595
transform 1 0 13616 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_148
timestamp 1604681595
transform 1 0 14720 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_160
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 2760 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1604681595
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_14
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_22
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_26
timestamp 1604681595
transform 1 0 3496 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604681595
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_38
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 5336 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_42
timestamp 1604681595
transform 1 0 4968 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_50
timestamp 1604681595
transform 1 0 5704 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_55
timestamp 1604681595
transform 1 0 6164 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1604681595
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_96
timestamp 1604681595
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_100
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_32_124
timestamp 1604681595
transform 1 0 12512 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_136
timestamp 1604681595
transform 1 0 13616 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1604681595
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1604681595
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_11
timestamp 1604681595
transform 1 0 2116 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_14
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_10
timestamp 1604681595
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2760 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 2852 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_28
timestamp 1604681595
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_24
timestamp 1604681595
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_40
timestamp 1604681595
transform 1 0 4784 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_36
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_36
timestamp 1604681595
transform 1 0 4416 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_48
timestamp 1604681595
transform 1 0 5520 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_48
timestamp 1604681595
transform 1 0 5520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_52
timestamp 1604681595
transform 1 0 5888 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_52
timestamp 1604681595
transform 1 0 5888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5980 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 5612 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_59
timestamp 1604681595
transform 1 0 6532 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_73
timestamp 1604681595
transform 1 0 7820 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_83
timestamp 1604681595
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_63
timestamp 1604681595
transform 1 0 6900 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1604681595
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_78
timestamp 1604681595
transform 1 0 8280 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_37.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_102
timestamp 1604681595
transform 1 0 10488 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_108
timestamp 1604681595
transform 1 0 11040 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_120
timestamp 1604681595
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_39.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 12880 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_142
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_131
timestamp 1604681595
transform 1 0 13156 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_143
timestamp 1604681595
transform 1 0 14260 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_154
timestamp 1604681595
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_166
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_151
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1604681595
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1604681595
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2944 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_12
timestamp 1604681595
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_16
timestamp 1604681595
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_26
timestamp 1604681595
transform 1 0 3496 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_30
timestamp 1604681595
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_38
timestamp 1604681595
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_54
timestamp 1604681595
transform 1 0 6072 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1604681595
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_76
timestamp 1604681595
transform 1 0 8096 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_88
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_100
timestamp 1604681595
transform 1 0 10304 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_112
timestamp 1604681595
transform 1 0 11408 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1604681595
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_12
timestamp 1604681595
transform 1 0 2208 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_24
timestamp 1604681595
transform 1 0 3312 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_30
timestamp 1604681595
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_36
timestamp 1604681595
transform 1 0 4416 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_48
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_60
timestamp 1604681595
transform 1 0 6624 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7912 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1604681595
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 2852 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2668 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_11
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_23
timestamp 1604681595
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_31
timestamp 1604681595
transform 1 0 3956 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_34
timestamp 1604681595
transform 1 0 4232 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_46
timestamp 1604681595
transform 1 0 5336 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_58
timestamp 1604681595
transform 1 0 6440 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604681595
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604681595
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_12
timestamp 1604681595
transform 1 0 2208 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_24
timestamp 1604681595
transform 1 0 3312 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_30
timestamp 1604681595
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_36
timestamp 1604681595
transform 1 0 4416 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_48
timestamp 1604681595
transform 1 0 5520 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_60
timestamp 1604681595
transform 1 0 6624 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_72
timestamp 1604681595
transform 1 0 7728 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_84
timestamp 1604681595
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1604681595
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604681595
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_16
timestamp 1604681595
transform 1 0 2576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_12
timestamp 1604681595
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 2944 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_24
timestamp 1604681595
transform 1 0 3312 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_28
timestamp 1604681595
transform 1 0 3680 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_40
timestamp 1604681595
transform 1 0 4784 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_52
timestamp 1604681595
transform 1 0 5888 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_60
timestamp 1604681595
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_66
timestamp 1604681595
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1604681595
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1604681595
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1604681595
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_106
timestamp 1604681595
transform 1 0 10856 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 19780 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_196
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_202
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_207
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_219
timestamp 1604681595
transform 1 0 21252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_231
timestamp 1604681595
transform 1 0 22356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1604681595
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1604681595
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 27066 0 27122 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 7010 27520 7066 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 27618 0 27674 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 20994 27520 21050 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 4 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 5 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_44_
port 6 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_45_
port 7 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_46_
port 8 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_47_
port 9 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_48_
port 10 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_left_grid_pin_49_
port 11 nsew default input
rlabel metal2 s 26514 0 26570 480 6 bottom_right_grid_pin_1_
port 12 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_head
port 13 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 ccff_tail
port 14 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[10]
port 16 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[11]
port 17 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[12]
port 18 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[13]
port 19 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[14]
port 20 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[15]
port 21 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[16]
port 22 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[17]
port 23 nsew default input
rlabel metal3 s 0 15104 480 15224 6 chanx_left_in[18]
port 24 nsew default input
rlabel metal3 s 0 15648 480 15768 6 chanx_left_in[19]
port 25 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[1]
port 26 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[2]
port 27 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[3]
port 28 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[4]
port 29 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[5]
port 30 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[6]
port 31 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[7]
port 32 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[8]
port 33 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[9]
port 34 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[0]
port 35 nsew default tristate
rlabel metal3 s 0 21904 480 22024 6 chanx_left_out[10]
port 36 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[11]
port 37 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[12]
port 38 nsew default tristate
rlabel metal3 s 0 23672 480 23792 6 chanx_left_out[13]
port 39 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[14]
port 40 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[15]
port 41 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[16]
port 42 nsew default tristate
rlabel metal3 s 0 25984 480 26104 6 chanx_left_out[17]
port 43 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[18]
port 44 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[19]
port 45 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[1]
port 46 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[2]
port 47 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[3]
port 48 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 49 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 50 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[6]
port 51 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 52 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[8]
port 53 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[9]
port 54 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[0]
port 55 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[10]
port 56 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[11]
port 57 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[12]
port 58 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[13]
port 59 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[14]
port 60 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[15]
port 61 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[16]
port 62 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[17]
port 63 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_in[18]
port 64 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[19]
port 65 nsew default input
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[1]
port 66 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chany_bottom_in[2]
port 67 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[3]
port 68 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[4]
port 69 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[5]
port 70 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[6]
port 71 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[7]
port 72 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[8]
port 73 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[9]
port 74 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[0]
port 75 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[10]
port 76 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[11]
port 77 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[12]
port 78 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[13]
port 79 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[14]
port 80 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[15]
port 81 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[16]
port 82 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[17]
port 83 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[18]
port 84 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[19]
port 85 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_out[1]
port 86 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[2]
port 87 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[3]
port 88 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[4]
port 89 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[5]
port 90 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[6]
port 91 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 92 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[8]
port 93 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[9]
port 94 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 95 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 96 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 97 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 98 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_38_
port 99 nsew default input
rlabel metal3 s 0 3136 480 3256 6 left_bottom_grid_pin_39_
port 100 nsew default input
rlabel metal3 s 0 3680 480 3800 6 left_bottom_grid_pin_40_
port 101 nsew default input
rlabel metal3 s 0 4224 480 4344 6 left_bottom_grid_pin_41_
port 102 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_1_
port 103 nsew default input
rlabel metal3 s 27520 4632 28000 4752 6 prog_clk
port 104 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 105 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 106 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
