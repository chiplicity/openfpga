magic
tech sky130A
magscale 1 2
timestamp 1605003321
<< locali >>
rect 22557 12699 22591 12937
rect 22097 2839 22131 3145
<< viali >>
rect 23845 24361 23879 24395
rect 24489 23817 24523 23851
rect 24305 23613 24339 23647
rect 24857 23613 24891 23647
rect 10689 23273 10723 23307
rect 24489 23273 24523 23307
rect 10505 23137 10539 23171
rect 24305 23137 24339 23171
rect 24857 22729 24891 22763
rect 23661 22593 23695 22627
rect 23385 22525 23419 22559
rect 24673 22525 24707 22559
rect 25225 22525 25259 22559
rect 23201 22457 23235 22491
rect 10505 22389 10539 22423
rect 24397 22389 24431 22423
rect 9769 22117 9803 22151
rect 9493 22049 9527 22083
rect 12161 22049 12195 22083
rect 24305 22049 24339 22083
rect 12437 21981 12471 22015
rect 24489 21913 24523 21947
rect 24489 21641 24523 21675
rect 14737 21437 14771 21471
rect 15473 21437 15507 21471
rect 24121 21437 24155 21471
rect 24305 21437 24339 21471
rect 24857 21437 24891 21471
rect 15013 21369 15047 21403
rect 9493 21301 9527 21335
rect 12345 21301 12379 21335
rect 24765 21097 24799 21131
rect 23569 21029 23603 21063
rect 23293 20961 23327 20995
rect 24581 20961 24615 20995
rect 23569 20553 23603 20587
rect 23201 20349 23235 20383
rect 23385 20349 23419 20383
rect 23937 20349 23971 20383
rect 24581 20213 24615 20247
rect 24489 20009 24523 20043
rect 21453 19941 21487 19975
rect 22741 19941 22775 19975
rect 21177 19873 21211 19907
rect 22465 19873 22499 19907
rect 24305 19873 24339 19907
rect 24305 19261 24339 19295
rect 24857 19261 24891 19295
rect 21177 19125 21211 19159
rect 22465 19125 22499 19159
rect 24121 19125 24155 19159
rect 24489 19125 24523 19159
rect 11149 18921 11183 18955
rect 10965 18785 10999 18819
rect 15473 18785 15507 18819
rect 15749 18785 15783 18819
rect 24857 18377 24891 18411
rect 23661 18241 23695 18275
rect 23385 18173 23419 18207
rect 24121 18173 24155 18207
rect 24673 18173 24707 18207
rect 25225 18173 25259 18207
rect 10965 18037 10999 18071
rect 15473 18037 15507 18071
rect 10321 17765 10355 17799
rect 10045 17697 10079 17731
rect 15841 17697 15875 17731
rect 16025 17561 16059 17595
rect 24489 17289 24523 17323
rect 12621 17085 12655 17119
rect 13357 17085 13391 17119
rect 24305 17085 24339 17119
rect 24857 17085 24891 17119
rect 12897 17017 12931 17051
rect 10045 16949 10079 16983
rect 15841 16949 15875 16983
rect 24489 16745 24523 16779
rect 15289 16677 15323 16711
rect 15013 16609 15047 16643
rect 24305 16609 24339 16643
rect 24489 16201 24523 16235
rect 18233 16065 18267 16099
rect 17957 15997 17991 16031
rect 24305 15997 24339 16031
rect 24857 15997 24891 16031
rect 15013 15861 15047 15895
rect 18785 15861 18819 15895
rect 24121 15861 24155 15895
rect 23385 15589 23419 15623
rect 23109 15521 23143 15555
rect 24397 15521 24431 15555
rect 24581 15317 24615 15351
rect 24397 15113 24431 15147
rect 25041 15113 25075 15147
rect 23845 14977 23879 15011
rect 23201 14909 23235 14943
rect 23569 14909 23603 14943
rect 24857 14909 24891 14943
rect 25409 14909 25443 14943
rect 22741 14773 22775 14807
rect 24581 14569 24615 14603
rect 23385 14501 23419 14535
rect 23109 14433 23143 14467
rect 24397 14433 24431 14467
rect 20625 14365 20659 14399
rect 24489 14025 24523 14059
rect 24857 13957 24891 13991
rect 18601 13889 18635 13923
rect 18325 13821 18359 13855
rect 19061 13821 19095 13855
rect 23109 13821 23143 13855
rect 24305 13821 24339 13855
rect 20165 13685 20199 13719
rect 21913 13685 21947 13719
rect 24121 13685 24155 13719
rect 20625 13481 20659 13515
rect 20993 13481 21027 13515
rect 22925 13481 22959 13515
rect 24489 13481 24523 13515
rect 22833 13345 22867 13379
rect 24305 13345 24339 13379
rect 19245 13277 19279 13311
rect 21085 13277 21119 13311
rect 21269 13277 21303 13311
rect 23109 13277 23143 13311
rect 19061 13141 19095 13175
rect 20441 13141 20475 13175
rect 22465 13141 22499 13175
rect 23477 13141 23511 13175
rect 18969 12937 19003 12971
rect 21545 12937 21579 12971
rect 22557 12937 22591 12971
rect 22833 12937 22867 12971
rect 23201 12937 23235 12971
rect 24857 12937 24891 12971
rect 25317 12937 25351 12971
rect 19429 12801 19463 12835
rect 19521 12801 19555 12835
rect 21177 12801 21211 12835
rect 21913 12801 21947 12835
rect 18509 12733 18543 12767
rect 20073 12733 20107 12767
rect 20993 12733 21027 12767
rect 24305 12869 24339 12903
rect 23661 12801 23695 12835
rect 23385 12733 23419 12767
rect 24673 12733 24707 12767
rect 18785 12665 18819 12699
rect 19337 12665 19371 12699
rect 20441 12665 20475 12699
rect 20901 12665 20935 12699
rect 22557 12665 22591 12699
rect 17957 12597 17991 12631
rect 20533 12597 20567 12631
rect 22281 12597 22315 12631
rect 20441 12393 20475 12427
rect 22649 12393 22683 12427
rect 24489 12393 24523 12427
rect 16669 12325 16703 12359
rect 17926 12325 17960 12359
rect 16393 12257 16427 12291
rect 17589 12257 17623 12291
rect 17681 12257 17715 12291
rect 20892 12257 20926 12291
rect 23376 12257 23410 12291
rect 20625 12189 20659 12223
rect 23109 12189 23143 12223
rect 22005 12121 22039 12155
rect 19061 12053 19095 12087
rect 19705 12053 19739 12087
rect 22925 12053 22959 12087
rect 20993 11849 21027 11883
rect 21545 11849 21579 11883
rect 22833 11849 22867 11883
rect 24489 11849 24523 11883
rect 24765 11849 24799 11883
rect 25133 11849 25167 11883
rect 16485 11781 16519 11815
rect 17773 11781 17807 11815
rect 15933 11713 15967 11747
rect 18325 11713 18359 11747
rect 18785 11713 18819 11747
rect 19613 11713 19647 11747
rect 23845 11713 23879 11747
rect 23937 11713 23971 11747
rect 15105 11645 15139 11679
rect 22189 11645 22223 11679
rect 24949 11645 24983 11679
rect 25501 11645 25535 11679
rect 15381 11577 15415 11611
rect 16669 11577 16703 11611
rect 17497 11577 17531 11611
rect 18141 11577 18175 11611
rect 19858 11577 19892 11611
rect 23753 11577 23787 11611
rect 17221 11509 17255 11543
rect 18233 11509 18267 11543
rect 19521 11509 19555 11543
rect 22005 11509 22039 11543
rect 22373 11509 22407 11543
rect 23201 11509 23235 11543
rect 23385 11509 23419 11543
rect 17865 11305 17899 11339
rect 18969 11305 19003 11339
rect 19337 11305 19371 11339
rect 20993 11305 21027 11339
rect 18877 11237 18911 11271
rect 21085 11237 21119 11271
rect 22548 11237 22582 11271
rect 13633 11169 13667 11203
rect 15013 11169 15047 11203
rect 15289 11169 15323 11203
rect 15841 11169 15875 11203
rect 16485 11169 16519 11203
rect 16741 11169 16775 11203
rect 19429 11169 19463 11203
rect 20073 11169 20107 11203
rect 20441 11169 20475 11203
rect 24765 11169 24799 11203
rect 13817 11101 13851 11135
rect 19521 11101 19555 11135
rect 21269 11101 21303 11135
rect 22281 11101 22315 11135
rect 18417 11033 18451 11067
rect 20625 11033 20659 11067
rect 24949 11033 24983 11067
rect 16209 10965 16243 10999
rect 21821 10965 21855 10999
rect 23661 10965 23695 10999
rect 24305 10965 24339 10999
rect 13357 10761 13391 10795
rect 16117 10761 16151 10795
rect 18693 10761 18727 10795
rect 20717 10761 20751 10795
rect 21177 10761 21211 10795
rect 21637 10761 21671 10795
rect 22741 10761 22775 10795
rect 25409 10761 25443 10795
rect 14185 10693 14219 10727
rect 15197 10693 15231 10727
rect 21729 10693 21763 10727
rect 13725 10625 13759 10659
rect 14737 10625 14771 10659
rect 16669 10625 16703 10659
rect 18785 10625 18819 10659
rect 22281 10625 22315 10659
rect 23109 10625 23143 10659
rect 16025 10557 16059 10591
rect 16485 10557 16519 10591
rect 17129 10557 17163 10591
rect 17589 10557 17623 10591
rect 19041 10557 19075 10591
rect 22189 10557 22223 10591
rect 23385 10557 23419 10591
rect 23641 10557 23675 10591
rect 14093 10489 14127 10523
rect 14553 10489 14587 10523
rect 15657 10489 15691 10523
rect 18325 10489 18359 10523
rect 22097 10489 22131 10523
rect 14645 10421 14679 10455
rect 16577 10421 16611 10455
rect 17773 10421 17807 10455
rect 20165 10421 20199 10455
rect 24765 10421 24799 10455
rect 13909 10217 13943 10251
rect 17405 10217 17439 10251
rect 18877 10217 18911 10251
rect 19889 10217 19923 10251
rect 20441 10217 20475 10251
rect 20809 10217 20843 10251
rect 21913 10217 21947 10251
rect 23201 10217 23235 10251
rect 15350 10149 15384 10183
rect 19337 10149 19371 10183
rect 23560 10149 23594 10183
rect 14829 10081 14863 10115
rect 15105 10081 15139 10115
rect 18785 10081 18819 10115
rect 19245 10081 19279 10115
rect 21177 10081 21211 10115
rect 17865 10013 17899 10047
rect 19429 10013 19463 10047
rect 21269 10013 21303 10047
rect 21453 10013 21487 10047
rect 23293 10013 23327 10047
rect 17773 9945 17807 9979
rect 13633 9877 13667 9911
rect 14369 9877 14403 9911
rect 16485 9877 16519 9911
rect 18325 9877 18359 9911
rect 22281 9877 22315 9911
rect 22741 9877 22775 9911
rect 24673 9877 24707 9911
rect 15013 9673 15047 9707
rect 15565 9673 15599 9707
rect 24765 9673 24799 9707
rect 16117 9605 16151 9639
rect 17773 9605 17807 9639
rect 21085 9605 21119 9639
rect 22833 9605 22867 9639
rect 24489 9605 24523 9639
rect 13633 9537 13667 9571
rect 16669 9537 16703 9571
rect 18417 9537 18451 9571
rect 23201 9537 23235 9571
rect 23845 9537 23879 9571
rect 24029 9537 24063 9571
rect 19521 9469 19555 9503
rect 19705 9469 19739 9503
rect 19961 9469 19995 9503
rect 22189 9469 22223 9503
rect 24949 9469 24983 9503
rect 25685 9469 25719 9503
rect 13541 9401 13575 9435
rect 13878 9401 13912 9435
rect 17497 9401 17531 9435
rect 18141 9401 18175 9435
rect 22005 9401 22039 9435
rect 23753 9401 23787 9435
rect 25225 9401 25259 9435
rect 11057 9333 11091 9367
rect 12621 9333 12655 9367
rect 15933 9333 15967 9367
rect 16485 9333 16519 9367
rect 16577 9333 16611 9367
rect 17221 9333 17255 9367
rect 18233 9333 18267 9367
rect 18877 9333 18911 9367
rect 19337 9333 19371 9367
rect 21729 9333 21763 9367
rect 22373 9333 22407 9367
rect 23385 9333 23419 9367
rect 10597 9129 10631 9163
rect 13541 9129 13575 9163
rect 14093 9129 14127 9163
rect 15013 9129 15047 9163
rect 16577 9129 16611 9163
rect 17037 9129 17071 9163
rect 18693 9129 18727 9163
rect 19797 9129 19831 9163
rect 20441 9129 20475 9163
rect 20625 9129 20659 9163
rect 21821 9129 21855 9163
rect 12069 9061 12103 9095
rect 12406 9061 12440 9095
rect 14829 9061 14863 9095
rect 16209 9061 16243 9095
rect 17580 9061 17614 9095
rect 23376 9061 23410 9095
rect 10965 8993 10999 9027
rect 15381 8993 15415 9027
rect 15473 8993 15507 9027
rect 17221 8993 17255 9027
rect 20993 8993 21027 9027
rect 11057 8925 11091 8959
rect 11241 8925 11275 8959
rect 12161 8925 12195 8959
rect 15565 8925 15599 8959
rect 17313 8925 17347 8959
rect 21085 8925 21119 8959
rect 21177 8925 21211 8959
rect 23109 8925 23143 8959
rect 16945 8857 16979 8891
rect 10505 8789 10539 8823
rect 19337 8789 19371 8823
rect 22189 8789 22223 8823
rect 22649 8789 22683 8823
rect 23017 8789 23051 8823
rect 24489 8789 24523 8823
rect 25041 8789 25075 8823
rect 11425 8585 11459 8619
rect 11793 8585 11827 8619
rect 12621 8585 12655 8619
rect 13541 8585 13575 8619
rect 15105 8585 15139 8619
rect 16577 8585 16611 8619
rect 17405 8585 17439 8619
rect 18509 8585 18543 8619
rect 19981 8585 20015 8619
rect 20625 8585 20659 8619
rect 21637 8585 21671 8619
rect 24765 8585 24799 8619
rect 21729 8517 21763 8551
rect 23201 8517 23235 8551
rect 14093 8449 14127 8483
rect 15197 8449 15231 8483
rect 18601 8449 18635 8483
rect 22189 8449 22223 8483
rect 22373 8449 22407 8483
rect 9033 8381 9067 8415
rect 9493 8381 9527 8415
rect 13081 8381 13115 8415
rect 14001 8381 14035 8415
rect 18857 8381 18891 8415
rect 22097 8381 22131 8415
rect 23385 8381 23419 8415
rect 9401 8313 9435 8347
rect 9738 8313 9772 8347
rect 13357 8313 13391 8347
rect 13909 8313 13943 8347
rect 14737 8313 14771 8347
rect 15464 8313 15498 8347
rect 17957 8313 17991 8347
rect 20993 8313 21027 8347
rect 22833 8313 22867 8347
rect 23652 8313 23686 8347
rect 10873 8245 10907 8279
rect 12161 8245 12195 8279
rect 12069 8041 12103 8075
rect 13173 8041 13207 8075
rect 14829 8041 14863 8075
rect 16393 8041 16427 8075
rect 17865 8041 17899 8075
rect 20073 8041 20107 8075
rect 23201 8041 23235 8075
rect 23661 8041 23695 8075
rect 24673 8041 24707 8075
rect 10597 7905 10631 7939
rect 10956 7905 10990 7939
rect 13541 7905 13575 7939
rect 15269 7905 15303 7939
rect 17405 7905 17439 7939
rect 19245 7905 19279 7939
rect 20625 7905 20659 7939
rect 20892 7905 20926 7939
rect 23569 7905 23603 7939
rect 24765 7905 24799 7939
rect 9401 7837 9435 7871
rect 10689 7837 10723 7871
rect 13633 7837 13667 7871
rect 13725 7837 13759 7871
rect 14461 7837 14495 7871
rect 15013 7837 15047 7871
rect 17957 7837 17991 7871
rect 18049 7837 18083 7871
rect 19521 7837 19555 7871
rect 23753 7837 23787 7871
rect 12805 7769 12839 7803
rect 17497 7769 17531 7803
rect 18877 7769 18911 7803
rect 24949 7769 24983 7803
rect 7837 7701 7871 7735
rect 17037 7701 17071 7735
rect 18509 7701 18543 7735
rect 20441 7701 20475 7735
rect 22005 7701 22039 7735
rect 22557 7701 22591 7735
rect 22925 7701 22959 7735
rect 24213 7701 24247 7735
rect 7745 7497 7779 7531
rect 10505 7497 10539 7531
rect 12529 7497 12563 7531
rect 15105 7497 15139 7531
rect 20809 7497 20843 7531
rect 20901 7497 20935 7531
rect 21913 7497 21947 7531
rect 22465 7497 22499 7531
rect 22833 7497 22867 7531
rect 24765 7497 24799 7531
rect 25685 7497 25719 7531
rect 9217 7429 9251 7463
rect 16485 7429 16519 7463
rect 19337 7429 19371 7463
rect 23109 7429 23143 7463
rect 11149 7361 11183 7395
rect 11517 7361 11551 7395
rect 11977 7361 12011 7395
rect 12713 7361 12747 7395
rect 18325 7361 18359 7395
rect 19981 7361 20015 7395
rect 21453 7361 21487 7395
rect 24029 7361 24063 7395
rect 7837 7293 7871 7327
rect 12980 7293 13014 7327
rect 15197 7293 15231 7327
rect 19797 7293 19831 7327
rect 20441 7293 20475 7327
rect 25041 7293 25075 7327
rect 8082 7225 8116 7259
rect 10321 7225 10355 7259
rect 10873 7225 10907 7259
rect 18233 7225 18267 7259
rect 19245 7225 19279 7259
rect 19705 7225 19739 7259
rect 10045 7157 10079 7191
rect 10965 7157 10999 7191
rect 14093 7157 14127 7191
rect 14645 7157 14679 7191
rect 17497 7157 17531 7191
rect 17773 7157 17807 7191
rect 18141 7157 18175 7191
rect 18877 7157 18911 7191
rect 21269 7157 21303 7191
rect 21361 7157 21395 7191
rect 23477 7157 23511 7191
rect 23845 7157 23879 7191
rect 23937 7157 23971 7191
rect 25225 7157 25259 7191
rect 9769 6953 9803 6987
rect 11149 6953 11183 6987
rect 12805 6953 12839 6987
rect 13357 6953 13391 6987
rect 16025 6953 16059 6987
rect 18325 6953 18359 6987
rect 19245 6953 19279 6987
rect 19981 6953 20015 6987
rect 20625 6953 20659 6987
rect 24581 6953 24615 6987
rect 11057 6885 11091 6919
rect 15933 6885 15967 6919
rect 6825 6817 6859 6851
rect 7081 6817 7115 6851
rect 10505 6817 10539 6851
rect 11333 6817 11367 6851
rect 11425 6817 11459 6851
rect 11692 6817 11726 6851
rect 15197 6817 15231 6851
rect 16649 6817 16683 6851
rect 20993 6817 21027 6851
rect 22537 6817 22571 6851
rect 24765 6817 24799 6851
rect 9861 6749 9895 6783
rect 9953 6749 9987 6783
rect 13909 6749 13943 6783
rect 16117 6749 16151 6783
rect 16393 6749 16427 6783
rect 19337 6749 19371 6783
rect 19429 6749 19463 6783
rect 21085 6749 21119 6783
rect 21177 6749 21211 6783
rect 22281 6749 22315 6783
rect 9401 6681 9435 6715
rect 15381 6681 15415 6715
rect 15565 6681 15599 6715
rect 17773 6681 17807 6715
rect 18877 6681 18911 6715
rect 20441 6681 20475 6715
rect 24213 6681 24247 6715
rect 8205 6613 8239 6647
rect 13725 6613 13759 6647
rect 14369 6613 14403 6647
rect 14829 6613 14863 6647
rect 18693 6613 18727 6647
rect 21821 6613 21855 6647
rect 22189 6613 22223 6647
rect 23661 6613 23695 6647
rect 24949 6613 24983 6647
rect 6917 6409 6951 6443
rect 10045 6409 10079 6443
rect 12253 6409 12287 6443
rect 13357 6409 13391 6443
rect 15197 6409 15231 6443
rect 17221 6409 17255 6443
rect 18509 6409 18543 6443
rect 20349 6409 20383 6443
rect 20901 6409 20935 6443
rect 21545 6409 21579 6443
rect 21729 6409 21763 6443
rect 22741 6409 22775 6443
rect 25409 6409 25443 6443
rect 24857 6341 24891 6375
rect 12897 6273 12931 6307
rect 22373 6273 22407 6307
rect 7285 6205 7319 6239
rect 7653 6205 7687 6239
rect 8113 6205 8147 6239
rect 13817 6205 13851 6239
rect 15841 6205 15875 6239
rect 16577 6205 16611 6239
rect 17865 6205 17899 6239
rect 18969 6205 19003 6239
rect 23477 6205 23511 6239
rect 8021 6137 8055 6171
rect 8358 6137 8392 6171
rect 10413 6137 10447 6171
rect 10965 6137 10999 6171
rect 14062 6137 14096 6171
rect 17497 6137 17531 6171
rect 18877 6137 18911 6171
rect 19236 6137 19270 6171
rect 22097 6137 22131 6171
rect 23722 6137 23756 6171
rect 9493 6069 9527 6103
rect 11057 6069 11091 6103
rect 11517 6069 11551 6103
rect 11977 6069 12011 6103
rect 12621 6069 12655 6103
rect 12713 6069 12747 6103
rect 13633 6069 13667 6103
rect 16117 6069 16151 6103
rect 16761 6069 16795 6103
rect 18049 6069 18083 6103
rect 22189 6069 22223 6103
rect 23109 6069 23143 6103
rect 25869 6069 25903 6103
rect 26145 6069 26179 6103
rect 8757 5865 8791 5899
rect 9585 5865 9619 5899
rect 9861 5865 9895 5899
rect 10229 5865 10263 5899
rect 13909 5865 13943 5899
rect 14737 5865 14771 5899
rect 15565 5865 15599 5899
rect 17129 5865 17163 5899
rect 18969 5865 19003 5899
rect 19521 5865 19555 5899
rect 19889 5865 19923 5899
rect 22005 5865 22039 5899
rect 11333 5797 11367 5831
rect 17856 5797 17890 5831
rect 20870 5797 20904 5831
rect 23722 5797 23756 5831
rect 8113 5729 8147 5763
rect 11681 5729 11715 5763
rect 15013 5729 15047 5763
rect 16393 5729 16427 5763
rect 8205 5661 8239 5695
rect 8297 5661 8331 5695
rect 9217 5661 9251 5695
rect 10321 5661 10355 5695
rect 10413 5661 10447 5695
rect 11425 5661 11459 5695
rect 16485 5661 16519 5695
rect 16577 5661 16611 5695
rect 17589 5661 17623 5695
rect 20625 5661 20659 5695
rect 22557 5661 22591 5695
rect 23477 5661 23511 5695
rect 7745 5593 7779 5627
rect 13357 5593 13391 5627
rect 13725 5593 13759 5627
rect 14369 5593 14403 5627
rect 16025 5593 16059 5627
rect 17405 5593 17439 5627
rect 10965 5525 10999 5559
rect 12805 5525 12839 5559
rect 20441 5525 20475 5559
rect 22925 5525 22959 5559
rect 23293 5525 23327 5559
rect 24857 5525 24891 5559
rect 7469 5321 7503 5355
rect 8573 5321 8607 5355
rect 9677 5321 9711 5355
rect 10505 5321 10539 5355
rect 13541 5321 13575 5355
rect 14185 5321 14219 5355
rect 17221 5321 17255 5355
rect 17497 5321 17531 5355
rect 17773 5321 17807 5355
rect 19337 5321 19371 5355
rect 20625 5321 20659 5355
rect 22189 5321 22223 5355
rect 23569 5321 23603 5355
rect 25685 5321 25719 5355
rect 18785 5253 18819 5287
rect 24581 5253 24615 5287
rect 7561 5185 7595 5219
rect 9125 5185 9159 5219
rect 11057 5185 11091 5219
rect 11517 5185 11551 5219
rect 11977 5185 12011 5219
rect 15197 5185 15231 5219
rect 18233 5185 18267 5219
rect 18325 5185 18359 5219
rect 20809 5185 20843 5219
rect 23201 5185 23235 5219
rect 24029 5185 24063 5219
rect 24213 5185 24247 5219
rect 12161 5117 12195 5151
rect 12428 5117 12462 5151
rect 14553 5117 14587 5151
rect 14829 5117 14863 5151
rect 18141 5117 18175 5151
rect 19521 5117 19555 5151
rect 19705 5117 19739 5151
rect 20349 5117 20383 5151
rect 21065 5117 21099 5151
rect 25133 5117 25167 5151
rect 10045 5049 10079 5083
rect 10965 5049 10999 5083
rect 15442 5049 15476 5083
rect 23937 5049 23971 5083
rect 24949 5049 24983 5083
rect 8021 4981 8055 5015
rect 8389 4981 8423 5015
rect 8941 4981 8975 5015
rect 9033 4981 9067 5015
rect 10321 4981 10355 5015
rect 10873 4981 10907 5015
rect 14645 4981 14679 5015
rect 16577 4981 16611 5015
rect 19245 4981 19279 5015
rect 19889 4981 19923 5015
rect 22833 4981 22867 5015
rect 25317 4981 25351 5015
rect 26053 4981 26087 5015
rect 7837 4777 7871 4811
rect 8113 4777 8147 4811
rect 9861 4777 9895 4811
rect 11517 4777 11551 4811
rect 13357 4777 13391 4811
rect 14369 4777 14403 4811
rect 15289 4777 15323 4811
rect 15657 4777 15691 4811
rect 16117 4777 16151 4811
rect 17221 4777 17255 4811
rect 18325 4777 18359 4811
rect 19153 4777 19187 4811
rect 19889 4777 19923 4811
rect 22097 4777 22131 4811
rect 23201 4777 23235 4811
rect 23569 4777 23603 4811
rect 24305 4777 24339 4811
rect 17037 4709 17071 4743
rect 17681 4709 17715 4743
rect 10404 4641 10438 4675
rect 12897 4641 12931 4675
rect 13725 4641 13759 4675
rect 14829 4641 14863 4675
rect 16025 4641 16059 4675
rect 17589 4641 17623 4675
rect 22005 4641 22039 4675
rect 24765 4641 24799 4675
rect 8297 4573 8331 4607
rect 10137 4573 10171 4607
rect 13817 4573 13851 4607
rect 14001 4573 14035 4607
rect 16301 4573 16335 4607
rect 17773 4573 17807 4607
rect 19245 4573 19279 4607
rect 19337 4573 19371 4607
rect 20625 4573 20659 4607
rect 22281 4573 22315 4607
rect 23661 4573 23695 4607
rect 23753 4573 23787 4607
rect 8849 4505 8883 4539
rect 12253 4505 12287 4539
rect 13265 4505 13299 4539
rect 16761 4505 16795 4539
rect 20165 4505 20199 4539
rect 21637 4505 21671 4539
rect 23017 4505 23051 4539
rect 24949 4505 24983 4539
rect 9217 4437 9251 4471
rect 12621 4437 12655 4471
rect 12713 4437 12747 4471
rect 18601 4437 18635 4471
rect 18785 4437 18819 4471
rect 21269 4437 21303 4471
rect 22649 4437 22683 4471
rect 24673 4437 24707 4471
rect 15289 4233 15323 4267
rect 15933 4233 15967 4267
rect 22189 4233 22223 4267
rect 23201 4233 23235 4267
rect 23937 4233 23971 4267
rect 24949 4233 24983 4267
rect 10137 4165 10171 4199
rect 22649 4165 22683 4199
rect 8113 4097 8147 4131
rect 9677 4097 9711 4131
rect 11609 4097 11643 4131
rect 12805 4097 12839 4131
rect 16301 4097 16335 4131
rect 18325 4097 18359 4131
rect 18877 4097 18911 4131
rect 20257 4097 20291 4131
rect 20717 4097 20751 4131
rect 21729 4097 21763 4131
rect 23753 4097 23787 4131
rect 24581 4097 24615 4131
rect 7101 4029 7135 4063
rect 9493 4029 9527 4063
rect 10965 4029 10999 4063
rect 11885 4029 11919 4063
rect 12529 4029 12563 4063
rect 13909 4029 13943 4063
rect 14176 4029 14210 4063
rect 16393 4029 16427 4063
rect 18233 4029 18267 4063
rect 20993 4029 21027 4063
rect 24305 4029 24339 4063
rect 6549 3961 6583 3995
rect 7377 3961 7411 3995
rect 7929 3961 7963 3995
rect 8021 3961 8055 3995
rect 10781 3961 10815 3995
rect 18141 3961 18175 3995
rect 19521 3961 19555 3995
rect 21637 3961 21671 3995
rect 24397 3961 24431 3995
rect 7561 3893 7595 3927
rect 8665 3893 8699 3927
rect 8941 3893 8975 3927
rect 9125 3893 9159 3927
rect 9585 3893 9619 3927
rect 11149 3893 11183 3927
rect 12161 3893 12195 3927
rect 12621 3893 12655 3927
rect 13357 3893 13391 3927
rect 13817 3893 13851 3927
rect 16577 3893 16611 3927
rect 17129 3893 17163 3927
rect 17497 3893 17531 3927
rect 17773 3893 17807 3927
rect 19613 3893 19647 3927
rect 19981 3893 20015 3927
rect 20073 3893 20107 3927
rect 21177 3893 21211 3927
rect 21545 3893 21579 3927
rect 7653 3689 7687 3723
rect 10781 3689 10815 3723
rect 11333 3689 11367 3723
rect 13265 3689 13299 3723
rect 14001 3689 14035 3723
rect 14369 3689 14403 3723
rect 14829 3689 14863 3723
rect 16025 3689 16059 3723
rect 16577 3689 16611 3723
rect 17037 3689 17071 3723
rect 17681 3689 17715 3723
rect 18141 3689 18175 3723
rect 18601 3689 18635 3723
rect 19981 3689 20015 3723
rect 20441 3689 20475 3723
rect 21177 3689 21211 3723
rect 21913 3689 21947 3723
rect 23201 3689 23235 3723
rect 9668 3621 9702 3655
rect 16945 3621 16979 3655
rect 18509 3621 18543 3655
rect 19153 3621 19187 3655
rect 23560 3621 23594 3655
rect 8205 3553 8239 3587
rect 11885 3553 11919 3587
rect 12152 3553 12186 3587
rect 15381 3553 15415 3587
rect 15473 3553 15507 3587
rect 18049 3553 18083 3587
rect 22281 3553 22315 3587
rect 22649 3553 22683 3587
rect 23293 3553 23327 3587
rect 9401 3485 9435 3519
rect 15565 3485 15599 3519
rect 17221 3485 17255 3519
rect 18693 3485 18727 3519
rect 21269 3485 21303 3519
rect 21361 3485 21395 3519
rect 8389 3349 8423 3383
rect 8757 3349 8791 3383
rect 9217 3349 9251 3383
rect 11793 3349 11827 3383
rect 15013 3349 15047 3383
rect 16485 3349 16519 3383
rect 19613 3349 19647 3383
rect 20809 3349 20843 3383
rect 24673 3349 24707 3383
rect 7745 3145 7779 3179
rect 8849 3145 8883 3179
rect 10689 3145 10723 3179
rect 12437 3145 12471 3179
rect 15381 3145 15415 3179
rect 16393 3145 16427 3179
rect 17405 3145 17439 3179
rect 19153 3145 19187 3179
rect 19705 3145 19739 3179
rect 22097 3145 22131 3179
rect 23201 3145 23235 3179
rect 8113 3077 8147 3111
rect 16669 3077 16703 3111
rect 17037 3077 17071 3111
rect 9217 3009 9251 3043
rect 11609 3009 11643 3043
rect 13081 3009 13115 3043
rect 14001 3009 14035 3043
rect 15933 3009 15967 3043
rect 20257 3009 20291 3043
rect 8205 2941 8239 2975
rect 9309 2941 9343 2975
rect 9576 2941 9610 2975
rect 13449 2941 13483 2975
rect 16485 2941 16519 2975
rect 17773 2941 17807 2975
rect 20524 2941 20558 2975
rect 7193 2873 7227 2907
rect 11885 2873 11919 2907
rect 12805 2873 12839 2907
rect 12897 2873 12931 2907
rect 13909 2873 13943 2907
rect 14246 2873 14280 2907
rect 18018 2873 18052 2907
rect 20165 2873 20199 2907
rect 22833 3009 22867 3043
rect 23937 3009 23971 3043
rect 24397 3009 24431 3043
rect 23753 2941 23787 2975
rect 23845 2873 23879 2907
rect 24857 2873 24891 2907
rect 8389 2805 8423 2839
rect 21637 2805 21671 2839
rect 22097 2805 22131 2839
rect 22281 2805 22315 2839
rect 23385 2805 23419 2839
rect 25133 2805 25167 2839
rect 25593 2805 25627 2839
rect 25869 2805 25903 2839
rect 9309 2601 9343 2635
rect 10689 2601 10723 2635
rect 11793 2601 11827 2635
rect 13725 2601 13759 2635
rect 16577 2601 16611 2635
rect 17221 2601 17255 2635
rect 19429 2601 19463 2635
rect 20717 2601 20751 2635
rect 22281 2601 22315 2635
rect 23753 2601 23787 2635
rect 24213 2601 24247 2635
rect 24765 2601 24799 2635
rect 25777 2601 25811 2635
rect 7009 2533 7043 2567
rect 10229 2533 10263 2567
rect 11149 2533 11183 2567
rect 12161 2533 12195 2567
rect 12612 2533 12646 2567
rect 14645 2533 14679 2567
rect 15013 2533 15047 2567
rect 15464 2533 15498 2567
rect 21146 2533 21180 2567
rect 7377 2465 7411 2499
rect 8205 2465 8239 2499
rect 8941 2465 8975 2499
rect 9585 2465 9619 2499
rect 11057 2465 11091 2499
rect 12345 2465 12379 2499
rect 15197 2465 15231 2499
rect 17865 2465 17899 2499
rect 18316 2465 18350 2499
rect 20901 2465 20935 2499
rect 23017 2465 23051 2499
rect 24121 2465 24155 2499
rect 25133 2465 25167 2499
rect 7745 2397 7779 2431
rect 8297 2397 8331 2431
rect 8481 2397 8515 2431
rect 11333 2397 11367 2431
rect 18049 2397 18083 2431
rect 24305 2397 24339 2431
rect 25317 2397 25351 2431
rect 7837 2329 7871 2363
rect 9769 2261 9803 2295
rect 10505 2261 10539 2295
rect 20257 2261 20291 2295
rect 23477 2261 23511 2295
<< metal1 >>
rect 816 25594 26576 25616
rect 816 25542 10027 25594
rect 10079 25542 10091 25594
rect 10143 25542 10155 25594
rect 10207 25542 10219 25594
rect 10271 25542 19360 25594
rect 19412 25542 19424 25594
rect 19476 25542 19488 25594
rect 19540 25542 19552 25594
rect 19604 25542 26576 25594
rect 816 25520 26576 25542
rect 816 25050 26576 25072
rect 816 24998 5360 25050
rect 5412 24998 5424 25050
rect 5476 24998 5488 25050
rect 5540 24998 5552 25050
rect 5604 24998 14694 25050
rect 14746 24998 14758 25050
rect 14810 24998 14822 25050
rect 14874 24998 14886 25050
rect 14938 24998 24027 25050
rect 24079 24998 24091 25050
rect 24143 24998 24155 25050
rect 24207 24998 24219 25050
rect 24271 24998 26576 25050
rect 816 24976 26576 24998
rect 816 24506 26576 24528
rect 816 24454 10027 24506
rect 10079 24454 10091 24506
rect 10143 24454 10155 24506
rect 10207 24454 10219 24506
rect 10271 24454 19360 24506
rect 19412 24454 19424 24506
rect 19476 24454 19488 24506
rect 19540 24454 19552 24506
rect 19604 24454 26576 24506
rect 816 24432 26576 24454
rect 23833 24395 23891 24401
rect 23833 24361 23845 24395
rect 23879 24392 23891 24395
rect 24842 24392 24848 24404
rect 23879 24364 24848 24392
rect 23879 24361 23891 24364
rect 23833 24355 23891 24361
rect 24842 24352 24848 24364
rect 24900 24352 24906 24404
rect 816 23962 26576 23984
rect 816 23910 5360 23962
rect 5412 23910 5424 23962
rect 5476 23910 5488 23962
rect 5540 23910 5552 23962
rect 5604 23910 14694 23962
rect 14746 23910 14758 23962
rect 14810 23910 14822 23962
rect 14874 23910 14886 23962
rect 14938 23910 24027 23962
rect 24079 23910 24091 23962
rect 24143 23910 24155 23962
rect 24207 23910 24219 23962
rect 24271 23910 26576 23962
rect 816 23888 26576 23910
rect 24474 23848 24480 23860
rect 24435 23820 24480 23848
rect 24474 23808 24480 23820
rect 24532 23808 24538 23860
rect 23646 23604 23652 23656
rect 23704 23644 23710 23656
rect 24293 23647 24351 23653
rect 24293 23644 24305 23647
rect 23704 23616 24305 23644
rect 23704 23604 23710 23616
rect 24293 23613 24305 23616
rect 24339 23644 24351 23647
rect 24845 23647 24903 23653
rect 24845 23644 24857 23647
rect 24339 23616 24857 23644
rect 24339 23613 24351 23616
rect 24293 23607 24351 23613
rect 24845 23613 24857 23616
rect 24891 23613 24903 23647
rect 24845 23607 24903 23613
rect 2486 23468 2492 23520
rect 2544 23508 2550 23520
rect 3774 23508 3780 23520
rect 2544 23480 3780 23508
rect 2544 23468 2550 23480
rect 3774 23468 3780 23480
rect 3832 23468 3838 23520
rect 816 23418 26576 23440
rect 816 23366 10027 23418
rect 10079 23366 10091 23418
rect 10143 23366 10155 23418
rect 10207 23366 10219 23418
rect 10271 23366 19360 23418
rect 19412 23366 19424 23418
rect 19476 23366 19488 23418
rect 19540 23366 19552 23418
rect 19604 23366 26576 23418
rect 816 23344 26576 23366
rect 10674 23304 10680 23316
rect 10635 23276 10680 23304
rect 10674 23264 10680 23276
rect 10732 23264 10738 23316
rect 24474 23304 24480 23316
rect 24435 23276 24480 23304
rect 24474 23264 24480 23276
rect 24532 23264 24538 23316
rect 10490 23168 10496 23180
rect 10451 23140 10496 23168
rect 10490 23128 10496 23140
rect 10548 23128 10554 23180
rect 23830 23128 23836 23180
rect 23888 23168 23894 23180
rect 24293 23171 24351 23177
rect 24293 23168 24305 23171
rect 23888 23140 24305 23168
rect 23888 23128 23894 23140
rect 24293 23137 24305 23140
rect 24339 23137 24351 23171
rect 24293 23131 24351 23137
rect 816 22874 26576 22896
rect 816 22822 5360 22874
rect 5412 22822 5424 22874
rect 5476 22822 5488 22874
rect 5540 22822 5552 22874
rect 5604 22822 14694 22874
rect 14746 22822 14758 22874
rect 14810 22822 14822 22874
rect 14874 22822 14886 22874
rect 14938 22822 24027 22874
rect 24079 22822 24091 22874
rect 24143 22822 24155 22874
rect 24207 22822 24219 22874
rect 24271 22822 26576 22874
rect 816 22800 26576 22822
rect 24566 22720 24572 22772
rect 24624 22760 24630 22772
rect 24845 22763 24903 22769
rect 24845 22760 24857 22763
rect 24624 22732 24857 22760
rect 24624 22720 24630 22732
rect 24845 22729 24857 22732
rect 24891 22729 24903 22763
rect 24845 22723 24903 22729
rect 23646 22624 23652 22636
rect 23607 22596 23652 22624
rect 23646 22584 23652 22596
rect 23704 22584 23710 22636
rect 23373 22559 23431 22565
rect 23373 22556 23385 22559
rect 23204 22528 23385 22556
rect 23204 22500 23232 22528
rect 23373 22525 23385 22528
rect 23419 22525 23431 22559
rect 24658 22556 24664 22568
rect 24619 22528 24664 22556
rect 23373 22519 23431 22525
rect 24658 22516 24664 22528
rect 24716 22556 24722 22568
rect 25213 22559 25271 22565
rect 25213 22556 25225 22559
rect 24716 22528 25225 22556
rect 24716 22516 24722 22528
rect 25213 22525 25225 22528
rect 25259 22525 25271 22559
rect 25213 22519 25271 22525
rect 23186 22488 23192 22500
rect 23147 22460 23192 22488
rect 23186 22448 23192 22460
rect 23244 22448 23250 22500
rect 9754 22380 9760 22432
rect 9812 22420 9818 22432
rect 10490 22420 10496 22432
rect 9812 22392 10496 22420
rect 9812 22380 9818 22392
rect 10490 22380 10496 22392
rect 10548 22380 10554 22432
rect 23830 22380 23836 22432
rect 23888 22420 23894 22432
rect 24382 22420 24388 22432
rect 23888 22392 24388 22420
rect 23888 22380 23894 22392
rect 24382 22380 24388 22392
rect 24440 22380 24446 22432
rect 816 22330 26576 22352
rect 816 22278 10027 22330
rect 10079 22278 10091 22330
rect 10143 22278 10155 22330
rect 10207 22278 10219 22330
rect 10271 22278 19360 22330
rect 19412 22278 19424 22330
rect 19476 22278 19488 22330
rect 19540 22278 19552 22330
rect 19604 22278 26576 22330
rect 816 22256 26576 22278
rect 9754 22148 9760 22160
rect 9715 22120 9760 22148
rect 9754 22108 9760 22120
rect 9812 22108 9818 22160
rect 9386 22040 9392 22092
rect 9444 22080 9450 22092
rect 9481 22083 9539 22089
rect 9481 22080 9493 22083
rect 9444 22052 9493 22080
rect 9444 22040 9450 22052
rect 9481 22049 9493 22052
rect 9527 22049 9539 22083
rect 9481 22043 9539 22049
rect 12149 22083 12207 22089
rect 12149 22049 12161 22083
rect 12195 22080 12207 22083
rect 12330 22080 12336 22092
rect 12195 22052 12336 22080
rect 12195 22049 12207 22052
rect 12149 22043 12207 22049
rect 12330 22040 12336 22052
rect 12388 22040 12394 22092
rect 24293 22083 24351 22089
rect 24293 22049 24305 22083
rect 24339 22080 24351 22083
rect 24382 22080 24388 22092
rect 24339 22052 24388 22080
rect 24339 22049 24351 22052
rect 24293 22043 24351 22049
rect 24382 22040 24388 22052
rect 24440 22040 24446 22092
rect 12422 22012 12428 22024
rect 12383 21984 12428 22012
rect 12422 21972 12428 21984
rect 12480 21972 12486 22024
rect 23738 21904 23744 21956
rect 23796 21944 23802 21956
rect 24477 21947 24535 21953
rect 24477 21944 24489 21947
rect 23796 21916 24489 21944
rect 23796 21904 23802 21916
rect 24477 21913 24489 21916
rect 24523 21913 24535 21947
rect 24477 21907 24535 21913
rect 816 21786 26576 21808
rect 816 21734 5360 21786
rect 5412 21734 5424 21786
rect 5476 21734 5488 21786
rect 5540 21734 5552 21786
rect 5604 21734 14694 21786
rect 14746 21734 14758 21786
rect 14810 21734 14822 21786
rect 14874 21734 14886 21786
rect 14938 21734 24027 21786
rect 24079 21734 24091 21786
rect 24143 21734 24155 21786
rect 24207 21734 24219 21786
rect 24271 21734 26576 21786
rect 816 21712 26576 21734
rect 24474 21672 24480 21684
rect 24435 21644 24480 21672
rect 24474 21632 24480 21644
rect 24532 21632 24538 21684
rect 24382 21536 24388 21548
rect 24124 21508 24388 21536
rect 24124 21480 24152 21508
rect 24382 21496 24388 21508
rect 24440 21496 24446 21548
rect 14722 21468 14728 21480
rect 14683 21440 14728 21468
rect 14722 21428 14728 21440
rect 14780 21468 14786 21480
rect 15461 21471 15519 21477
rect 15461 21468 15473 21471
rect 14780 21440 15473 21468
rect 14780 21428 14786 21440
rect 15461 21437 15473 21440
rect 15507 21437 15519 21471
rect 24106 21468 24112 21480
rect 24067 21440 24112 21468
rect 15461 21431 15519 21437
rect 24106 21428 24112 21440
rect 24164 21428 24170 21480
rect 24290 21468 24296 21480
rect 24203 21440 24296 21468
rect 24290 21428 24296 21440
rect 24348 21468 24354 21480
rect 24845 21471 24903 21477
rect 24845 21468 24857 21471
rect 24348 21440 24857 21468
rect 24348 21428 24354 21440
rect 24845 21437 24857 21440
rect 24891 21437 24903 21471
rect 24845 21431 24903 21437
rect 14998 21400 15004 21412
rect 14959 21372 15004 21400
rect 14998 21360 15004 21372
rect 15056 21360 15062 21412
rect 9386 21292 9392 21344
rect 9444 21332 9450 21344
rect 9481 21335 9539 21341
rect 9481 21332 9493 21335
rect 9444 21304 9493 21332
rect 9444 21292 9450 21304
rect 9481 21301 9493 21304
rect 9527 21301 9539 21335
rect 12330 21332 12336 21344
rect 12291 21304 12336 21332
rect 9481 21295 9539 21301
rect 12330 21292 12336 21304
rect 12388 21292 12394 21344
rect 816 21242 26576 21264
rect 816 21190 10027 21242
rect 10079 21190 10091 21242
rect 10143 21190 10155 21242
rect 10207 21190 10219 21242
rect 10271 21190 19360 21242
rect 19412 21190 19424 21242
rect 19476 21190 19488 21242
rect 19540 21190 19552 21242
rect 19604 21190 26576 21242
rect 816 21168 26576 21190
rect 24750 21128 24756 21140
rect 24711 21100 24756 21128
rect 24750 21088 24756 21100
rect 24808 21088 24814 21140
rect 23557 21063 23615 21069
rect 23557 21029 23569 21063
rect 23603 21060 23615 21063
rect 24290 21060 24296 21072
rect 23603 21032 24296 21060
rect 23603 21029 23615 21032
rect 23557 21023 23615 21029
rect 24290 21020 24296 21032
rect 24348 21020 24354 21072
rect 23186 20952 23192 21004
rect 23244 20992 23250 21004
rect 23281 20995 23339 21001
rect 23281 20992 23293 20995
rect 23244 20964 23293 20992
rect 23244 20952 23250 20964
rect 23281 20961 23293 20964
rect 23327 20961 23339 20995
rect 24566 20992 24572 21004
rect 24527 20964 24572 20992
rect 23281 20955 23339 20961
rect 24566 20952 24572 20964
rect 24624 20952 24630 21004
rect 816 20698 26576 20720
rect 816 20646 5360 20698
rect 5412 20646 5424 20698
rect 5476 20646 5488 20698
rect 5540 20646 5552 20698
rect 5604 20646 14694 20698
rect 14746 20646 14758 20698
rect 14810 20646 14822 20698
rect 14874 20646 14886 20698
rect 14938 20646 24027 20698
rect 24079 20646 24091 20698
rect 24143 20646 24155 20698
rect 24207 20646 24219 20698
rect 24271 20646 26576 20698
rect 816 20624 26576 20646
rect 23554 20584 23560 20596
rect 23515 20556 23560 20584
rect 23554 20544 23560 20556
rect 23612 20544 23618 20596
rect 23186 20380 23192 20392
rect 23147 20352 23192 20380
rect 23186 20340 23192 20352
rect 23244 20340 23250 20392
rect 23370 20380 23376 20392
rect 23283 20352 23376 20380
rect 23370 20340 23376 20352
rect 23428 20380 23434 20392
rect 23925 20383 23983 20389
rect 23925 20380 23937 20383
rect 23428 20352 23937 20380
rect 23428 20340 23434 20352
rect 23925 20349 23937 20352
rect 23971 20349 23983 20383
rect 23925 20343 23983 20349
rect 24566 20244 24572 20256
rect 24527 20216 24572 20244
rect 24566 20204 24572 20216
rect 24624 20204 24630 20256
rect 816 20154 26576 20176
rect 816 20102 10027 20154
rect 10079 20102 10091 20154
rect 10143 20102 10155 20154
rect 10207 20102 10219 20154
rect 10271 20102 19360 20154
rect 19412 20102 19424 20154
rect 19476 20102 19488 20154
rect 19540 20102 19552 20154
rect 19604 20102 26576 20154
rect 816 20080 26576 20102
rect 24382 20000 24388 20052
rect 24440 20040 24446 20052
rect 24477 20043 24535 20049
rect 24477 20040 24489 20043
rect 24440 20012 24489 20040
rect 24440 20000 24446 20012
rect 24477 20009 24489 20012
rect 24523 20009 24535 20043
rect 24477 20003 24535 20009
rect 21438 19972 21444 19984
rect 21399 19944 21444 19972
rect 21438 19932 21444 19944
rect 21496 19932 21502 19984
rect 22729 19975 22787 19981
rect 22729 19941 22741 19975
rect 22775 19972 22787 19975
rect 23370 19972 23376 19984
rect 22775 19944 23376 19972
rect 22775 19941 22787 19944
rect 22729 19935 22787 19941
rect 23370 19932 23376 19944
rect 23428 19932 23434 19984
rect 21162 19904 21168 19916
rect 21123 19876 21168 19904
rect 21162 19864 21168 19876
rect 21220 19864 21226 19916
rect 22450 19904 22456 19916
rect 22411 19876 22456 19904
rect 22450 19864 22456 19876
rect 22508 19864 22514 19916
rect 24293 19907 24351 19913
rect 24293 19873 24305 19907
rect 24339 19904 24351 19907
rect 24382 19904 24388 19916
rect 24339 19876 24388 19904
rect 24339 19873 24351 19876
rect 24293 19867 24351 19873
rect 24382 19864 24388 19876
rect 24440 19864 24446 19916
rect 816 19610 26576 19632
rect 816 19558 5360 19610
rect 5412 19558 5424 19610
rect 5476 19558 5488 19610
rect 5540 19558 5552 19610
rect 5604 19558 14694 19610
rect 14746 19558 14758 19610
rect 14810 19558 14822 19610
rect 14874 19558 14886 19610
rect 14938 19558 24027 19610
rect 24079 19558 24091 19610
rect 24143 19558 24155 19610
rect 24207 19558 24219 19610
rect 24271 19558 26576 19610
rect 816 19536 26576 19558
rect 23646 19252 23652 19304
rect 23704 19292 23710 19304
rect 24293 19295 24351 19301
rect 24293 19292 24305 19295
rect 23704 19264 24305 19292
rect 23704 19252 23710 19264
rect 24293 19261 24305 19264
rect 24339 19292 24351 19295
rect 24845 19295 24903 19301
rect 24845 19292 24857 19295
rect 24339 19264 24857 19292
rect 24339 19261 24351 19264
rect 24293 19255 24351 19261
rect 24845 19261 24857 19264
rect 24891 19261 24903 19295
rect 24845 19255 24903 19261
rect 20610 19116 20616 19168
rect 20668 19156 20674 19168
rect 21162 19156 21168 19168
rect 20668 19128 21168 19156
rect 20668 19116 20674 19128
rect 21162 19116 21168 19128
rect 21220 19116 21226 19168
rect 22450 19156 22456 19168
rect 22411 19128 22456 19156
rect 22450 19116 22456 19128
rect 22508 19116 22514 19168
rect 24106 19156 24112 19168
rect 24067 19128 24112 19156
rect 24106 19116 24112 19128
rect 24164 19156 24170 19168
rect 24382 19156 24388 19168
rect 24164 19128 24388 19156
rect 24164 19116 24170 19128
rect 24382 19116 24388 19128
rect 24440 19116 24446 19168
rect 24474 19116 24480 19168
rect 24532 19156 24538 19168
rect 24532 19128 24577 19156
rect 24532 19116 24538 19128
rect 816 19066 26576 19088
rect 816 19014 10027 19066
rect 10079 19014 10091 19066
rect 10143 19014 10155 19066
rect 10207 19014 10219 19066
rect 10271 19014 19360 19066
rect 19412 19014 19424 19066
rect 19476 19014 19488 19066
rect 19540 19014 19552 19066
rect 19604 19014 26576 19066
rect 816 18992 26576 19014
rect 11134 18952 11140 18964
rect 11095 18924 11140 18952
rect 11134 18912 11140 18924
rect 11192 18912 11198 18964
rect 10766 18776 10772 18828
rect 10824 18816 10830 18828
rect 10953 18819 11011 18825
rect 10953 18816 10965 18819
rect 10824 18788 10965 18816
rect 10824 18776 10830 18788
rect 10953 18785 10965 18788
rect 10999 18785 11011 18819
rect 10953 18779 11011 18785
rect 15366 18776 15372 18828
rect 15424 18816 15430 18828
rect 15461 18819 15519 18825
rect 15461 18816 15473 18819
rect 15424 18788 15473 18816
rect 15424 18776 15430 18788
rect 15461 18785 15473 18788
rect 15507 18785 15519 18819
rect 15734 18816 15740 18828
rect 15695 18788 15740 18816
rect 15461 18779 15519 18785
rect 15734 18776 15740 18788
rect 15792 18776 15798 18828
rect 816 18522 26576 18544
rect 816 18470 5360 18522
rect 5412 18470 5424 18522
rect 5476 18470 5488 18522
rect 5540 18470 5552 18522
rect 5604 18470 14694 18522
rect 14746 18470 14758 18522
rect 14810 18470 14822 18522
rect 14874 18470 14886 18522
rect 14938 18470 24027 18522
rect 24079 18470 24091 18522
rect 24143 18470 24155 18522
rect 24207 18470 24219 18522
rect 24271 18470 26576 18522
rect 816 18448 26576 18470
rect 24842 18408 24848 18420
rect 24803 18380 24848 18408
rect 24842 18368 24848 18380
rect 24900 18368 24906 18420
rect 23646 18272 23652 18284
rect 23607 18244 23652 18272
rect 23646 18232 23652 18244
rect 23704 18232 23710 18284
rect 23186 18164 23192 18216
rect 23244 18204 23250 18216
rect 23373 18207 23431 18213
rect 23373 18204 23385 18207
rect 23244 18176 23385 18204
rect 23244 18164 23250 18176
rect 23373 18173 23385 18176
rect 23419 18204 23431 18207
rect 24109 18207 24167 18213
rect 24109 18204 24121 18207
rect 23419 18176 24121 18204
rect 23419 18173 23431 18176
rect 23373 18167 23431 18173
rect 24109 18173 24121 18176
rect 24155 18173 24167 18207
rect 24658 18204 24664 18216
rect 24619 18176 24664 18204
rect 24109 18167 24167 18173
rect 24658 18164 24664 18176
rect 24716 18204 24722 18216
rect 25213 18207 25271 18213
rect 25213 18204 25225 18207
rect 24716 18176 25225 18204
rect 24716 18164 24722 18176
rect 25213 18173 25225 18176
rect 25259 18173 25271 18207
rect 25213 18167 25271 18173
rect 10766 18028 10772 18080
rect 10824 18068 10830 18080
rect 10953 18071 11011 18077
rect 10953 18068 10965 18071
rect 10824 18040 10965 18068
rect 10824 18028 10830 18040
rect 10953 18037 10965 18040
rect 10999 18037 11011 18071
rect 10953 18031 11011 18037
rect 15366 18028 15372 18080
rect 15424 18068 15430 18080
rect 15461 18071 15519 18077
rect 15461 18068 15473 18071
rect 15424 18040 15473 18068
rect 15424 18028 15430 18040
rect 15461 18037 15473 18040
rect 15507 18037 15519 18071
rect 15461 18031 15519 18037
rect 816 17978 26576 18000
rect 816 17926 10027 17978
rect 10079 17926 10091 17978
rect 10143 17926 10155 17978
rect 10207 17926 10219 17978
rect 10271 17926 19360 17978
rect 19412 17926 19424 17978
rect 19476 17926 19488 17978
rect 19540 17926 19552 17978
rect 19604 17926 26576 17978
rect 816 17904 26576 17926
rect 10309 17799 10367 17805
rect 10309 17765 10321 17799
rect 10355 17796 10367 17799
rect 10674 17796 10680 17808
rect 10355 17768 10680 17796
rect 10355 17765 10367 17768
rect 10309 17759 10367 17765
rect 10674 17756 10680 17768
rect 10732 17756 10738 17808
rect 9846 17688 9852 17740
rect 9904 17728 9910 17740
rect 10033 17731 10091 17737
rect 10033 17728 10045 17731
rect 9904 17700 10045 17728
rect 9904 17688 9910 17700
rect 10033 17697 10045 17700
rect 10079 17697 10091 17731
rect 15826 17728 15832 17740
rect 15787 17700 15832 17728
rect 10033 17691 10091 17697
rect 15826 17688 15832 17700
rect 15884 17688 15890 17740
rect 16010 17592 16016 17604
rect 15971 17564 16016 17592
rect 16010 17552 16016 17564
rect 16068 17552 16074 17604
rect 816 17434 26576 17456
rect 816 17382 5360 17434
rect 5412 17382 5424 17434
rect 5476 17382 5488 17434
rect 5540 17382 5552 17434
rect 5604 17382 14694 17434
rect 14746 17382 14758 17434
rect 14810 17382 14822 17434
rect 14874 17382 14886 17434
rect 14938 17382 24027 17434
rect 24079 17382 24091 17434
rect 24143 17382 24155 17434
rect 24207 17382 24219 17434
rect 24271 17382 26576 17434
rect 816 17360 26576 17382
rect 24382 17280 24388 17332
rect 24440 17320 24446 17332
rect 24477 17323 24535 17329
rect 24477 17320 24489 17323
rect 24440 17292 24489 17320
rect 24440 17280 24446 17292
rect 24477 17289 24489 17292
rect 24523 17289 24535 17323
rect 24477 17283 24535 17289
rect 12146 17076 12152 17128
rect 12204 17116 12210 17128
rect 12609 17119 12667 17125
rect 12609 17116 12621 17119
rect 12204 17088 12621 17116
rect 12204 17076 12210 17088
rect 12609 17085 12621 17088
rect 12655 17116 12667 17119
rect 13345 17119 13403 17125
rect 13345 17116 13357 17119
rect 12655 17088 13357 17116
rect 12655 17085 12667 17088
rect 12609 17079 12667 17085
rect 13345 17085 13357 17088
rect 13391 17085 13403 17119
rect 24290 17116 24296 17128
rect 24251 17088 24296 17116
rect 13345 17079 13403 17085
rect 24290 17076 24296 17088
rect 24348 17116 24354 17128
rect 24845 17119 24903 17125
rect 24845 17116 24857 17119
rect 24348 17088 24857 17116
rect 24348 17076 24354 17088
rect 24845 17085 24857 17088
rect 24891 17085 24903 17119
rect 24845 17079 24903 17085
rect 12882 17048 12888 17060
rect 12843 17020 12888 17048
rect 12882 17008 12888 17020
rect 12940 17008 12946 17060
rect 9846 16940 9852 16992
rect 9904 16980 9910 16992
rect 10033 16983 10091 16989
rect 10033 16980 10045 16983
rect 9904 16952 10045 16980
rect 9904 16940 9910 16952
rect 10033 16949 10045 16952
rect 10079 16949 10091 16983
rect 15826 16980 15832 16992
rect 15787 16952 15832 16980
rect 10033 16943 10091 16949
rect 15826 16940 15832 16952
rect 15884 16940 15890 16992
rect 816 16890 26576 16912
rect 816 16838 10027 16890
rect 10079 16838 10091 16890
rect 10143 16838 10155 16890
rect 10207 16838 10219 16890
rect 10271 16838 19360 16890
rect 19412 16838 19424 16890
rect 19476 16838 19488 16890
rect 19540 16838 19552 16890
rect 19604 16838 26576 16890
rect 816 16816 26576 16838
rect 24474 16776 24480 16788
rect 24435 16748 24480 16776
rect 24474 16736 24480 16748
rect 24532 16736 24538 16788
rect 15277 16711 15335 16717
rect 15277 16677 15289 16711
rect 15323 16708 15335 16711
rect 15826 16708 15832 16720
rect 15323 16680 15832 16708
rect 15323 16677 15335 16680
rect 15277 16671 15335 16677
rect 15826 16668 15832 16680
rect 15884 16668 15890 16720
rect 14998 16640 15004 16652
rect 14959 16612 15004 16640
rect 14998 16600 15004 16612
rect 15056 16600 15062 16652
rect 24293 16643 24351 16649
rect 24293 16609 24305 16643
rect 24339 16640 24351 16643
rect 24382 16640 24388 16652
rect 24339 16612 24388 16640
rect 24339 16609 24351 16612
rect 24293 16603 24351 16609
rect 24382 16600 24388 16612
rect 24440 16600 24446 16652
rect 816 16346 26576 16368
rect 816 16294 5360 16346
rect 5412 16294 5424 16346
rect 5476 16294 5488 16346
rect 5540 16294 5552 16346
rect 5604 16294 14694 16346
rect 14746 16294 14758 16346
rect 14810 16294 14822 16346
rect 14874 16294 14886 16346
rect 14938 16294 24027 16346
rect 24079 16294 24091 16346
rect 24143 16294 24155 16346
rect 24207 16294 24219 16346
rect 24271 16294 26576 16346
rect 816 16272 26576 16294
rect 23830 16192 23836 16244
rect 23888 16232 23894 16244
rect 24477 16235 24535 16241
rect 24477 16232 24489 16235
rect 23888 16204 24489 16232
rect 23888 16192 23894 16204
rect 24477 16201 24489 16204
rect 24523 16201 24535 16235
rect 24477 16195 24535 16201
rect 18218 16096 18224 16108
rect 18179 16068 18224 16096
rect 18218 16056 18224 16068
rect 18276 16056 18282 16108
rect 17945 16031 18003 16037
rect 17945 15997 17957 16031
rect 17991 16028 18003 16031
rect 17991 16000 18816 16028
rect 17991 15997 18003 16000
rect 17945 15991 18003 15997
rect 14998 15892 15004 15904
rect 14959 15864 15004 15892
rect 14998 15852 15004 15864
rect 15056 15852 15062 15904
rect 18788 15901 18816 16000
rect 23830 15988 23836 16040
rect 23888 16028 23894 16040
rect 24293 16031 24351 16037
rect 24293 16028 24305 16031
rect 23888 16000 24305 16028
rect 23888 15988 23894 16000
rect 24293 15997 24305 16000
rect 24339 16028 24351 16031
rect 24845 16031 24903 16037
rect 24845 16028 24857 16031
rect 24339 16000 24857 16028
rect 24339 15997 24351 16000
rect 24293 15991 24351 15997
rect 24845 15997 24857 16000
rect 24891 15997 24903 16031
rect 24845 15991 24903 15997
rect 18773 15895 18831 15901
rect 18773 15861 18785 15895
rect 18819 15892 18831 15895
rect 18862 15892 18868 15904
rect 18819 15864 18868 15892
rect 18819 15861 18831 15864
rect 18773 15855 18831 15861
rect 18862 15852 18868 15864
rect 18920 15852 18926 15904
rect 24106 15892 24112 15904
rect 24067 15864 24112 15892
rect 24106 15852 24112 15864
rect 24164 15892 24170 15904
rect 24382 15892 24388 15904
rect 24164 15864 24388 15892
rect 24164 15852 24170 15864
rect 24382 15852 24388 15864
rect 24440 15852 24446 15904
rect 816 15802 26576 15824
rect 816 15750 10027 15802
rect 10079 15750 10091 15802
rect 10143 15750 10155 15802
rect 10207 15750 10219 15802
rect 10271 15750 19360 15802
rect 19412 15750 19424 15802
rect 19476 15750 19488 15802
rect 19540 15750 19552 15802
rect 19604 15750 26576 15802
rect 816 15728 26576 15750
rect 23373 15623 23431 15629
rect 23373 15589 23385 15623
rect 23419 15620 23431 15623
rect 24106 15620 24112 15632
rect 23419 15592 24112 15620
rect 23419 15589 23431 15592
rect 23373 15583 23431 15589
rect 24106 15580 24112 15592
rect 24164 15580 24170 15632
rect 22726 15512 22732 15564
rect 22784 15552 22790 15564
rect 23097 15555 23155 15561
rect 23097 15552 23109 15555
rect 22784 15524 23109 15552
rect 22784 15512 22790 15524
rect 23097 15521 23109 15524
rect 23143 15521 23155 15555
rect 24382 15552 24388 15564
rect 24343 15524 24388 15552
rect 23097 15515 23155 15521
rect 24382 15512 24388 15524
rect 24440 15512 24446 15564
rect 24569 15351 24627 15357
rect 24569 15317 24581 15351
rect 24615 15348 24627 15351
rect 26314 15348 26320 15360
rect 24615 15320 26320 15348
rect 24615 15317 24627 15320
rect 24569 15311 24627 15317
rect 26314 15308 26320 15320
rect 26372 15308 26378 15360
rect 816 15258 26576 15280
rect 816 15206 5360 15258
rect 5412 15206 5424 15258
rect 5476 15206 5488 15258
rect 5540 15206 5552 15258
rect 5604 15206 14694 15258
rect 14746 15206 14758 15258
rect 14810 15206 14822 15258
rect 14874 15206 14886 15258
rect 14938 15206 24027 15258
rect 24079 15206 24091 15258
rect 24143 15206 24155 15258
rect 24207 15206 24219 15258
rect 24271 15206 26576 15258
rect 816 15184 26576 15206
rect 24382 15144 24388 15156
rect 24343 15116 24388 15144
rect 24382 15104 24388 15116
rect 24440 15104 24446 15156
rect 24566 15104 24572 15156
rect 24624 15144 24630 15156
rect 25029 15147 25087 15153
rect 25029 15144 25041 15147
rect 24624 15116 25041 15144
rect 24624 15104 24630 15116
rect 25029 15113 25041 15116
rect 25075 15113 25087 15147
rect 25029 15107 25087 15113
rect 23830 15008 23836 15020
rect 23791 14980 23836 15008
rect 23830 14968 23836 14980
rect 23888 14968 23894 15020
rect 23189 14943 23247 14949
rect 23189 14909 23201 14943
rect 23235 14940 23247 14943
rect 23554 14940 23560 14952
rect 23235 14912 23560 14940
rect 23235 14909 23247 14912
rect 23189 14903 23247 14909
rect 23554 14900 23560 14912
rect 23612 14900 23618 14952
rect 24842 14940 24848 14952
rect 24803 14912 24848 14940
rect 24842 14900 24848 14912
rect 24900 14940 24906 14952
rect 25397 14943 25455 14949
rect 25397 14940 25409 14943
rect 24900 14912 25409 14940
rect 24900 14900 24906 14912
rect 25397 14909 25409 14912
rect 25443 14909 25455 14943
rect 25397 14903 25455 14909
rect 22726 14804 22732 14816
rect 22687 14776 22732 14804
rect 22726 14764 22732 14776
rect 22784 14764 22790 14816
rect 816 14714 26576 14736
rect 816 14662 10027 14714
rect 10079 14662 10091 14714
rect 10143 14662 10155 14714
rect 10207 14662 10219 14714
rect 10271 14662 19360 14714
rect 19412 14662 19424 14714
rect 19476 14662 19488 14714
rect 19540 14662 19552 14714
rect 19604 14662 26576 14714
rect 816 14640 26576 14662
rect 24569 14603 24627 14609
rect 24569 14569 24581 14603
rect 24615 14600 24627 14603
rect 24658 14600 24664 14612
rect 24615 14572 24664 14600
rect 24615 14569 24627 14572
rect 24569 14563 24627 14569
rect 24658 14560 24664 14572
rect 24716 14560 24722 14612
rect 23373 14535 23431 14541
rect 23373 14501 23385 14535
rect 23419 14532 23431 14535
rect 24842 14532 24848 14544
rect 23419 14504 24848 14532
rect 23419 14501 23431 14504
rect 23373 14495 23431 14501
rect 24842 14492 24848 14504
rect 24900 14492 24906 14544
rect 23094 14464 23100 14476
rect 23055 14436 23100 14464
rect 23094 14424 23100 14436
rect 23152 14424 23158 14476
rect 24382 14464 24388 14476
rect 24343 14436 24388 14464
rect 24382 14424 24388 14436
rect 24440 14424 24446 14476
rect 20613 14399 20671 14405
rect 20613 14365 20625 14399
rect 20659 14396 20671 14399
rect 20978 14396 20984 14408
rect 20659 14368 20984 14396
rect 20659 14365 20671 14368
rect 20613 14359 20671 14365
rect 20978 14356 20984 14368
rect 21036 14356 21042 14408
rect 816 14170 26576 14192
rect 816 14118 5360 14170
rect 5412 14118 5424 14170
rect 5476 14118 5488 14170
rect 5540 14118 5552 14170
rect 5604 14118 14694 14170
rect 14746 14118 14758 14170
rect 14810 14118 14822 14170
rect 14874 14118 14886 14170
rect 14938 14118 24027 14170
rect 24079 14118 24091 14170
rect 24143 14118 24155 14170
rect 24207 14118 24219 14170
rect 24271 14118 26576 14170
rect 816 14096 26576 14118
rect 23462 14016 23468 14068
rect 23520 14056 23526 14068
rect 24477 14059 24535 14065
rect 24477 14056 24489 14059
rect 23520 14028 24489 14056
rect 23520 14016 23526 14028
rect 24477 14025 24489 14028
rect 24523 14025 24535 14059
rect 24477 14019 24535 14025
rect 24842 13988 24848 14000
rect 24803 13960 24848 13988
rect 24842 13948 24848 13960
rect 24900 13948 24906 14000
rect 18586 13920 18592 13932
rect 18547 13892 18592 13920
rect 18586 13880 18592 13892
rect 18644 13880 18650 13932
rect 18313 13855 18371 13861
rect 18313 13821 18325 13855
rect 18359 13852 18371 13855
rect 18770 13852 18776 13864
rect 18359 13824 18776 13852
rect 18359 13821 18371 13824
rect 18313 13815 18371 13821
rect 18770 13812 18776 13824
rect 18828 13852 18834 13864
rect 19049 13855 19107 13861
rect 19049 13852 19061 13855
rect 18828 13824 19061 13852
rect 18828 13812 18834 13824
rect 19049 13821 19061 13824
rect 19095 13821 19107 13855
rect 19049 13815 19107 13821
rect 21806 13812 21812 13864
rect 21864 13852 21870 13864
rect 23094 13852 23100 13864
rect 21864 13824 23100 13852
rect 21864 13812 21870 13824
rect 23094 13812 23100 13824
rect 23152 13812 23158 13864
rect 24293 13855 24351 13861
rect 24293 13852 24305 13855
rect 24124 13824 24305 13852
rect 20153 13719 20211 13725
rect 20153 13685 20165 13719
rect 20199 13716 20211 13719
rect 20426 13716 20432 13728
rect 20199 13688 20432 13716
rect 20199 13685 20211 13688
rect 20153 13679 20211 13685
rect 20426 13676 20432 13688
rect 20484 13676 20490 13728
rect 21898 13716 21904 13728
rect 21859 13688 21904 13716
rect 21898 13676 21904 13688
rect 21956 13676 21962 13728
rect 23646 13676 23652 13728
rect 23704 13716 23710 13728
rect 24124 13725 24152 13824
rect 24293 13821 24305 13824
rect 24339 13821 24351 13855
rect 24293 13815 24351 13821
rect 24109 13719 24167 13725
rect 24109 13716 24121 13719
rect 23704 13688 24121 13716
rect 23704 13676 23710 13688
rect 24109 13685 24121 13688
rect 24155 13685 24167 13719
rect 24109 13679 24167 13685
rect 816 13626 26576 13648
rect 816 13574 10027 13626
rect 10079 13574 10091 13626
rect 10143 13574 10155 13626
rect 10207 13574 10219 13626
rect 10271 13574 19360 13626
rect 19412 13574 19424 13626
rect 19476 13574 19488 13626
rect 19540 13574 19552 13626
rect 19604 13574 26576 13626
rect 816 13552 26576 13574
rect 20610 13512 20616 13524
rect 20571 13484 20616 13512
rect 20610 13472 20616 13484
rect 20668 13472 20674 13524
rect 20978 13512 20984 13524
rect 20939 13484 20984 13512
rect 20978 13472 20984 13484
rect 21036 13472 21042 13524
rect 22913 13515 22971 13521
rect 22913 13481 22925 13515
rect 22959 13512 22971 13515
rect 23186 13512 23192 13524
rect 22959 13484 23192 13512
rect 22959 13481 22971 13484
rect 22913 13475 22971 13481
rect 23186 13472 23192 13484
rect 23244 13472 23250 13524
rect 23278 13472 23284 13524
rect 23336 13512 23342 13524
rect 24477 13515 24535 13521
rect 24477 13512 24489 13515
rect 23336 13484 24489 13512
rect 23336 13472 23342 13484
rect 24477 13481 24489 13484
rect 24523 13481 24535 13515
rect 24477 13475 24535 13481
rect 22821 13379 22879 13385
rect 22821 13345 22833 13379
rect 22867 13376 22879 13379
rect 22910 13376 22916 13388
rect 22867 13348 22916 13376
rect 22867 13345 22879 13348
rect 22821 13339 22879 13345
rect 22910 13336 22916 13348
rect 22968 13336 22974 13388
rect 24293 13379 24351 13385
rect 24293 13345 24305 13379
rect 24339 13376 24351 13379
rect 24382 13376 24388 13388
rect 24339 13348 24388 13376
rect 24339 13345 24351 13348
rect 24293 13339 24351 13345
rect 24382 13336 24388 13348
rect 24440 13336 24446 13388
rect 19230 13308 19236 13320
rect 19191 13280 19236 13308
rect 19230 13268 19236 13280
rect 19288 13268 19294 13320
rect 21073 13311 21131 13317
rect 21073 13277 21085 13311
rect 21119 13277 21131 13311
rect 21073 13271 21131 13277
rect 21257 13311 21315 13317
rect 21257 13277 21269 13311
rect 21303 13308 21315 13311
rect 21346 13308 21352 13320
rect 21303 13280 21352 13308
rect 21303 13277 21315 13280
rect 21257 13271 21315 13277
rect 19049 13175 19107 13181
rect 19049 13141 19061 13175
rect 19095 13172 19107 13175
rect 19414 13172 19420 13184
rect 19095 13144 19420 13172
rect 19095 13141 19107 13144
rect 19049 13135 19107 13141
rect 19414 13132 19420 13144
rect 19472 13132 19478 13184
rect 20429 13175 20487 13181
rect 20429 13141 20441 13175
rect 20475 13172 20487 13175
rect 20518 13172 20524 13184
rect 20475 13144 20524 13172
rect 20475 13141 20487 13144
rect 20429 13135 20487 13141
rect 20518 13132 20524 13144
rect 20576 13172 20582 13184
rect 21088 13172 21116 13271
rect 21346 13268 21352 13280
rect 21404 13268 21410 13320
rect 23094 13308 23100 13320
rect 23055 13280 23100 13308
rect 23094 13268 23100 13280
rect 23152 13268 23158 13320
rect 20576 13144 21116 13172
rect 20576 13132 20582 13144
rect 22174 13132 22180 13184
rect 22232 13172 22238 13184
rect 22453 13175 22511 13181
rect 22453 13172 22465 13175
rect 22232 13144 22465 13172
rect 22232 13132 22238 13144
rect 22453 13141 22465 13144
rect 22499 13141 22511 13175
rect 22453 13135 22511 13141
rect 23370 13132 23376 13184
rect 23428 13172 23434 13184
rect 23465 13175 23523 13181
rect 23465 13172 23477 13175
rect 23428 13144 23477 13172
rect 23428 13132 23434 13144
rect 23465 13141 23477 13144
rect 23511 13141 23523 13175
rect 23465 13135 23523 13141
rect 816 13082 26576 13104
rect 816 13030 5360 13082
rect 5412 13030 5424 13082
rect 5476 13030 5488 13082
rect 5540 13030 5552 13082
rect 5604 13030 14694 13082
rect 14746 13030 14758 13082
rect 14810 13030 14822 13082
rect 14874 13030 14886 13082
rect 14938 13030 24027 13082
rect 24079 13030 24091 13082
rect 24143 13030 24155 13082
rect 24207 13030 24219 13082
rect 24271 13030 26576 13082
rect 816 13008 26576 13030
rect 18954 12968 18960 12980
rect 18915 12940 18960 12968
rect 18954 12928 18960 12940
rect 19012 12928 19018 12980
rect 20978 12928 20984 12980
rect 21036 12968 21042 12980
rect 21533 12971 21591 12977
rect 21533 12968 21545 12971
rect 21036 12940 21545 12968
rect 21036 12928 21042 12940
rect 21533 12937 21545 12940
rect 21579 12937 21591 12971
rect 21533 12931 21591 12937
rect 22545 12971 22603 12977
rect 22545 12937 22557 12971
rect 22591 12968 22603 12971
rect 22821 12971 22879 12977
rect 22821 12968 22833 12971
rect 22591 12940 22833 12968
rect 22591 12937 22603 12940
rect 22545 12931 22603 12937
rect 22821 12937 22833 12940
rect 22867 12968 22879 12971
rect 22910 12968 22916 12980
rect 22867 12940 22916 12968
rect 22867 12937 22879 12940
rect 22821 12931 22879 12937
rect 22910 12928 22916 12940
rect 22968 12928 22974 12980
rect 23186 12968 23192 12980
rect 23147 12940 23192 12968
rect 23186 12928 23192 12940
rect 23244 12928 23250 12980
rect 24842 12968 24848 12980
rect 24803 12940 24848 12968
rect 24842 12928 24848 12940
rect 24900 12928 24906 12980
rect 25302 12968 25308 12980
rect 25263 12940 25308 12968
rect 25302 12928 25308 12940
rect 25360 12928 25366 12980
rect 24290 12900 24296 12912
rect 24251 12872 24296 12900
rect 24290 12860 24296 12872
rect 24348 12860 24354 12912
rect 19138 12792 19144 12844
rect 19196 12832 19202 12844
rect 19414 12832 19420 12844
rect 19196 12804 19420 12832
rect 19196 12792 19202 12804
rect 19414 12792 19420 12804
rect 19472 12792 19478 12844
rect 19509 12835 19567 12841
rect 19509 12801 19521 12835
rect 19555 12801 19567 12835
rect 21162 12832 21168 12844
rect 21123 12804 21168 12832
rect 19509 12795 19567 12801
rect 18497 12767 18555 12773
rect 18497 12733 18509 12767
rect 18543 12764 18555 12767
rect 19524 12764 19552 12795
rect 21162 12792 21168 12804
rect 21220 12832 21226 12844
rect 21901 12835 21959 12841
rect 21901 12832 21913 12835
rect 21220 12804 21913 12832
rect 21220 12792 21226 12804
rect 21901 12801 21913 12804
rect 21947 12801 21959 12835
rect 23646 12832 23652 12844
rect 23607 12804 23652 12832
rect 21901 12795 21959 12801
rect 23646 12792 23652 12804
rect 23704 12792 23710 12844
rect 19782 12764 19788 12776
rect 18543 12736 19788 12764
rect 18543 12733 18555 12736
rect 18497 12727 18555 12733
rect 19782 12724 19788 12736
rect 19840 12724 19846 12776
rect 20061 12767 20119 12773
rect 20061 12733 20073 12767
rect 20107 12764 20119 12767
rect 20981 12767 21039 12773
rect 20981 12764 20993 12767
rect 20107 12736 20993 12764
rect 20107 12733 20119 12736
rect 20061 12727 20119 12733
rect 20981 12733 20993 12736
rect 21027 12764 21039 12767
rect 21070 12764 21076 12776
rect 21027 12736 21076 12764
rect 21027 12733 21039 12736
rect 20981 12727 21039 12733
rect 21070 12724 21076 12736
rect 21128 12724 21134 12776
rect 23370 12764 23376 12776
rect 23331 12736 23376 12764
rect 23370 12724 23376 12736
rect 23428 12724 23434 12776
rect 24661 12767 24719 12773
rect 24661 12733 24673 12767
rect 24707 12764 24719 12767
rect 25302 12764 25308 12776
rect 24707 12736 25308 12764
rect 24707 12733 24719 12736
rect 24661 12727 24719 12733
rect 25302 12724 25308 12736
rect 25360 12724 25366 12776
rect 18586 12656 18592 12708
rect 18644 12696 18650 12708
rect 18773 12699 18831 12705
rect 18773 12696 18785 12699
rect 18644 12668 18785 12696
rect 18644 12656 18650 12668
rect 18773 12665 18785 12668
rect 18819 12696 18831 12699
rect 19325 12699 19383 12705
rect 19325 12696 19337 12699
rect 18819 12668 19337 12696
rect 18819 12665 18831 12668
rect 18773 12659 18831 12665
rect 19325 12665 19337 12668
rect 19371 12665 19383 12699
rect 19325 12659 19383 12665
rect 20429 12699 20487 12705
rect 20429 12665 20441 12699
rect 20475 12696 20487 12699
rect 20889 12699 20947 12705
rect 20889 12696 20901 12699
rect 20475 12668 20901 12696
rect 20475 12665 20487 12668
rect 20429 12659 20487 12665
rect 20889 12665 20901 12668
rect 20935 12696 20947 12699
rect 22545 12699 22603 12705
rect 22545 12696 22557 12699
rect 20935 12668 22557 12696
rect 20935 12665 20947 12668
rect 20889 12659 20947 12665
rect 22545 12665 22557 12668
rect 22591 12665 22603 12699
rect 22545 12659 22603 12665
rect 16470 12588 16476 12640
rect 16528 12628 16534 12640
rect 17945 12631 18003 12637
rect 17945 12628 17957 12631
rect 16528 12600 17957 12628
rect 16528 12588 16534 12600
rect 17945 12597 17957 12600
rect 17991 12597 18003 12631
rect 20518 12628 20524 12640
rect 20479 12600 20524 12628
rect 17945 12591 18003 12597
rect 20518 12588 20524 12600
rect 20576 12588 20582 12640
rect 21806 12588 21812 12640
rect 21864 12628 21870 12640
rect 22269 12631 22327 12637
rect 22269 12628 22281 12631
rect 21864 12600 22281 12628
rect 21864 12588 21870 12600
rect 22269 12597 22281 12600
rect 22315 12597 22327 12631
rect 22269 12591 22327 12597
rect 816 12538 26576 12560
rect 816 12486 10027 12538
rect 10079 12486 10091 12538
rect 10143 12486 10155 12538
rect 10207 12486 10219 12538
rect 10271 12486 19360 12538
rect 19412 12486 19424 12538
rect 19476 12486 19488 12538
rect 19540 12486 19552 12538
rect 19604 12486 26576 12538
rect 816 12464 26576 12486
rect 18494 12384 18500 12436
rect 18552 12424 18558 12436
rect 18862 12424 18868 12436
rect 18552 12396 18868 12424
rect 18552 12384 18558 12396
rect 18862 12384 18868 12396
rect 18920 12384 18926 12436
rect 20429 12427 20487 12433
rect 20429 12393 20441 12427
rect 20475 12424 20487 12427
rect 21346 12424 21352 12436
rect 20475 12396 21352 12424
rect 20475 12393 20487 12396
rect 20429 12387 20487 12393
rect 21346 12384 21352 12396
rect 21404 12384 21410 12436
rect 22634 12424 22640 12436
rect 22547 12396 22640 12424
rect 22634 12384 22640 12396
rect 22692 12424 22698 12436
rect 23094 12424 23100 12436
rect 22692 12396 23100 12424
rect 22692 12384 22698 12396
rect 23094 12384 23100 12396
rect 23152 12424 23158 12436
rect 24477 12427 24535 12433
rect 24477 12424 24489 12427
rect 23152 12396 24489 12424
rect 23152 12384 23158 12396
rect 24477 12393 24489 12396
rect 24523 12393 24535 12427
rect 24477 12387 24535 12393
rect 16654 12356 16660 12368
rect 16615 12328 16660 12356
rect 16654 12316 16660 12328
rect 16712 12316 16718 12368
rect 17850 12316 17856 12368
rect 17908 12365 17914 12368
rect 17908 12359 17972 12365
rect 17908 12325 17926 12359
rect 17960 12325 17972 12359
rect 17908 12319 17972 12325
rect 17908 12316 17914 12319
rect 16378 12288 16384 12300
rect 16339 12260 16384 12288
rect 16378 12248 16384 12260
rect 16436 12248 16442 12300
rect 17577 12291 17635 12297
rect 17577 12257 17589 12291
rect 17623 12288 17635 12291
rect 17669 12291 17727 12297
rect 17669 12288 17681 12291
rect 17623 12260 17681 12288
rect 17623 12257 17635 12260
rect 17577 12251 17635 12257
rect 17669 12257 17681 12260
rect 17715 12288 17727 12291
rect 18678 12288 18684 12300
rect 17715 12260 18684 12288
rect 17715 12257 17727 12260
rect 17669 12251 17727 12257
rect 18678 12248 18684 12260
rect 18736 12248 18742 12300
rect 20880 12291 20938 12297
rect 20880 12257 20892 12291
rect 20926 12288 20938 12291
rect 21162 12288 21168 12300
rect 20926 12260 21168 12288
rect 20926 12257 20938 12260
rect 20880 12251 20938 12257
rect 21162 12248 21168 12260
rect 21220 12248 21226 12300
rect 23364 12291 23422 12297
rect 23364 12288 23376 12291
rect 22008 12260 23376 12288
rect 20613 12223 20671 12229
rect 20613 12189 20625 12223
rect 20659 12189 20671 12223
rect 20613 12183 20671 12189
rect 18862 12044 18868 12096
rect 18920 12084 18926 12096
rect 19049 12087 19107 12093
rect 19049 12084 19061 12087
rect 18920 12056 19061 12084
rect 18920 12044 18926 12056
rect 19049 12053 19061 12056
rect 19095 12053 19107 12087
rect 19049 12047 19107 12053
rect 19598 12044 19604 12096
rect 19656 12084 19662 12096
rect 19693 12087 19751 12093
rect 19693 12084 19705 12087
rect 19656 12056 19705 12084
rect 19656 12044 19662 12056
rect 19693 12053 19705 12056
rect 19739 12084 19751 12087
rect 20628 12084 20656 12183
rect 22008 12164 22036 12260
rect 23364 12257 23376 12260
rect 23410 12288 23422 12291
rect 24750 12288 24756 12300
rect 23410 12260 24756 12288
rect 23410 12257 23422 12260
rect 23364 12251 23422 12257
rect 24750 12248 24756 12260
rect 24808 12248 24814 12300
rect 23097 12223 23155 12229
rect 23097 12220 23109 12223
rect 22928 12192 23109 12220
rect 21990 12152 21996 12164
rect 21903 12124 21996 12152
rect 21990 12112 21996 12124
rect 22048 12112 22054 12164
rect 22082 12084 22088 12096
rect 19739 12056 22088 12084
rect 19739 12053 19751 12056
rect 19693 12047 19751 12053
rect 22082 12044 22088 12056
rect 22140 12084 22146 12096
rect 22928 12093 22956 12192
rect 23097 12189 23109 12192
rect 23143 12189 23155 12223
rect 23097 12183 23155 12189
rect 22913 12087 22971 12093
rect 22913 12084 22925 12087
rect 22140 12056 22925 12084
rect 22140 12044 22146 12056
rect 22913 12053 22925 12056
rect 22959 12053 22971 12087
rect 22913 12047 22971 12053
rect 816 11994 26576 12016
rect 816 11942 5360 11994
rect 5412 11942 5424 11994
rect 5476 11942 5488 11994
rect 5540 11942 5552 11994
rect 5604 11942 14694 11994
rect 14746 11942 14758 11994
rect 14810 11942 14822 11994
rect 14874 11942 14886 11994
rect 14938 11942 24027 11994
rect 24079 11942 24091 11994
rect 24143 11942 24155 11994
rect 24207 11942 24219 11994
rect 24271 11942 26576 11994
rect 816 11920 26576 11942
rect 20981 11883 21039 11889
rect 20981 11849 20993 11883
rect 21027 11880 21039 11883
rect 21162 11880 21168 11892
rect 21027 11852 21168 11880
rect 21027 11849 21039 11852
rect 20981 11843 21039 11849
rect 21162 11840 21168 11852
rect 21220 11880 21226 11892
rect 21533 11883 21591 11889
rect 21533 11880 21545 11883
rect 21220 11852 21545 11880
rect 21220 11840 21226 11852
rect 21533 11849 21545 11852
rect 21579 11849 21591 11883
rect 22818 11880 22824 11892
rect 22779 11852 22824 11880
rect 21533 11843 21591 11849
rect 22818 11840 22824 11852
rect 22876 11840 22882 11892
rect 24474 11880 24480 11892
rect 23848 11852 24480 11880
rect 16378 11772 16384 11824
rect 16436 11812 16442 11824
rect 16473 11815 16531 11821
rect 16473 11812 16485 11815
rect 16436 11784 16485 11812
rect 16436 11772 16442 11784
rect 16473 11781 16485 11784
rect 16519 11812 16531 11815
rect 17761 11815 17819 11821
rect 17761 11812 17773 11815
rect 16519 11784 17773 11812
rect 16519 11781 16531 11784
rect 16473 11775 16531 11781
rect 17761 11781 17773 11784
rect 17807 11781 17819 11815
rect 17761 11775 17819 11781
rect 15918 11744 15924 11756
rect 15108 11716 15924 11744
rect 15108 11685 15136 11716
rect 15918 11704 15924 11716
rect 15976 11704 15982 11756
rect 17850 11704 17856 11756
rect 17908 11744 17914 11756
rect 18313 11747 18371 11753
rect 18313 11744 18325 11747
rect 17908 11716 18325 11744
rect 17908 11704 17914 11716
rect 18313 11713 18325 11716
rect 18359 11744 18371 11747
rect 18773 11747 18831 11753
rect 18773 11744 18785 11747
rect 18359 11716 18785 11744
rect 18359 11713 18371 11716
rect 18313 11707 18371 11713
rect 18773 11713 18785 11716
rect 18819 11713 18831 11747
rect 19598 11744 19604 11756
rect 19559 11716 19604 11744
rect 18773 11707 18831 11713
rect 19598 11704 19604 11716
rect 19656 11704 19662 11756
rect 23848 11753 23876 11852
rect 24474 11840 24480 11852
rect 24532 11840 24538 11892
rect 24750 11880 24756 11892
rect 24711 11852 24756 11880
rect 24750 11840 24756 11852
rect 24808 11840 24814 11892
rect 25118 11880 25124 11892
rect 25079 11852 25124 11880
rect 25118 11840 25124 11852
rect 25176 11840 25182 11892
rect 23833 11747 23891 11753
rect 23833 11713 23845 11747
rect 23879 11713 23891 11747
rect 23833 11707 23891 11713
rect 23922 11704 23928 11756
rect 23980 11744 23986 11756
rect 23980 11716 24025 11744
rect 23980 11704 23986 11716
rect 15093 11679 15151 11685
rect 15093 11645 15105 11679
rect 15139 11645 15151 11679
rect 15093 11639 15151 11645
rect 18678 11636 18684 11688
rect 18736 11676 18742 11688
rect 19616 11676 19644 11704
rect 18736 11648 19644 11676
rect 22177 11679 22235 11685
rect 18736 11636 18742 11648
rect 22177 11645 22189 11679
rect 22223 11676 22235 11679
rect 22818 11676 22824 11688
rect 22223 11648 22824 11676
rect 22223 11645 22235 11648
rect 22177 11639 22235 11645
rect 22818 11636 22824 11648
rect 22876 11636 22882 11688
rect 24934 11676 24940 11688
rect 24895 11648 24940 11676
rect 24934 11636 24940 11648
rect 24992 11676 24998 11688
rect 25489 11679 25547 11685
rect 25489 11676 25501 11679
rect 24992 11648 25501 11676
rect 24992 11636 24998 11648
rect 25489 11645 25501 11648
rect 25535 11645 25547 11679
rect 25489 11639 25547 11645
rect 15369 11611 15427 11617
rect 15369 11577 15381 11611
rect 15415 11608 15427 11611
rect 16010 11608 16016 11620
rect 15415 11580 16016 11608
rect 15415 11577 15427 11580
rect 15369 11571 15427 11577
rect 16010 11568 16016 11580
rect 16068 11568 16074 11620
rect 16657 11611 16715 11617
rect 16657 11577 16669 11611
rect 16703 11608 16715 11611
rect 17485 11611 17543 11617
rect 17485 11608 17497 11611
rect 16703 11580 17497 11608
rect 16703 11577 16715 11580
rect 16657 11571 16715 11577
rect 17485 11577 17497 11580
rect 17531 11608 17543 11611
rect 18129 11611 18187 11617
rect 18129 11608 18141 11611
rect 17531 11580 18141 11608
rect 17531 11577 17543 11580
rect 17485 11571 17543 11577
rect 18129 11577 18141 11580
rect 18175 11577 18187 11611
rect 19846 11611 19904 11617
rect 19846 11608 19858 11611
rect 18129 11571 18187 11577
rect 19708 11580 19858 11608
rect 19708 11552 19736 11580
rect 19846 11577 19858 11580
rect 19892 11577 19904 11611
rect 19846 11571 19904 11577
rect 22910 11568 22916 11620
rect 22968 11608 22974 11620
rect 23741 11611 23799 11617
rect 23741 11608 23753 11611
rect 22968 11580 23753 11608
rect 22968 11568 22974 11580
rect 23204 11552 23232 11580
rect 23741 11577 23753 11580
rect 23787 11577 23799 11611
rect 23741 11571 23799 11577
rect 17209 11543 17267 11549
rect 17209 11509 17221 11543
rect 17255 11540 17267 11543
rect 17850 11540 17856 11552
rect 17255 11512 17856 11540
rect 17255 11509 17267 11512
rect 17209 11503 17267 11509
rect 17850 11500 17856 11512
rect 17908 11500 17914 11552
rect 18221 11543 18279 11549
rect 18221 11509 18233 11543
rect 18267 11540 18279 11543
rect 18310 11540 18316 11552
rect 18267 11512 18316 11540
rect 18267 11509 18279 11512
rect 18221 11503 18279 11509
rect 18310 11500 18316 11512
rect 18368 11500 18374 11552
rect 19509 11543 19567 11549
rect 19509 11509 19521 11543
rect 19555 11540 19567 11543
rect 19690 11540 19696 11552
rect 19555 11512 19696 11540
rect 19555 11509 19567 11512
rect 19509 11503 19567 11509
rect 19690 11500 19696 11512
rect 19748 11500 19754 11552
rect 21993 11543 22051 11549
rect 21993 11509 22005 11543
rect 22039 11540 22051 11543
rect 22082 11540 22088 11552
rect 22039 11512 22088 11540
rect 22039 11509 22051 11512
rect 21993 11503 22051 11509
rect 22082 11500 22088 11512
rect 22140 11500 22146 11552
rect 22358 11540 22364 11552
rect 22319 11512 22364 11540
rect 22358 11500 22364 11512
rect 22416 11500 22422 11552
rect 23186 11540 23192 11552
rect 23147 11512 23192 11540
rect 23186 11500 23192 11512
rect 23244 11500 23250 11552
rect 23370 11540 23376 11552
rect 23331 11512 23376 11540
rect 23370 11500 23376 11512
rect 23428 11500 23434 11552
rect 816 11450 26576 11472
rect 816 11398 10027 11450
rect 10079 11398 10091 11450
rect 10143 11398 10155 11450
rect 10207 11398 10219 11450
rect 10271 11398 19360 11450
rect 19412 11398 19424 11450
rect 19476 11398 19488 11450
rect 19540 11398 19552 11450
rect 19604 11398 26576 11450
rect 816 11376 26576 11398
rect 17850 11336 17856 11348
rect 17811 11308 17856 11336
rect 17850 11296 17856 11308
rect 17908 11296 17914 11348
rect 18954 11336 18960 11348
rect 18915 11308 18960 11336
rect 18954 11296 18960 11308
rect 19012 11296 19018 11348
rect 19046 11296 19052 11348
rect 19104 11336 19110 11348
rect 19230 11336 19236 11348
rect 19104 11308 19236 11336
rect 19104 11296 19110 11308
rect 19230 11296 19236 11308
rect 19288 11336 19294 11348
rect 19325 11339 19383 11345
rect 19325 11336 19337 11339
rect 19288 11308 19337 11336
rect 19288 11296 19294 11308
rect 19325 11305 19337 11308
rect 19371 11305 19383 11339
rect 19325 11299 19383 11305
rect 20426 11296 20432 11348
rect 20484 11336 20490 11348
rect 20981 11339 21039 11345
rect 20981 11336 20993 11339
rect 20484 11308 20993 11336
rect 20484 11296 20490 11308
rect 20981 11305 20993 11308
rect 21027 11305 21039 11339
rect 20981 11299 21039 11305
rect 17390 11268 17396 11280
rect 16488 11240 17396 11268
rect 13618 11200 13624 11212
rect 13579 11172 13624 11200
rect 13618 11160 13624 11172
rect 13676 11160 13682 11212
rect 14998 11200 15004 11212
rect 14959 11172 15004 11200
rect 14998 11160 15004 11172
rect 15056 11160 15062 11212
rect 15274 11200 15280 11212
rect 15235 11172 15280 11200
rect 15274 11160 15280 11172
rect 15332 11160 15338 11212
rect 15826 11200 15832 11212
rect 15739 11172 15832 11200
rect 15826 11160 15832 11172
rect 15884 11200 15890 11212
rect 16488 11209 16516 11240
rect 17390 11228 17396 11240
rect 17448 11228 17454 11280
rect 18862 11268 18868 11280
rect 18823 11240 18868 11268
rect 18862 11228 18868 11240
rect 18920 11228 18926 11280
rect 20518 11228 20524 11280
rect 20576 11268 20582 11280
rect 21073 11271 21131 11277
rect 21073 11268 21085 11271
rect 20576 11240 21085 11268
rect 20576 11228 20582 11240
rect 21073 11237 21085 11240
rect 21119 11237 21131 11271
rect 21073 11231 21131 11237
rect 22536 11271 22594 11277
rect 22536 11237 22548 11271
rect 22582 11268 22594 11271
rect 22634 11268 22640 11280
rect 22582 11240 22640 11268
rect 22582 11237 22594 11240
rect 22536 11231 22594 11237
rect 22634 11228 22640 11240
rect 22692 11228 22698 11280
rect 16473 11203 16531 11209
rect 16473 11200 16485 11203
rect 15884 11172 16485 11200
rect 15884 11160 15890 11172
rect 16473 11169 16485 11172
rect 16519 11169 16531 11203
rect 16473 11163 16531 11169
rect 16562 11160 16568 11212
rect 16620 11200 16626 11212
rect 16729 11203 16787 11209
rect 16729 11200 16741 11203
rect 16620 11172 16741 11200
rect 16620 11160 16626 11172
rect 16729 11169 16741 11172
rect 16775 11169 16787 11203
rect 16729 11163 16787 11169
rect 19417 11203 19475 11209
rect 19417 11169 19429 11203
rect 19463 11200 19475 11203
rect 19874 11200 19880 11212
rect 19463 11172 19880 11200
rect 19463 11169 19475 11172
rect 19417 11163 19475 11169
rect 19874 11160 19880 11172
rect 19932 11160 19938 11212
rect 20061 11203 20119 11209
rect 20061 11169 20073 11203
rect 20107 11200 20119 11203
rect 20429 11203 20487 11209
rect 20429 11200 20441 11203
rect 20107 11172 20441 11200
rect 20107 11169 20119 11172
rect 20061 11163 20119 11169
rect 20429 11169 20441 11172
rect 20475 11200 20487 11203
rect 24753 11203 24811 11209
rect 20475 11172 22128 11200
rect 20475 11169 20487 11172
rect 20429 11163 20487 11169
rect 22100 11144 22128 11172
rect 24753 11169 24765 11203
rect 24799 11200 24811 11203
rect 25394 11200 25400 11212
rect 24799 11172 25400 11200
rect 24799 11169 24811 11172
rect 24753 11163 24811 11169
rect 25394 11160 25400 11172
rect 25452 11160 25458 11212
rect 13710 11092 13716 11144
rect 13768 11132 13774 11144
rect 13805 11135 13863 11141
rect 13805 11132 13817 11135
rect 13768 11104 13817 11132
rect 13768 11092 13774 11104
rect 13805 11101 13817 11104
rect 13851 11101 13863 11135
rect 19506 11132 19512 11144
rect 19467 11104 19512 11132
rect 13805 11095 13863 11101
rect 19506 11092 19512 11104
rect 19564 11092 19570 11144
rect 21162 11092 21168 11144
rect 21220 11132 21226 11144
rect 21257 11135 21315 11141
rect 21257 11132 21269 11135
rect 21220 11104 21269 11132
rect 21220 11092 21226 11104
rect 21257 11101 21269 11104
rect 21303 11132 21315 11135
rect 21990 11132 21996 11144
rect 21303 11104 21996 11132
rect 21303 11101 21315 11104
rect 21257 11095 21315 11101
rect 21990 11092 21996 11104
rect 22048 11092 22054 11144
rect 22082 11092 22088 11144
rect 22140 11132 22146 11144
rect 22269 11135 22327 11141
rect 22269 11132 22281 11135
rect 22140 11104 22281 11132
rect 22140 11092 22146 11104
rect 22269 11101 22281 11104
rect 22315 11101 22327 11135
rect 22269 11095 22327 11101
rect 18310 11024 18316 11076
rect 18368 11064 18374 11076
rect 18405 11067 18463 11073
rect 18405 11064 18417 11067
rect 18368 11036 18417 11064
rect 18368 11024 18374 11036
rect 18405 11033 18417 11036
rect 18451 11033 18463 11067
rect 20610 11064 20616 11076
rect 20571 11036 20616 11064
rect 18405 11027 18463 11033
rect 20610 11024 20616 11036
rect 20668 11024 20674 11076
rect 24934 11064 24940 11076
rect 24895 11036 24940 11064
rect 24934 11024 24940 11036
rect 24992 11024 24998 11076
rect 16197 10999 16255 11005
rect 16197 10965 16209 10999
rect 16243 10996 16255 10999
rect 16654 10996 16660 11008
rect 16243 10968 16660 10996
rect 16243 10965 16255 10968
rect 16197 10959 16255 10965
rect 16654 10956 16660 10968
rect 16712 10956 16718 11008
rect 21809 10999 21867 11005
rect 21809 10965 21821 10999
rect 21855 10996 21867 10999
rect 22266 10996 22272 11008
rect 21855 10968 22272 10996
rect 21855 10965 21867 10968
rect 21809 10959 21867 10965
rect 22266 10956 22272 10968
rect 22324 10996 22330 11008
rect 23649 10999 23707 11005
rect 23649 10996 23661 10999
rect 22324 10968 23661 10996
rect 22324 10956 22330 10968
rect 23649 10965 23661 10968
rect 23695 10965 23707 10999
rect 23649 10959 23707 10965
rect 23922 10956 23928 11008
rect 23980 10996 23986 11008
rect 24293 10999 24351 11005
rect 24293 10996 24305 10999
rect 23980 10968 24305 10996
rect 23980 10956 23986 10968
rect 24293 10965 24305 10968
rect 24339 10996 24351 10999
rect 24750 10996 24756 11008
rect 24339 10968 24756 10996
rect 24339 10965 24351 10968
rect 24293 10959 24351 10965
rect 24750 10956 24756 10968
rect 24808 10956 24814 11008
rect 816 10906 26576 10928
rect 816 10854 5360 10906
rect 5412 10854 5424 10906
rect 5476 10854 5488 10906
rect 5540 10854 5552 10906
rect 5604 10854 14694 10906
rect 14746 10854 14758 10906
rect 14810 10854 14822 10906
rect 14874 10854 14886 10906
rect 14938 10854 24027 10906
rect 24079 10854 24091 10906
rect 24143 10854 24155 10906
rect 24207 10854 24219 10906
rect 24271 10854 26576 10906
rect 816 10832 26576 10854
rect 13345 10795 13403 10801
rect 13345 10761 13357 10795
rect 13391 10792 13403 10795
rect 13434 10792 13440 10804
rect 13391 10764 13440 10792
rect 13391 10761 13403 10764
rect 13345 10755 13403 10761
rect 13434 10752 13440 10764
rect 13492 10752 13498 10804
rect 16102 10792 16108 10804
rect 16063 10764 16108 10792
rect 16102 10752 16108 10764
rect 16160 10752 16166 10804
rect 18681 10795 18739 10801
rect 18681 10761 18693 10795
rect 18727 10792 18739 10795
rect 18954 10792 18960 10804
rect 18727 10764 18960 10792
rect 18727 10761 18739 10764
rect 18681 10755 18739 10761
rect 18954 10752 18960 10764
rect 19012 10752 19018 10804
rect 20426 10752 20432 10804
rect 20484 10792 20490 10804
rect 20705 10795 20763 10801
rect 20705 10792 20717 10795
rect 20484 10764 20717 10792
rect 20484 10752 20490 10764
rect 20705 10761 20717 10764
rect 20751 10761 20763 10795
rect 21162 10792 21168 10804
rect 21123 10764 21168 10792
rect 20705 10755 20763 10761
rect 21162 10752 21168 10764
rect 21220 10752 21226 10804
rect 21625 10795 21683 10801
rect 21625 10761 21637 10795
rect 21671 10792 21683 10795
rect 21898 10792 21904 10804
rect 21671 10764 21904 10792
rect 21671 10761 21683 10764
rect 21625 10755 21683 10761
rect 21898 10752 21904 10764
rect 21956 10752 21962 10804
rect 22634 10752 22640 10804
rect 22692 10792 22698 10804
rect 22729 10795 22787 10801
rect 22729 10792 22741 10795
rect 22692 10764 22741 10792
rect 22692 10752 22698 10764
rect 22729 10761 22741 10764
rect 22775 10761 22787 10795
rect 25394 10792 25400 10804
rect 25355 10764 25400 10792
rect 22729 10755 22787 10761
rect 25394 10752 25400 10764
rect 25452 10752 25458 10804
rect 14173 10727 14231 10733
rect 14173 10693 14185 10727
rect 14219 10724 14231 10727
rect 14998 10724 15004 10736
rect 14219 10696 15004 10724
rect 14219 10693 14231 10696
rect 14173 10687 14231 10693
rect 14998 10684 15004 10696
rect 15056 10724 15062 10736
rect 15185 10727 15243 10733
rect 15185 10724 15197 10727
rect 15056 10696 15197 10724
rect 15056 10684 15062 10696
rect 15185 10693 15197 10696
rect 15231 10693 15243 10727
rect 21714 10724 21720 10736
rect 21675 10696 21720 10724
rect 15185 10687 15243 10693
rect 21714 10684 21720 10696
rect 21772 10684 21778 10736
rect 13713 10659 13771 10665
rect 13713 10625 13725 10659
rect 13759 10656 13771 10659
rect 14722 10656 14728 10668
rect 13759 10628 14728 10656
rect 13759 10625 13771 10628
rect 13713 10619 13771 10625
rect 14722 10616 14728 10628
rect 14780 10616 14786 10668
rect 16654 10656 16660 10668
rect 16615 10628 16660 10656
rect 16654 10616 16660 10628
rect 16712 10656 16718 10668
rect 17666 10656 17672 10668
rect 16712 10628 17672 10656
rect 16712 10616 16718 10628
rect 17666 10616 17672 10628
rect 17724 10616 17730 10668
rect 18678 10616 18684 10668
rect 18736 10656 18742 10668
rect 18773 10659 18831 10665
rect 18773 10656 18785 10659
rect 18736 10628 18785 10656
rect 18736 10616 18742 10628
rect 18773 10625 18785 10628
rect 18819 10625 18831 10659
rect 22266 10656 22272 10668
rect 22227 10628 22272 10656
rect 18773 10619 18831 10625
rect 22266 10616 22272 10628
rect 22324 10656 22330 10668
rect 23097 10659 23155 10665
rect 23097 10656 23109 10659
rect 22324 10628 23109 10656
rect 22324 10616 22330 10628
rect 23097 10625 23109 10628
rect 23143 10656 23155 10659
rect 23143 10628 23508 10656
rect 23143 10625 23155 10628
rect 23097 10619 23155 10625
rect 16013 10591 16071 10597
rect 16013 10557 16025 10591
rect 16059 10588 16071 10591
rect 16470 10588 16476 10600
rect 16059 10560 16476 10588
rect 16059 10557 16071 10560
rect 16013 10551 16071 10557
rect 16470 10548 16476 10560
rect 16528 10548 16534 10600
rect 16562 10548 16568 10600
rect 16620 10588 16626 10600
rect 17117 10591 17175 10597
rect 17117 10588 17129 10591
rect 16620 10560 17129 10588
rect 16620 10548 16626 10560
rect 17117 10557 17129 10560
rect 17163 10557 17175 10591
rect 17117 10551 17175 10557
rect 17390 10548 17396 10600
rect 17448 10588 17454 10600
rect 17577 10591 17635 10597
rect 17577 10588 17589 10591
rect 17448 10560 17589 10588
rect 17448 10548 17454 10560
rect 17577 10557 17589 10560
rect 17623 10588 17635 10591
rect 18696 10588 18724 10616
rect 17623 10560 18724 10588
rect 17623 10557 17635 10560
rect 17577 10551 17635 10557
rect 18862 10548 18868 10600
rect 18920 10588 18926 10600
rect 19029 10591 19087 10597
rect 19029 10588 19041 10591
rect 18920 10560 19041 10588
rect 18920 10548 18926 10560
rect 19029 10557 19041 10560
rect 19075 10557 19087 10591
rect 22174 10588 22180 10600
rect 22135 10560 22180 10588
rect 19029 10551 19087 10557
rect 22174 10548 22180 10560
rect 22232 10548 22238 10600
rect 23278 10548 23284 10600
rect 23336 10588 23342 10600
rect 23373 10591 23431 10597
rect 23373 10588 23385 10591
rect 23336 10560 23385 10588
rect 23336 10548 23342 10560
rect 23373 10557 23385 10560
rect 23419 10557 23431 10591
rect 23480 10588 23508 10628
rect 23629 10591 23687 10597
rect 23629 10588 23641 10591
rect 23480 10560 23641 10588
rect 23373 10551 23431 10557
rect 23629 10557 23641 10560
rect 23675 10557 23687 10591
rect 23629 10551 23687 10557
rect 13894 10480 13900 10532
rect 13952 10520 13958 10532
rect 14081 10523 14139 10529
rect 14081 10520 14093 10523
rect 13952 10492 14093 10520
rect 13952 10480 13958 10492
rect 14081 10489 14093 10492
rect 14127 10520 14139 10523
rect 14541 10523 14599 10529
rect 14541 10520 14553 10523
rect 14127 10492 14553 10520
rect 14127 10489 14139 10492
rect 14081 10483 14139 10489
rect 14541 10489 14553 10492
rect 14587 10489 14599 10523
rect 14541 10483 14599 10489
rect 15645 10523 15703 10529
rect 15645 10489 15657 10523
rect 15691 10520 15703 10523
rect 18313 10523 18371 10529
rect 15691 10492 16608 10520
rect 15691 10489 15703 10492
rect 15645 10483 15703 10489
rect 14354 10412 14360 10464
rect 14412 10452 14418 10464
rect 16580 10461 16608 10492
rect 18313 10489 18325 10523
rect 18359 10520 18371 10523
rect 19506 10520 19512 10532
rect 18359 10492 19512 10520
rect 18359 10489 18371 10492
rect 18313 10483 18371 10489
rect 19506 10480 19512 10492
rect 19564 10520 19570 10532
rect 19564 10492 20196 10520
rect 19564 10480 19570 10492
rect 14633 10455 14691 10461
rect 14633 10452 14645 10455
rect 14412 10424 14645 10452
rect 14412 10412 14418 10424
rect 14633 10421 14645 10424
rect 14679 10421 14691 10455
rect 14633 10415 14691 10421
rect 16565 10455 16623 10461
rect 16565 10421 16577 10455
rect 16611 10452 16623 10455
rect 16654 10452 16660 10464
rect 16611 10424 16660 10452
rect 16611 10421 16623 10424
rect 16565 10415 16623 10421
rect 16654 10412 16660 10424
rect 16712 10412 16718 10464
rect 17758 10452 17764 10464
rect 17719 10424 17764 10452
rect 17758 10412 17764 10424
rect 17816 10412 17822 10464
rect 20168 10461 20196 10492
rect 21898 10480 21904 10532
rect 21956 10520 21962 10532
rect 22085 10523 22143 10529
rect 22085 10520 22097 10523
rect 21956 10492 22097 10520
rect 21956 10480 21962 10492
rect 22085 10489 22097 10492
rect 22131 10489 22143 10523
rect 22085 10483 22143 10489
rect 20153 10455 20211 10461
rect 20153 10421 20165 10455
rect 20199 10421 20211 10455
rect 24750 10452 24756 10464
rect 24711 10424 24756 10452
rect 20153 10415 20211 10421
rect 24750 10412 24756 10424
rect 24808 10412 24814 10464
rect 816 10362 26576 10384
rect 816 10310 10027 10362
rect 10079 10310 10091 10362
rect 10143 10310 10155 10362
rect 10207 10310 10219 10362
rect 10271 10310 19360 10362
rect 19412 10310 19424 10362
rect 19476 10310 19488 10362
rect 19540 10310 19552 10362
rect 19604 10310 26576 10362
rect 816 10288 26576 10310
rect 13894 10248 13900 10260
rect 13855 10220 13900 10248
rect 13894 10208 13900 10220
rect 13952 10208 13958 10260
rect 17390 10248 17396 10260
rect 17351 10220 17396 10248
rect 17390 10208 17396 10220
rect 17448 10208 17454 10260
rect 18865 10251 18923 10257
rect 18865 10217 18877 10251
rect 18911 10248 18923 10251
rect 19874 10248 19880 10260
rect 18911 10220 19880 10248
rect 18911 10217 18923 10220
rect 18865 10211 18923 10217
rect 19874 10208 19880 10220
rect 19932 10208 19938 10260
rect 20429 10251 20487 10257
rect 20429 10217 20441 10251
rect 20475 10248 20487 10251
rect 20518 10248 20524 10260
rect 20475 10220 20524 10248
rect 20475 10217 20487 10220
rect 20429 10211 20487 10217
rect 20518 10208 20524 10220
rect 20576 10208 20582 10260
rect 20797 10251 20855 10257
rect 20797 10217 20809 10251
rect 20843 10248 20855 10251
rect 21622 10248 21628 10260
rect 20843 10220 21628 10248
rect 20843 10217 20855 10220
rect 20797 10211 20855 10217
rect 21622 10208 21628 10220
rect 21680 10208 21686 10260
rect 21901 10251 21959 10257
rect 21901 10217 21913 10251
rect 21947 10248 21959 10251
rect 22174 10248 22180 10260
rect 21947 10220 22180 10248
rect 21947 10217 21959 10220
rect 21901 10211 21959 10217
rect 22174 10208 22180 10220
rect 22232 10208 22238 10260
rect 23189 10251 23247 10257
rect 23189 10217 23201 10251
rect 23235 10248 23247 10251
rect 23370 10248 23376 10260
rect 23235 10220 23376 10248
rect 23235 10217 23247 10220
rect 23189 10211 23247 10217
rect 23370 10208 23376 10220
rect 23428 10208 23434 10260
rect 14722 10140 14728 10192
rect 14780 10180 14786 10192
rect 14998 10180 15004 10192
rect 14780 10152 15004 10180
rect 14780 10140 14786 10152
rect 14998 10140 15004 10152
rect 15056 10180 15062 10192
rect 15338 10183 15396 10189
rect 15338 10180 15350 10183
rect 15056 10152 15350 10180
rect 15056 10140 15062 10152
rect 15338 10149 15350 10152
rect 15384 10149 15396 10183
rect 15338 10143 15396 10149
rect 19138 10140 19144 10192
rect 19196 10180 19202 10192
rect 19325 10183 19383 10189
rect 19325 10180 19337 10183
rect 19196 10152 19337 10180
rect 19196 10140 19202 10152
rect 19325 10149 19337 10152
rect 19371 10149 19383 10183
rect 19325 10143 19383 10149
rect 23548 10183 23606 10189
rect 23548 10149 23560 10183
rect 23594 10180 23606 10183
rect 24750 10180 24756 10192
rect 23594 10152 24756 10180
rect 23594 10149 23606 10152
rect 23548 10143 23606 10149
rect 24750 10140 24756 10152
rect 24808 10140 24814 10192
rect 14817 10115 14875 10121
rect 14817 10081 14829 10115
rect 14863 10112 14875 10115
rect 15090 10112 15096 10124
rect 14863 10084 15096 10112
rect 14863 10081 14875 10084
rect 14817 10075 14875 10081
rect 15090 10072 15096 10084
rect 15148 10112 15154 10124
rect 15826 10112 15832 10124
rect 15148 10084 15832 10112
rect 15148 10072 15154 10084
rect 15826 10072 15832 10084
rect 15884 10072 15890 10124
rect 18773 10115 18831 10121
rect 18773 10081 18785 10115
rect 18819 10112 18831 10115
rect 18862 10112 18868 10124
rect 18819 10084 18868 10112
rect 18819 10081 18831 10084
rect 18773 10075 18831 10081
rect 18862 10072 18868 10084
rect 18920 10072 18926 10124
rect 19046 10072 19052 10124
rect 19104 10112 19110 10124
rect 19233 10115 19291 10121
rect 19233 10112 19245 10115
rect 19104 10084 19245 10112
rect 19104 10072 19110 10084
rect 19233 10081 19245 10084
rect 19279 10081 19291 10115
rect 21162 10112 21168 10124
rect 21123 10084 21168 10112
rect 19233 10075 19291 10081
rect 21162 10072 21168 10084
rect 21220 10072 21226 10124
rect 17850 10044 17856 10056
rect 17811 10016 17856 10044
rect 17850 10004 17856 10016
rect 17908 10004 17914 10056
rect 17574 9936 17580 9988
rect 17632 9976 17638 9988
rect 17761 9979 17819 9985
rect 17761 9976 17773 9979
rect 17632 9948 17773 9976
rect 17632 9936 17638 9948
rect 17761 9945 17773 9948
rect 17807 9976 17819 9979
rect 18880 9976 18908 10072
rect 19417 10047 19475 10053
rect 19417 10013 19429 10047
rect 19463 10013 19475 10047
rect 21254 10044 21260 10056
rect 21215 10016 21260 10044
rect 19417 10007 19475 10013
rect 19432 9976 19460 10007
rect 21254 10004 21260 10016
rect 21312 10004 21318 10056
rect 21441 10047 21499 10053
rect 21441 10013 21453 10047
rect 21487 10044 21499 10047
rect 21714 10044 21720 10056
rect 21487 10016 21720 10044
rect 21487 10013 21499 10016
rect 21441 10007 21499 10013
rect 21714 10004 21720 10016
rect 21772 10004 21778 10056
rect 23278 10044 23284 10056
rect 22744 10016 23284 10044
rect 17807 9948 18816 9976
rect 18880 9948 19460 9976
rect 17807 9945 17819 9948
rect 17761 9939 17819 9945
rect 13618 9908 13624 9920
rect 13579 9880 13624 9908
rect 13618 9868 13624 9880
rect 13676 9868 13682 9920
rect 14354 9908 14360 9920
rect 14315 9880 14360 9908
rect 14354 9868 14360 9880
rect 14412 9868 14418 9920
rect 16473 9911 16531 9917
rect 16473 9877 16485 9911
rect 16519 9908 16531 9911
rect 16562 9908 16568 9920
rect 16519 9880 16568 9908
rect 16519 9877 16531 9880
rect 16473 9871 16531 9877
rect 16562 9868 16568 9880
rect 16620 9868 16626 9920
rect 18310 9908 18316 9920
rect 18271 9880 18316 9908
rect 18310 9868 18316 9880
rect 18368 9868 18374 9920
rect 18788 9908 18816 9948
rect 18954 9908 18960 9920
rect 18788 9880 18960 9908
rect 18954 9868 18960 9880
rect 19012 9868 19018 9920
rect 22266 9908 22272 9920
rect 22227 9880 22272 9908
rect 22266 9868 22272 9880
rect 22324 9908 22330 9920
rect 22744 9917 22772 10016
rect 23278 10004 23284 10016
rect 23336 10004 23342 10056
rect 22729 9911 22787 9917
rect 22729 9908 22741 9911
rect 22324 9880 22741 9908
rect 22324 9868 22330 9880
rect 22729 9877 22741 9880
rect 22775 9877 22787 9911
rect 22729 9871 22787 9877
rect 24474 9868 24480 9920
rect 24532 9908 24538 9920
rect 24661 9911 24719 9917
rect 24661 9908 24673 9911
rect 24532 9880 24673 9908
rect 24532 9868 24538 9880
rect 24661 9877 24673 9880
rect 24707 9877 24719 9911
rect 24661 9871 24719 9877
rect 816 9818 26576 9840
rect 816 9766 5360 9818
rect 5412 9766 5424 9818
rect 5476 9766 5488 9818
rect 5540 9766 5552 9818
rect 5604 9766 14694 9818
rect 14746 9766 14758 9818
rect 14810 9766 14822 9818
rect 14874 9766 14886 9818
rect 14938 9766 24027 9818
rect 24079 9766 24091 9818
rect 24143 9766 24155 9818
rect 24207 9766 24219 9818
rect 24271 9766 26576 9818
rect 816 9744 26576 9766
rect 14998 9704 15004 9716
rect 14959 9676 15004 9704
rect 14998 9664 15004 9676
rect 15056 9704 15062 9716
rect 15553 9707 15611 9713
rect 15553 9704 15565 9707
rect 15056 9676 15565 9704
rect 15056 9664 15062 9676
rect 15553 9673 15565 9676
rect 15599 9673 15611 9707
rect 15553 9667 15611 9673
rect 16654 9664 16660 9716
rect 16712 9704 16718 9716
rect 24750 9704 24756 9716
rect 16712 9676 17620 9704
rect 24711 9676 24756 9704
rect 16712 9664 16718 9676
rect 16105 9639 16163 9645
rect 16105 9605 16117 9639
rect 16151 9636 16163 9639
rect 16194 9636 16200 9648
rect 16151 9608 16200 9636
rect 16151 9605 16163 9608
rect 16105 9599 16163 9605
rect 16194 9596 16200 9608
rect 16252 9596 16258 9648
rect 17592 9636 17620 9676
rect 24750 9664 24756 9676
rect 24808 9664 24814 9716
rect 17761 9639 17819 9645
rect 17761 9636 17773 9639
rect 17592 9608 17773 9636
rect 17761 9605 17773 9608
rect 17807 9605 17819 9639
rect 17761 9599 17819 9605
rect 18310 9596 18316 9648
rect 18368 9596 18374 9648
rect 21073 9639 21131 9645
rect 21073 9605 21085 9639
rect 21119 9636 21131 9639
rect 21346 9636 21352 9648
rect 21119 9608 21352 9636
rect 21119 9605 21131 9608
rect 21073 9599 21131 9605
rect 21346 9596 21352 9608
rect 21404 9596 21410 9648
rect 22818 9636 22824 9648
rect 22779 9608 22824 9636
rect 22818 9596 22824 9608
rect 22876 9596 22882 9648
rect 23370 9596 23376 9648
rect 23428 9636 23434 9648
rect 24474 9636 24480 9648
rect 23428 9608 23876 9636
rect 23428 9596 23434 9608
rect 13618 9568 13624 9580
rect 13579 9540 13624 9568
rect 13618 9528 13624 9540
rect 13676 9528 13682 9580
rect 16562 9528 16568 9580
rect 16620 9568 16626 9580
rect 16657 9571 16715 9577
rect 16657 9568 16669 9571
rect 16620 9540 16669 9568
rect 16620 9528 16626 9540
rect 16657 9537 16669 9540
rect 16703 9537 16715 9571
rect 16657 9531 16715 9537
rect 17942 9528 17948 9580
rect 18000 9568 18006 9580
rect 18328 9568 18356 9596
rect 18405 9571 18463 9577
rect 18405 9568 18417 9571
rect 18000 9540 18417 9568
rect 18000 9528 18006 9540
rect 18405 9537 18417 9540
rect 18451 9537 18463 9571
rect 18405 9531 18463 9537
rect 18954 9460 18960 9512
rect 19012 9500 19018 9512
rect 19509 9503 19567 9509
rect 19509 9500 19521 9503
rect 19012 9472 19521 9500
rect 19012 9460 19018 9472
rect 19509 9469 19521 9472
rect 19555 9500 19567 9503
rect 19598 9500 19604 9512
rect 19555 9472 19604 9500
rect 19555 9469 19567 9472
rect 19509 9463 19567 9469
rect 19598 9460 19604 9472
rect 19656 9460 19662 9512
rect 19693 9503 19751 9509
rect 19693 9469 19705 9503
rect 19739 9469 19751 9503
rect 19693 9463 19751 9469
rect 13526 9432 13532 9444
rect 13439 9404 13532 9432
rect 13526 9392 13532 9404
rect 13584 9432 13590 9444
rect 13866 9435 13924 9441
rect 13866 9432 13878 9435
rect 13584 9404 13878 9432
rect 13584 9392 13590 9404
rect 13866 9401 13878 9404
rect 13912 9401 13924 9435
rect 17482 9432 17488 9444
rect 17443 9404 17488 9432
rect 13866 9395 13924 9401
rect 17482 9392 17488 9404
rect 17540 9432 17546 9444
rect 18129 9435 18187 9441
rect 18129 9432 18141 9435
rect 17540 9404 18141 9432
rect 17540 9392 17546 9404
rect 18129 9401 18141 9404
rect 18175 9401 18187 9435
rect 18129 9395 18187 9401
rect 18586 9392 18592 9444
rect 18644 9432 18650 9444
rect 19708 9432 19736 9463
rect 19782 9460 19788 9512
rect 19840 9500 19846 9512
rect 19949 9503 20007 9509
rect 19949 9500 19961 9503
rect 19840 9472 19961 9500
rect 19840 9460 19846 9472
rect 19949 9469 19961 9472
rect 19995 9469 20007 9503
rect 19949 9463 20007 9469
rect 22177 9503 22235 9509
rect 22177 9469 22189 9503
rect 22223 9500 22235 9503
rect 22836 9500 22864 9596
rect 23186 9568 23192 9580
rect 23147 9540 23192 9568
rect 23186 9528 23192 9540
rect 23244 9568 23250 9580
rect 23738 9568 23744 9580
rect 23244 9540 23744 9568
rect 23244 9528 23250 9540
rect 23738 9528 23744 9540
rect 23796 9528 23802 9580
rect 23848 9577 23876 9608
rect 24032 9608 24480 9636
rect 24032 9580 24060 9608
rect 24474 9596 24480 9608
rect 24532 9596 24538 9648
rect 23833 9571 23891 9577
rect 23833 9537 23845 9571
rect 23879 9537 23891 9571
rect 24014 9568 24020 9580
rect 23927 9540 24020 9568
rect 23833 9531 23891 9537
rect 24014 9528 24020 9540
rect 24072 9528 24078 9580
rect 24937 9503 24995 9509
rect 24937 9500 24949 9503
rect 22223 9472 22864 9500
rect 23388 9472 24949 9500
rect 22223 9469 22235 9472
rect 22177 9463 22235 9469
rect 20334 9432 20340 9444
rect 18644 9404 20340 9432
rect 18644 9392 18650 9404
rect 10950 9324 10956 9376
rect 11008 9364 11014 9376
rect 11045 9367 11103 9373
rect 11045 9364 11057 9367
rect 11008 9336 11057 9364
rect 11008 9324 11014 9336
rect 11045 9333 11057 9336
rect 11091 9333 11103 9367
rect 12606 9364 12612 9376
rect 12567 9336 12612 9364
rect 11045 9327 11103 9333
rect 12606 9324 12612 9336
rect 12664 9324 12670 9376
rect 15918 9364 15924 9376
rect 15879 9336 15924 9364
rect 15918 9324 15924 9336
rect 15976 9364 15982 9376
rect 16473 9367 16531 9373
rect 16473 9364 16485 9367
rect 15976 9336 16485 9364
rect 15976 9324 15982 9336
rect 16473 9333 16485 9336
rect 16519 9333 16531 9367
rect 16473 9327 16531 9333
rect 16565 9367 16623 9373
rect 16565 9333 16577 9367
rect 16611 9364 16623 9367
rect 16654 9364 16660 9376
rect 16611 9336 16660 9364
rect 16611 9333 16623 9336
rect 16565 9327 16623 9333
rect 16654 9324 16660 9336
rect 16712 9364 16718 9376
rect 17209 9367 17267 9373
rect 17209 9364 17221 9367
rect 16712 9336 17221 9364
rect 16712 9324 16718 9336
rect 17209 9333 17221 9336
rect 17255 9364 17267 9367
rect 18218 9364 18224 9376
rect 17255 9336 18224 9364
rect 17255 9333 17267 9336
rect 17209 9327 17267 9333
rect 18218 9324 18224 9336
rect 18276 9324 18282 9376
rect 18310 9324 18316 9376
rect 18368 9364 18374 9376
rect 18494 9364 18500 9376
rect 18368 9336 18500 9364
rect 18368 9324 18374 9336
rect 18494 9324 18500 9336
rect 18552 9324 18558 9376
rect 18862 9364 18868 9376
rect 18823 9336 18868 9364
rect 18862 9324 18868 9336
rect 18920 9324 18926 9376
rect 19340 9373 19368 9404
rect 20334 9392 20340 9404
rect 20392 9392 20398 9444
rect 21254 9392 21260 9444
rect 21312 9432 21318 9444
rect 21993 9435 22051 9441
rect 21993 9432 22005 9435
rect 21312 9404 22005 9432
rect 21312 9392 21318 9404
rect 21993 9401 22005 9404
rect 22039 9401 22051 9435
rect 21993 9395 22051 9401
rect 19325 9367 19383 9373
rect 19325 9333 19337 9367
rect 19371 9333 19383 9367
rect 21714 9364 21720 9376
rect 21675 9336 21720 9364
rect 19325 9327 19383 9333
rect 21714 9324 21720 9336
rect 21772 9324 21778 9376
rect 22358 9364 22364 9376
rect 22319 9336 22364 9364
rect 22358 9324 22364 9336
rect 22416 9324 22422 9376
rect 23388 9373 23416 9472
rect 24937 9469 24949 9472
rect 24983 9500 24995 9503
rect 25673 9503 25731 9509
rect 25673 9500 25685 9503
rect 24983 9472 25685 9500
rect 24983 9469 24995 9472
rect 24937 9463 24995 9469
rect 25673 9469 25685 9472
rect 25719 9469 25731 9503
rect 25673 9463 25731 9469
rect 23738 9432 23744 9444
rect 23699 9404 23744 9432
rect 23738 9392 23744 9404
rect 23796 9392 23802 9444
rect 25213 9435 25271 9441
rect 25213 9401 25225 9435
rect 25259 9401 25271 9435
rect 25213 9395 25271 9401
rect 23373 9367 23431 9373
rect 23373 9333 23385 9367
rect 23419 9333 23431 9367
rect 23373 9327 23431 9333
rect 23462 9324 23468 9376
rect 23520 9364 23526 9376
rect 25228 9364 25256 9395
rect 23520 9336 25256 9364
rect 23520 9324 23526 9336
rect 816 9274 26576 9296
rect 816 9222 10027 9274
rect 10079 9222 10091 9274
rect 10143 9222 10155 9274
rect 10207 9222 10219 9274
rect 10271 9222 19360 9274
rect 19412 9222 19424 9274
rect 19476 9222 19488 9274
rect 19540 9222 19552 9274
rect 19604 9222 26576 9274
rect 816 9200 26576 9222
rect 10582 9160 10588 9172
rect 10543 9132 10588 9160
rect 10582 9120 10588 9132
rect 10640 9120 10646 9172
rect 13526 9160 13532 9172
rect 12256 9132 12560 9160
rect 13487 9132 13532 9160
rect 12057 9095 12115 9101
rect 12057 9061 12069 9095
rect 12103 9092 12115 9095
rect 12256 9092 12284 9132
rect 12103 9064 12284 9092
rect 12103 9061 12115 9064
rect 12057 9055 12115 9061
rect 10950 9024 10956 9036
rect 10911 8996 10956 9024
rect 10950 8984 10956 8996
rect 11008 8984 11014 9036
rect 11045 8959 11103 8965
rect 11045 8925 11057 8959
rect 11091 8925 11103 8959
rect 11045 8919 11103 8925
rect 11229 8959 11287 8965
rect 11229 8925 11241 8959
rect 11275 8956 11287 8959
rect 11778 8956 11784 8968
rect 11275 8928 11784 8956
rect 11275 8925 11287 8928
rect 11229 8919 11287 8925
rect 10490 8820 10496 8832
rect 10451 8792 10496 8820
rect 10490 8780 10496 8792
rect 10548 8820 10554 8832
rect 11060 8820 11088 8919
rect 11778 8916 11784 8928
rect 11836 8916 11842 8968
rect 12054 8916 12060 8968
rect 12112 8956 12118 8968
rect 12164 8965 12192 9064
rect 12330 9052 12336 9104
rect 12388 9101 12394 9104
rect 12388 9095 12452 9101
rect 12388 9061 12406 9095
rect 12440 9061 12452 9095
rect 12532 9092 12560 9132
rect 13526 9120 13532 9132
rect 13584 9160 13590 9172
rect 14078 9160 14084 9172
rect 13584 9132 14084 9160
rect 13584 9120 13590 9132
rect 14078 9120 14084 9132
rect 14136 9120 14142 9172
rect 15001 9163 15059 9169
rect 15001 9129 15013 9163
rect 15047 9160 15059 9163
rect 15366 9160 15372 9172
rect 15047 9132 15372 9160
rect 15047 9129 15059 9132
rect 15001 9123 15059 9129
rect 15366 9120 15372 9132
rect 15424 9120 15430 9172
rect 16562 9160 16568 9172
rect 16523 9132 16568 9160
rect 16562 9120 16568 9132
rect 16620 9120 16626 9172
rect 17025 9163 17083 9169
rect 17025 9129 17037 9163
rect 17071 9160 17083 9163
rect 17482 9160 17488 9172
rect 17071 9132 17488 9160
rect 17071 9129 17083 9132
rect 17025 9123 17083 9129
rect 17482 9120 17488 9132
rect 17540 9120 17546 9172
rect 17666 9120 17672 9172
rect 17724 9160 17730 9172
rect 18494 9160 18500 9172
rect 17724 9132 18500 9160
rect 17724 9120 17730 9132
rect 18494 9120 18500 9132
rect 18552 9160 18558 9172
rect 18681 9163 18739 9169
rect 18681 9160 18693 9163
rect 18552 9132 18693 9160
rect 18552 9120 18558 9132
rect 18681 9129 18693 9132
rect 18727 9129 18739 9163
rect 19782 9160 19788 9172
rect 19743 9132 19788 9160
rect 18681 9123 18739 9129
rect 19782 9120 19788 9132
rect 19840 9120 19846 9172
rect 20429 9163 20487 9169
rect 20429 9129 20441 9163
rect 20475 9160 20487 9163
rect 20613 9163 20671 9169
rect 20613 9160 20625 9163
rect 20475 9132 20625 9160
rect 20475 9129 20487 9132
rect 20429 9123 20487 9129
rect 20613 9129 20625 9132
rect 20659 9160 20671 9163
rect 21162 9160 21168 9172
rect 20659 9132 21168 9160
rect 20659 9129 20671 9132
rect 20613 9123 20671 9129
rect 21162 9120 21168 9132
rect 21220 9120 21226 9172
rect 21806 9120 21812 9172
rect 21864 9160 21870 9172
rect 21864 9132 21909 9160
rect 21864 9120 21870 9132
rect 13618 9092 13624 9104
rect 12532 9064 13624 9092
rect 12388 9055 12452 9061
rect 12388 9052 12394 9055
rect 13618 9052 13624 9064
rect 13676 9052 13682 9104
rect 14817 9095 14875 9101
rect 14817 9061 14829 9095
rect 14863 9092 14875 9095
rect 16197 9095 16255 9101
rect 14863 9064 15504 9092
rect 14863 9061 14875 9064
rect 14817 9055 14875 9061
rect 15476 9036 15504 9064
rect 16197 9061 16209 9095
rect 16243 9092 16255 9095
rect 16654 9092 16660 9104
rect 16243 9064 16660 9092
rect 16243 9061 16255 9064
rect 16197 9055 16255 9061
rect 16654 9052 16660 9064
rect 16712 9052 16718 9104
rect 17390 9052 17396 9104
rect 17448 9092 17454 9104
rect 17568 9095 17626 9101
rect 17568 9092 17580 9095
rect 17448 9064 17580 9092
rect 17448 9052 17454 9064
rect 17568 9061 17580 9064
rect 17614 9092 17626 9095
rect 17942 9092 17948 9104
rect 17614 9064 17948 9092
rect 17614 9061 17626 9064
rect 17568 9055 17626 9061
rect 17942 9052 17948 9064
rect 18000 9052 18006 9104
rect 23186 9052 23192 9104
rect 23244 9092 23250 9104
rect 23364 9095 23422 9101
rect 23364 9092 23376 9095
rect 23244 9064 23376 9092
rect 23244 9052 23250 9064
rect 23364 9061 23376 9064
rect 23410 9092 23422 9095
rect 24014 9092 24020 9104
rect 23410 9064 24020 9092
rect 23410 9061 23422 9064
rect 23364 9055 23422 9061
rect 24014 9052 24020 9064
rect 24072 9052 24078 9104
rect 15366 9024 15372 9036
rect 15327 8996 15372 9024
rect 15366 8984 15372 8996
rect 15424 8984 15430 9036
rect 15458 8984 15464 9036
rect 15516 9024 15522 9036
rect 15516 8996 15561 9024
rect 15516 8984 15522 8996
rect 16746 8984 16752 9036
rect 16804 9024 16810 9036
rect 17209 9027 17267 9033
rect 17209 9024 17221 9027
rect 16804 8996 17221 9024
rect 16804 8984 16810 8996
rect 17209 8993 17221 8996
rect 17255 8993 17267 9027
rect 20978 9024 20984 9036
rect 20939 8996 20984 9024
rect 17209 8987 17267 8993
rect 20978 8984 20984 8996
rect 21036 8984 21042 9036
rect 12149 8959 12207 8965
rect 12149 8956 12161 8959
rect 12112 8928 12161 8956
rect 12112 8916 12118 8928
rect 12149 8925 12161 8928
rect 12195 8925 12207 8959
rect 15550 8956 15556 8968
rect 15511 8928 15556 8956
rect 12149 8919 12207 8925
rect 15550 8916 15556 8928
rect 15608 8916 15614 8968
rect 17301 8959 17359 8965
rect 17301 8925 17313 8959
rect 17347 8925 17359 8959
rect 17301 8919 17359 8925
rect 16933 8891 16991 8897
rect 16933 8857 16945 8891
rect 16979 8888 16991 8891
rect 17206 8888 17212 8900
rect 16979 8860 17212 8888
rect 16979 8857 16991 8860
rect 16933 8851 16991 8857
rect 17206 8848 17212 8860
rect 17264 8888 17270 8900
rect 17316 8888 17344 8919
rect 20610 8916 20616 8968
rect 20668 8956 20674 8968
rect 21073 8959 21131 8965
rect 21073 8956 21085 8959
rect 20668 8928 21085 8956
rect 20668 8916 20674 8928
rect 21073 8925 21085 8928
rect 21119 8925 21131 8959
rect 21073 8919 21131 8925
rect 21165 8959 21223 8965
rect 21165 8925 21177 8959
rect 21211 8925 21223 8959
rect 21165 8919 21223 8925
rect 23097 8959 23155 8965
rect 23097 8925 23109 8959
rect 23143 8925 23155 8959
rect 23097 8919 23155 8925
rect 17264 8860 17344 8888
rect 17264 8848 17270 8860
rect 20794 8848 20800 8900
rect 20852 8888 20858 8900
rect 21180 8888 21208 8919
rect 20852 8860 21208 8888
rect 20852 8848 20858 8860
rect 21622 8848 21628 8900
rect 21680 8888 21686 8900
rect 22266 8888 22272 8900
rect 21680 8860 22272 8888
rect 21680 8848 21686 8860
rect 22266 8848 22272 8860
rect 22324 8888 22330 8900
rect 22324 8860 22680 8888
rect 22324 8848 22330 8860
rect 10548 8792 11088 8820
rect 10548 8780 10554 8792
rect 19138 8780 19144 8832
rect 19196 8820 19202 8832
rect 19325 8823 19383 8829
rect 19325 8820 19337 8823
rect 19196 8792 19337 8820
rect 19196 8780 19202 8792
rect 19325 8789 19337 8792
rect 19371 8820 19383 8823
rect 20886 8820 20892 8832
rect 19371 8792 20892 8820
rect 19371 8789 19383 8792
rect 19325 8783 19383 8789
rect 20886 8780 20892 8792
rect 20944 8780 20950 8832
rect 22174 8820 22180 8832
rect 22135 8792 22180 8820
rect 22174 8780 22180 8792
rect 22232 8780 22238 8832
rect 22652 8829 22680 8860
rect 22637 8823 22695 8829
rect 22637 8789 22649 8823
rect 22683 8820 22695 8823
rect 23005 8823 23063 8829
rect 23005 8820 23017 8823
rect 22683 8792 23017 8820
rect 22683 8789 22695 8792
rect 22637 8783 22695 8789
rect 23005 8789 23017 8792
rect 23051 8820 23063 8823
rect 23112 8820 23140 8919
rect 23370 8820 23376 8832
rect 23051 8792 23376 8820
rect 23051 8789 23063 8792
rect 23005 8783 23063 8789
rect 23370 8780 23376 8792
rect 23428 8780 23434 8832
rect 23738 8780 23744 8832
rect 23796 8820 23802 8832
rect 24477 8823 24535 8829
rect 24477 8820 24489 8823
rect 23796 8792 24489 8820
rect 23796 8780 23802 8792
rect 24477 8789 24489 8792
rect 24523 8789 24535 8823
rect 24477 8783 24535 8789
rect 24658 8780 24664 8832
rect 24716 8820 24722 8832
rect 25029 8823 25087 8829
rect 25029 8820 25041 8823
rect 24716 8792 25041 8820
rect 24716 8780 24722 8792
rect 25029 8789 25041 8792
rect 25075 8789 25087 8823
rect 25029 8783 25087 8789
rect 816 8730 26576 8752
rect 816 8678 5360 8730
rect 5412 8678 5424 8730
rect 5476 8678 5488 8730
rect 5540 8678 5552 8730
rect 5604 8678 14694 8730
rect 14746 8678 14758 8730
rect 14810 8678 14822 8730
rect 14874 8678 14886 8730
rect 14938 8678 24027 8730
rect 24079 8678 24091 8730
rect 24143 8678 24155 8730
rect 24207 8678 24219 8730
rect 24271 8678 26576 8730
rect 816 8656 26576 8678
rect 10950 8576 10956 8628
rect 11008 8616 11014 8628
rect 11413 8619 11471 8625
rect 11413 8616 11425 8619
rect 11008 8588 11425 8616
rect 11008 8576 11014 8588
rect 11413 8585 11425 8588
rect 11459 8585 11471 8619
rect 11778 8616 11784 8628
rect 11739 8588 11784 8616
rect 11413 8579 11471 8585
rect 11778 8576 11784 8588
rect 11836 8616 11842 8628
rect 12330 8616 12336 8628
rect 11836 8588 12336 8616
rect 11836 8576 11842 8588
rect 12330 8576 12336 8588
rect 12388 8616 12394 8628
rect 12609 8619 12667 8625
rect 12609 8616 12621 8619
rect 12388 8588 12621 8616
rect 12388 8576 12394 8588
rect 12609 8585 12621 8588
rect 12655 8585 12667 8619
rect 12609 8579 12667 8585
rect 13529 8619 13587 8625
rect 13529 8585 13541 8619
rect 13575 8616 13587 8619
rect 14354 8616 14360 8628
rect 13575 8588 14360 8616
rect 13575 8585 13587 8588
rect 13529 8579 13587 8585
rect 14354 8576 14360 8588
rect 14412 8576 14418 8628
rect 15093 8619 15151 8625
rect 15093 8585 15105 8619
rect 15139 8616 15151 8619
rect 15366 8616 15372 8628
rect 15139 8588 15372 8616
rect 15139 8585 15151 8588
rect 15093 8579 15151 8585
rect 15366 8576 15372 8588
rect 15424 8576 15430 8628
rect 16565 8619 16623 8625
rect 16565 8585 16577 8619
rect 16611 8616 16623 8619
rect 17390 8616 17396 8628
rect 16611 8588 17396 8616
rect 16611 8585 16623 8588
rect 16565 8579 16623 8585
rect 17390 8576 17396 8588
rect 17448 8576 17454 8628
rect 18494 8616 18500 8628
rect 18455 8588 18500 8616
rect 18494 8576 18500 8588
rect 18552 8576 18558 8628
rect 19782 8576 19788 8628
rect 19840 8616 19846 8628
rect 19969 8619 20027 8625
rect 19969 8616 19981 8619
rect 19840 8588 19981 8616
rect 19840 8576 19846 8588
rect 19969 8585 19981 8588
rect 20015 8585 20027 8619
rect 20610 8616 20616 8628
rect 20571 8588 20616 8616
rect 19969 8579 20027 8585
rect 20610 8576 20616 8588
rect 20668 8576 20674 8628
rect 21530 8576 21536 8628
rect 21588 8616 21594 8628
rect 21625 8619 21683 8625
rect 21625 8616 21637 8619
rect 21588 8588 21637 8616
rect 21588 8576 21594 8588
rect 21625 8585 21637 8588
rect 21671 8616 21683 8619
rect 24753 8619 24811 8625
rect 24753 8616 24765 8619
rect 21671 8588 22404 8616
rect 21671 8585 21683 8588
rect 21625 8579 21683 8585
rect 20334 8508 20340 8560
rect 20392 8548 20398 8560
rect 21717 8551 21775 8557
rect 21717 8548 21729 8551
rect 20392 8520 21729 8548
rect 20392 8508 20398 8520
rect 21717 8517 21729 8520
rect 21763 8517 21775 8551
rect 21717 8511 21775 8517
rect 14078 8480 14084 8492
rect 14039 8452 14084 8480
rect 14078 8440 14084 8452
rect 14136 8440 14142 8492
rect 15090 8440 15096 8492
rect 15148 8480 15154 8492
rect 15185 8483 15243 8489
rect 15185 8480 15197 8483
rect 15148 8452 15197 8480
rect 15148 8440 15154 8452
rect 15185 8449 15197 8452
rect 15231 8449 15243 8483
rect 18586 8480 18592 8492
rect 18547 8452 18592 8480
rect 15185 8443 15243 8449
rect 18586 8440 18592 8452
rect 18644 8440 18650 8492
rect 22174 8480 22180 8492
rect 22135 8452 22180 8480
rect 22174 8440 22180 8452
rect 22232 8440 22238 8492
rect 22376 8489 22404 8588
rect 22928 8588 24765 8616
rect 22361 8483 22419 8489
rect 22361 8449 22373 8483
rect 22407 8480 22419 8483
rect 22928 8480 22956 8588
rect 24753 8585 24765 8588
rect 24799 8585 24811 8619
rect 24753 8579 24811 8585
rect 23186 8548 23192 8560
rect 23147 8520 23192 8548
rect 23186 8508 23192 8520
rect 23244 8508 23250 8560
rect 22407 8452 22956 8480
rect 22407 8449 22419 8452
rect 22361 8443 22419 8449
rect 9021 8415 9079 8421
rect 9021 8381 9033 8415
rect 9067 8412 9079 8415
rect 9481 8415 9539 8421
rect 9481 8412 9493 8415
rect 9067 8384 9493 8412
rect 9067 8381 9079 8384
rect 9021 8375 9079 8381
rect 9481 8381 9493 8384
rect 9527 8412 9539 8415
rect 10674 8412 10680 8424
rect 9527 8384 10680 8412
rect 9527 8381 9539 8384
rect 9481 8375 9539 8381
rect 10674 8372 10680 8384
rect 10732 8372 10738 8424
rect 13069 8415 13127 8421
rect 13069 8381 13081 8415
rect 13115 8412 13127 8415
rect 13989 8415 14047 8421
rect 13989 8412 14001 8415
rect 13115 8384 14001 8412
rect 13115 8381 13127 8384
rect 13069 8375 13127 8381
rect 13989 8381 14001 8384
rect 14035 8412 14047 8415
rect 14262 8412 14268 8424
rect 14035 8384 14268 8412
rect 14035 8381 14047 8384
rect 13989 8375 14047 8381
rect 14262 8372 14268 8384
rect 14320 8372 14326 8424
rect 18494 8372 18500 8424
rect 18552 8412 18558 8424
rect 18845 8415 18903 8421
rect 18845 8412 18857 8415
rect 18552 8384 18857 8412
rect 18552 8372 18558 8384
rect 18845 8381 18857 8384
rect 18891 8381 18903 8415
rect 18845 8375 18903 8381
rect 21898 8372 21904 8424
rect 21956 8412 21962 8424
rect 22085 8415 22143 8421
rect 22085 8412 22097 8415
rect 21956 8384 22097 8412
rect 21956 8372 21962 8384
rect 22085 8381 22097 8384
rect 22131 8381 22143 8415
rect 22192 8412 22220 8440
rect 23186 8412 23192 8424
rect 22192 8384 23192 8412
rect 22085 8375 22143 8381
rect 23186 8372 23192 8384
rect 23244 8372 23250 8424
rect 23370 8412 23376 8424
rect 23283 8384 23376 8412
rect 23370 8372 23376 8384
rect 23428 8412 23434 8424
rect 24658 8412 24664 8424
rect 23428 8384 24664 8412
rect 23428 8372 23434 8384
rect 24658 8372 24664 8384
rect 24716 8372 24722 8424
rect 9389 8347 9447 8353
rect 9389 8313 9401 8347
rect 9435 8344 9447 8347
rect 9570 8344 9576 8356
rect 9435 8316 9576 8344
rect 9435 8313 9447 8316
rect 9389 8307 9447 8313
rect 9570 8304 9576 8316
rect 9628 8344 9634 8356
rect 9726 8347 9784 8353
rect 9726 8344 9738 8347
rect 9628 8316 9738 8344
rect 9628 8304 9634 8316
rect 9726 8313 9738 8316
rect 9772 8313 9784 8347
rect 13342 8344 13348 8356
rect 13303 8316 13348 8344
rect 9726 8307 9784 8313
rect 13342 8304 13348 8316
rect 13400 8344 13406 8356
rect 13897 8347 13955 8353
rect 13897 8344 13909 8347
rect 13400 8316 13909 8344
rect 13400 8304 13406 8316
rect 13897 8313 13909 8316
rect 13943 8313 13955 8347
rect 13897 8307 13955 8313
rect 14725 8347 14783 8353
rect 14725 8313 14737 8347
rect 14771 8344 14783 8347
rect 14814 8344 14820 8356
rect 14771 8316 14820 8344
rect 14771 8313 14783 8316
rect 14725 8307 14783 8313
rect 14814 8304 14820 8316
rect 14872 8344 14878 8356
rect 15452 8347 15510 8353
rect 15452 8344 15464 8347
rect 14872 8316 15464 8344
rect 14872 8304 14878 8316
rect 15452 8313 15464 8316
rect 15498 8344 15510 8347
rect 15550 8344 15556 8356
rect 15498 8316 15556 8344
rect 15498 8313 15510 8316
rect 15452 8307 15510 8313
rect 15550 8304 15556 8316
rect 15608 8344 15614 8356
rect 15608 8316 16240 8344
rect 15608 8304 15614 8316
rect 10861 8279 10919 8285
rect 10861 8245 10873 8279
rect 10907 8276 10919 8279
rect 10950 8276 10956 8288
rect 10907 8248 10956 8276
rect 10907 8245 10919 8248
rect 10861 8239 10919 8245
rect 10950 8236 10956 8248
rect 11008 8236 11014 8288
rect 12149 8279 12207 8285
rect 12149 8245 12161 8279
rect 12195 8276 12207 8279
rect 12514 8276 12520 8288
rect 12195 8248 12520 8276
rect 12195 8245 12207 8248
rect 12149 8239 12207 8245
rect 12514 8236 12520 8248
rect 12572 8236 12578 8288
rect 16212 8276 16240 8316
rect 16746 8304 16752 8356
rect 16804 8344 16810 8356
rect 17945 8347 18003 8353
rect 17945 8344 17957 8347
rect 16804 8316 17957 8344
rect 16804 8304 16810 8316
rect 17945 8313 17957 8316
rect 17991 8313 18003 8347
rect 20978 8344 20984 8356
rect 20939 8316 20984 8344
rect 17945 8307 18003 8313
rect 20978 8304 20984 8316
rect 21036 8304 21042 8356
rect 22450 8304 22456 8356
rect 22508 8344 22514 8356
rect 22821 8347 22879 8353
rect 22821 8344 22833 8347
rect 22508 8316 22833 8344
rect 22508 8304 22514 8316
rect 22821 8313 22833 8316
rect 22867 8344 22879 8347
rect 23640 8347 23698 8353
rect 23640 8344 23652 8347
rect 22867 8316 23652 8344
rect 22867 8313 22879 8316
rect 22821 8307 22879 8313
rect 23640 8313 23652 8316
rect 23686 8344 23698 8347
rect 23738 8344 23744 8356
rect 23686 8316 23744 8344
rect 23686 8313 23698 8316
rect 23640 8307 23698 8313
rect 23738 8304 23744 8316
rect 23796 8304 23802 8356
rect 16378 8276 16384 8288
rect 16212 8248 16384 8276
rect 16378 8236 16384 8248
rect 16436 8236 16442 8288
rect 816 8186 26576 8208
rect 816 8134 10027 8186
rect 10079 8134 10091 8186
rect 10143 8134 10155 8186
rect 10207 8134 10219 8186
rect 10271 8134 19360 8186
rect 19412 8134 19424 8186
rect 19476 8134 19488 8186
rect 19540 8134 19552 8186
rect 19604 8134 26576 8186
rect 816 8112 26576 8134
rect 11778 8032 11784 8084
rect 11836 8072 11842 8084
rect 12057 8075 12115 8081
rect 12057 8072 12069 8075
rect 11836 8044 12069 8072
rect 11836 8032 11842 8044
rect 12057 8041 12069 8044
rect 12103 8041 12115 8075
rect 13158 8072 13164 8084
rect 13119 8044 13164 8072
rect 12057 8035 12115 8041
rect 13158 8032 13164 8044
rect 13216 8032 13222 8084
rect 14814 8072 14820 8084
rect 14775 8044 14820 8072
rect 14814 8032 14820 8044
rect 14872 8032 14878 8084
rect 16378 8072 16384 8084
rect 16339 8044 16384 8072
rect 16378 8032 16384 8044
rect 16436 8032 16442 8084
rect 17758 8032 17764 8084
rect 17816 8072 17822 8084
rect 17853 8075 17911 8081
rect 17853 8072 17865 8075
rect 17816 8044 17865 8072
rect 17816 8032 17822 8044
rect 17853 8041 17865 8044
rect 17899 8041 17911 8075
rect 17853 8035 17911 8041
rect 20061 8075 20119 8081
rect 20061 8041 20073 8075
rect 20107 8072 20119 8075
rect 20334 8072 20340 8084
rect 20107 8044 20340 8072
rect 20107 8041 20119 8044
rect 20061 8035 20119 8041
rect 10950 7945 10956 7948
rect 10585 7939 10643 7945
rect 10585 7905 10597 7939
rect 10631 7936 10643 7939
rect 10944 7936 10956 7945
rect 10631 7908 10956 7936
rect 10631 7905 10643 7908
rect 10585 7899 10643 7905
rect 10944 7899 10956 7908
rect 10950 7896 10956 7899
rect 11008 7896 11014 7948
rect 12514 7896 12520 7948
rect 12572 7936 12578 7948
rect 13529 7939 13587 7945
rect 13529 7936 13541 7939
rect 12572 7908 13541 7936
rect 12572 7896 12578 7908
rect 13529 7905 13541 7908
rect 13575 7905 13587 7939
rect 13529 7899 13587 7905
rect 14538 7896 14544 7948
rect 14596 7936 14602 7948
rect 15257 7939 15315 7945
rect 15257 7936 15269 7939
rect 14596 7908 15269 7936
rect 14596 7896 14602 7908
rect 15257 7905 15269 7908
rect 15303 7905 15315 7939
rect 15257 7899 15315 7905
rect 17393 7939 17451 7945
rect 17393 7905 17405 7939
rect 17439 7936 17451 7939
rect 17850 7936 17856 7948
rect 17439 7908 17856 7936
rect 17439 7905 17451 7908
rect 17393 7899 17451 7905
rect 17850 7896 17856 7908
rect 17908 7936 17914 7948
rect 19233 7939 19291 7945
rect 17908 7908 18080 7936
rect 17908 7896 17914 7908
rect 9389 7871 9447 7877
rect 9389 7837 9401 7871
rect 9435 7868 9447 7871
rect 9754 7868 9760 7880
rect 9435 7840 9760 7868
rect 9435 7837 9447 7840
rect 9389 7831 9447 7837
rect 9754 7828 9760 7840
rect 9812 7828 9818 7880
rect 10674 7868 10680 7880
rect 10635 7840 10680 7868
rect 10674 7828 10680 7840
rect 10732 7828 10738 7880
rect 13618 7868 13624 7880
rect 13579 7840 13624 7868
rect 13618 7828 13624 7840
rect 13676 7828 13682 7880
rect 13713 7871 13771 7877
rect 13713 7837 13725 7871
rect 13759 7837 13771 7871
rect 13713 7831 13771 7837
rect 14449 7871 14507 7877
rect 14449 7837 14461 7871
rect 14495 7868 14507 7871
rect 14998 7868 15004 7880
rect 14495 7840 15004 7868
rect 14495 7837 14507 7840
rect 14449 7831 14507 7837
rect 12793 7803 12851 7809
rect 12793 7769 12805 7803
rect 12839 7800 12851 7803
rect 12974 7800 12980 7812
rect 12839 7772 12980 7800
rect 12839 7769 12851 7772
rect 12793 7763 12851 7769
rect 12974 7760 12980 7772
rect 13032 7800 13038 7812
rect 13728 7800 13756 7831
rect 14998 7828 15004 7840
rect 15056 7828 15062 7880
rect 18052 7877 18080 7908
rect 19233 7905 19245 7939
rect 19279 7936 19291 7939
rect 20076 7936 20104 8035
rect 20334 8032 20340 8044
rect 20392 8032 20398 8084
rect 23186 8072 23192 8084
rect 23147 8044 23192 8072
rect 23186 8032 23192 8044
rect 23244 8032 23250 8084
rect 23646 8072 23652 8084
rect 23607 8044 23652 8072
rect 23646 8032 23652 8044
rect 23704 8032 23710 8084
rect 24658 8072 24664 8084
rect 24619 8044 24664 8072
rect 24658 8032 24664 8044
rect 24716 8032 24722 8084
rect 20426 7964 20432 8016
rect 20484 8004 20490 8016
rect 21622 8004 21628 8016
rect 20484 7976 21628 8004
rect 20484 7964 20490 7976
rect 20628 7945 20656 7976
rect 21622 7964 21628 7976
rect 21680 7964 21686 8016
rect 19279 7908 20104 7936
rect 20613 7939 20671 7945
rect 19279 7905 19291 7908
rect 19233 7899 19291 7905
rect 20613 7905 20625 7939
rect 20659 7905 20671 7939
rect 20613 7899 20671 7905
rect 20880 7939 20938 7945
rect 20880 7905 20892 7939
rect 20926 7936 20938 7939
rect 21346 7936 21352 7948
rect 20926 7908 21352 7936
rect 20926 7905 20938 7908
rect 20880 7899 20938 7905
rect 21346 7896 21352 7908
rect 21404 7896 21410 7948
rect 23094 7896 23100 7948
rect 23152 7936 23158 7948
rect 23557 7939 23615 7945
rect 23557 7936 23569 7939
rect 23152 7908 23569 7936
rect 23152 7896 23158 7908
rect 23557 7905 23569 7908
rect 23603 7905 23615 7939
rect 23557 7899 23615 7905
rect 24566 7896 24572 7948
rect 24624 7936 24630 7948
rect 24753 7939 24811 7945
rect 24753 7936 24765 7939
rect 24624 7908 24765 7936
rect 24624 7896 24630 7908
rect 24753 7905 24765 7908
rect 24799 7905 24811 7939
rect 24753 7899 24811 7905
rect 17945 7871 18003 7877
rect 17945 7868 17957 7871
rect 17224 7840 17957 7868
rect 13032 7772 13756 7800
rect 13032 7760 13038 7772
rect 17224 7744 17252 7840
rect 17945 7837 17957 7840
rect 17991 7837 18003 7871
rect 17945 7831 18003 7837
rect 18037 7871 18095 7877
rect 18037 7837 18049 7871
rect 18083 7837 18095 7871
rect 18037 7831 18095 7837
rect 18310 7828 18316 7880
rect 18368 7868 18374 7880
rect 18586 7868 18592 7880
rect 18368 7840 18592 7868
rect 18368 7828 18374 7840
rect 18586 7828 18592 7840
rect 18644 7828 18650 7880
rect 19509 7871 19567 7877
rect 19509 7837 19521 7871
rect 19555 7868 19567 7871
rect 19874 7868 19880 7880
rect 19555 7840 19880 7868
rect 19555 7837 19567 7840
rect 19509 7831 19567 7837
rect 19874 7828 19880 7840
rect 19932 7828 19938 7880
rect 23738 7828 23744 7880
rect 23796 7868 23802 7880
rect 23796 7840 23841 7868
rect 23796 7828 23802 7840
rect 23922 7828 23928 7880
rect 23980 7868 23986 7880
rect 24658 7868 24664 7880
rect 23980 7840 24664 7868
rect 23980 7828 23986 7840
rect 24658 7828 24664 7840
rect 24716 7828 24722 7880
rect 17485 7803 17543 7809
rect 17485 7769 17497 7803
rect 17531 7800 17543 7803
rect 18865 7803 18923 7809
rect 18865 7800 18877 7803
rect 17531 7772 18877 7800
rect 17531 7769 17543 7772
rect 17485 7763 17543 7769
rect 18865 7769 18877 7772
rect 18911 7800 18923 7803
rect 19230 7800 19236 7812
rect 18911 7772 19236 7800
rect 18911 7769 18923 7772
rect 18865 7763 18923 7769
rect 19230 7760 19236 7772
rect 19288 7760 19294 7812
rect 23940 7800 23968 7828
rect 24934 7800 24940 7812
rect 21548 7772 23968 7800
rect 24895 7772 24940 7800
rect 7822 7732 7828 7744
rect 7783 7704 7828 7732
rect 7822 7692 7828 7704
rect 7880 7692 7886 7744
rect 17025 7735 17083 7741
rect 17025 7701 17037 7735
rect 17071 7732 17083 7735
rect 17206 7732 17212 7744
rect 17071 7704 17212 7732
rect 17071 7701 17083 7704
rect 17025 7695 17083 7701
rect 17206 7692 17212 7704
rect 17264 7692 17270 7744
rect 18310 7692 18316 7744
rect 18368 7732 18374 7744
rect 18497 7735 18555 7741
rect 18497 7732 18509 7735
rect 18368 7704 18509 7732
rect 18368 7692 18374 7704
rect 18497 7701 18509 7704
rect 18543 7701 18555 7735
rect 18497 7695 18555 7701
rect 20429 7735 20487 7741
rect 20429 7701 20441 7735
rect 20475 7732 20487 7735
rect 20794 7732 20800 7744
rect 20475 7704 20800 7732
rect 20475 7701 20487 7704
rect 20429 7695 20487 7701
rect 20794 7692 20800 7704
rect 20852 7692 20858 7744
rect 20886 7692 20892 7744
rect 20944 7732 20950 7744
rect 21548 7732 21576 7772
rect 24934 7760 24940 7772
rect 24992 7760 24998 7812
rect 21990 7732 21996 7744
rect 20944 7704 21576 7732
rect 21951 7704 21996 7732
rect 20944 7692 20950 7704
rect 21990 7692 21996 7704
rect 22048 7692 22054 7744
rect 22174 7692 22180 7744
rect 22232 7732 22238 7744
rect 22545 7735 22603 7741
rect 22545 7732 22557 7735
rect 22232 7704 22557 7732
rect 22232 7692 22238 7704
rect 22545 7701 22557 7704
rect 22591 7701 22603 7735
rect 22910 7732 22916 7744
rect 22871 7704 22916 7732
rect 22545 7695 22603 7701
rect 22910 7692 22916 7704
rect 22968 7692 22974 7744
rect 23922 7692 23928 7744
rect 23980 7732 23986 7744
rect 24201 7735 24259 7741
rect 24201 7732 24213 7735
rect 23980 7704 24213 7732
rect 23980 7692 23986 7704
rect 24201 7701 24213 7704
rect 24247 7701 24259 7735
rect 24201 7695 24259 7701
rect 816 7642 26576 7664
rect 816 7590 5360 7642
rect 5412 7590 5424 7642
rect 5476 7590 5488 7642
rect 5540 7590 5552 7642
rect 5604 7590 14694 7642
rect 14746 7590 14758 7642
rect 14810 7590 14822 7642
rect 14874 7590 14886 7642
rect 14938 7590 24027 7642
rect 24079 7590 24091 7642
rect 24143 7590 24155 7642
rect 24207 7590 24219 7642
rect 24271 7590 26576 7642
rect 816 7568 26576 7590
rect 3866 7488 3872 7540
rect 3924 7528 3930 7540
rect 5154 7528 5160 7540
rect 3924 7500 5160 7528
rect 3924 7488 3930 7500
rect 5154 7488 5160 7500
rect 5212 7488 5218 7540
rect 7733 7531 7791 7537
rect 7733 7497 7745 7531
rect 7779 7528 7791 7531
rect 8006 7528 8012 7540
rect 7779 7500 8012 7528
rect 7779 7497 7791 7500
rect 7733 7491 7791 7497
rect 8006 7488 8012 7500
rect 8064 7488 8070 7540
rect 10490 7528 10496 7540
rect 10451 7500 10496 7528
rect 10490 7488 10496 7500
rect 10548 7488 10554 7540
rect 12514 7528 12520 7540
rect 12475 7500 12520 7528
rect 12514 7488 12520 7500
rect 12572 7488 12578 7540
rect 15093 7531 15151 7537
rect 15093 7497 15105 7531
rect 15139 7528 15151 7531
rect 15182 7528 15188 7540
rect 15139 7500 15188 7528
rect 15139 7497 15151 7500
rect 15093 7491 15151 7497
rect 15182 7488 15188 7500
rect 15240 7488 15246 7540
rect 20794 7528 20800 7540
rect 20755 7500 20800 7528
rect 20794 7488 20800 7500
rect 20852 7488 20858 7540
rect 20889 7531 20947 7537
rect 20889 7497 20901 7531
rect 20935 7528 20947 7531
rect 21254 7528 21260 7540
rect 20935 7500 21260 7528
rect 20935 7497 20947 7500
rect 20889 7491 20947 7497
rect 21254 7488 21260 7500
rect 21312 7488 21318 7540
rect 21346 7488 21352 7540
rect 21404 7528 21410 7540
rect 21901 7531 21959 7537
rect 21901 7528 21913 7531
rect 21404 7500 21913 7528
rect 21404 7488 21410 7500
rect 21901 7497 21913 7500
rect 21947 7497 21959 7531
rect 22450 7528 22456 7540
rect 22411 7500 22456 7528
rect 21901 7491 21959 7497
rect 22450 7488 22456 7500
rect 22508 7488 22514 7540
rect 22821 7531 22879 7537
rect 22821 7497 22833 7531
rect 22867 7528 22879 7531
rect 23646 7528 23652 7540
rect 22867 7500 23652 7528
rect 22867 7497 22879 7500
rect 22821 7491 22879 7497
rect 23646 7488 23652 7500
rect 23704 7488 23710 7540
rect 24566 7488 24572 7540
rect 24624 7528 24630 7540
rect 24753 7531 24811 7537
rect 24753 7528 24765 7531
rect 24624 7500 24765 7528
rect 24624 7488 24630 7500
rect 24753 7497 24765 7500
rect 24799 7497 24811 7531
rect 25670 7528 25676 7540
rect 25631 7500 25676 7528
rect 24753 7491 24811 7497
rect 25670 7488 25676 7500
rect 25728 7488 25734 7540
rect 25946 7488 25952 7540
rect 26004 7528 26010 7540
rect 26590 7528 26596 7540
rect 26004 7500 26596 7528
rect 26004 7488 26010 7500
rect 26590 7488 26596 7500
rect 26648 7488 26654 7540
rect 9202 7460 9208 7472
rect 9163 7432 9208 7460
rect 9202 7420 9208 7432
rect 9260 7420 9266 7472
rect 14354 7420 14360 7472
rect 14412 7460 14418 7472
rect 16473 7463 16531 7469
rect 16473 7460 16485 7463
rect 14412 7432 16485 7460
rect 14412 7420 14418 7432
rect 16473 7429 16485 7432
rect 16519 7460 16531 7463
rect 16746 7460 16752 7472
rect 16519 7432 16752 7460
rect 16519 7429 16531 7432
rect 16473 7423 16531 7429
rect 16746 7420 16752 7432
rect 16804 7420 16810 7472
rect 19138 7420 19144 7472
rect 19196 7460 19202 7472
rect 19325 7463 19383 7469
rect 19325 7460 19337 7463
rect 19196 7432 19337 7460
rect 19196 7420 19202 7432
rect 19325 7429 19337 7432
rect 19371 7429 19383 7463
rect 19325 7423 19383 7429
rect 10950 7352 10956 7404
rect 11008 7392 11014 7404
rect 11137 7395 11195 7401
rect 11137 7392 11149 7395
rect 11008 7364 11149 7392
rect 11008 7352 11014 7364
rect 11137 7361 11149 7364
rect 11183 7392 11195 7395
rect 11505 7395 11563 7401
rect 11505 7392 11517 7395
rect 11183 7364 11517 7392
rect 11183 7361 11195 7364
rect 11137 7355 11195 7361
rect 11505 7361 11517 7364
rect 11551 7361 11563 7395
rect 11505 7355 11563 7361
rect 11965 7395 12023 7401
rect 11965 7361 11977 7395
rect 12011 7392 12023 7395
rect 12054 7392 12060 7404
rect 12011 7364 12060 7392
rect 12011 7361 12023 7364
rect 11965 7355 12023 7361
rect 12054 7352 12060 7364
rect 12112 7392 12118 7404
rect 12701 7395 12759 7401
rect 12701 7392 12713 7395
rect 12112 7364 12713 7392
rect 12112 7352 12118 7364
rect 12701 7361 12713 7364
rect 12747 7361 12759 7395
rect 18310 7392 18316 7404
rect 18271 7364 18316 7392
rect 12701 7355 12759 7361
rect 18310 7352 18316 7364
rect 18368 7352 18374 7404
rect 19966 7392 19972 7404
rect 19927 7364 19972 7392
rect 19966 7352 19972 7364
rect 20024 7392 20030 7404
rect 20150 7392 20156 7404
rect 20024 7364 20156 7392
rect 20024 7352 20030 7364
rect 20150 7352 20156 7364
rect 20208 7352 20214 7404
rect 20812 7392 20840 7488
rect 23094 7460 23100 7472
rect 23055 7432 23100 7460
rect 23094 7420 23100 7432
rect 23152 7420 23158 7472
rect 21438 7392 21444 7404
rect 20812 7364 21444 7392
rect 21438 7352 21444 7364
rect 21496 7352 21502 7404
rect 24014 7392 24020 7404
rect 23975 7364 24020 7392
rect 24014 7352 24020 7364
rect 24072 7352 24078 7404
rect 7822 7324 7828 7336
rect 7783 7296 7828 7324
rect 7822 7284 7828 7296
rect 7880 7284 7886 7336
rect 12974 7333 12980 7336
rect 12968 7324 12980 7333
rect 12935 7296 12980 7324
rect 12968 7287 12980 7296
rect 12974 7284 12980 7287
rect 13032 7284 13038 7336
rect 15182 7324 15188 7336
rect 15143 7296 15188 7324
rect 15182 7284 15188 7296
rect 15240 7284 15246 7336
rect 19785 7327 19843 7333
rect 19785 7293 19797 7327
rect 19831 7324 19843 7327
rect 20058 7324 20064 7336
rect 19831 7296 20064 7324
rect 19831 7293 19843 7296
rect 19785 7287 19843 7293
rect 20058 7284 20064 7296
rect 20116 7324 20122 7336
rect 20429 7327 20487 7333
rect 20429 7324 20441 7327
rect 20116 7296 20441 7324
rect 20116 7284 20122 7296
rect 20429 7293 20441 7296
rect 20475 7324 20487 7327
rect 20886 7324 20892 7336
rect 20475 7296 20892 7324
rect 20475 7293 20487 7296
rect 20429 7287 20487 7293
rect 20886 7284 20892 7296
rect 20944 7284 20950 7336
rect 22910 7324 22916 7336
rect 21272 7296 22916 7324
rect 8006 7216 8012 7268
rect 8064 7265 8070 7268
rect 8064 7259 8128 7265
rect 8064 7225 8082 7259
rect 8116 7225 8128 7259
rect 10306 7256 10312 7268
rect 10267 7228 10312 7256
rect 8064 7219 8128 7225
rect 8064 7216 8070 7219
rect 10306 7216 10312 7228
rect 10364 7256 10370 7268
rect 10861 7259 10919 7265
rect 10861 7256 10873 7259
rect 10364 7228 10873 7256
rect 10364 7216 10370 7228
rect 10861 7225 10873 7228
rect 10907 7225 10919 7259
rect 18221 7259 18279 7265
rect 18221 7256 18233 7259
rect 10861 7219 10919 7225
rect 17500 7228 18233 7256
rect 9202 7148 9208 7200
rect 9260 7188 9266 7200
rect 10033 7191 10091 7197
rect 10033 7188 10045 7191
rect 9260 7160 10045 7188
rect 9260 7148 9266 7160
rect 10033 7157 10045 7160
rect 10079 7188 10091 7191
rect 10674 7188 10680 7200
rect 10079 7160 10680 7188
rect 10079 7157 10091 7160
rect 10033 7151 10091 7157
rect 10674 7148 10680 7160
rect 10732 7148 10738 7200
rect 10766 7148 10772 7200
rect 10824 7188 10830 7200
rect 10953 7191 11011 7197
rect 10953 7188 10965 7191
rect 10824 7160 10965 7188
rect 10824 7148 10830 7160
rect 10953 7157 10965 7160
rect 10999 7157 11011 7191
rect 10953 7151 11011 7157
rect 14081 7191 14139 7197
rect 14081 7157 14093 7191
rect 14127 7188 14139 7191
rect 14538 7188 14544 7200
rect 14127 7160 14544 7188
rect 14127 7157 14139 7160
rect 14081 7151 14139 7157
rect 14538 7148 14544 7160
rect 14596 7188 14602 7200
rect 14633 7191 14691 7197
rect 14633 7188 14645 7191
rect 14596 7160 14645 7188
rect 14596 7148 14602 7160
rect 14633 7157 14645 7160
rect 14679 7157 14691 7191
rect 14633 7151 14691 7157
rect 17114 7148 17120 7200
rect 17172 7188 17178 7200
rect 17500 7197 17528 7228
rect 18221 7225 18233 7228
rect 18267 7225 18279 7259
rect 18221 7219 18279 7225
rect 19233 7259 19291 7265
rect 19233 7225 19245 7259
rect 19279 7256 19291 7259
rect 19693 7259 19751 7265
rect 19693 7256 19705 7259
rect 19279 7228 19705 7256
rect 19279 7225 19291 7228
rect 19233 7219 19291 7225
rect 19693 7225 19705 7228
rect 19739 7256 19751 7259
rect 19966 7256 19972 7268
rect 19739 7228 19972 7256
rect 19739 7225 19751 7228
rect 19693 7219 19751 7225
rect 19966 7216 19972 7228
rect 20024 7216 20030 7268
rect 21272 7200 21300 7296
rect 22910 7284 22916 7296
rect 22968 7284 22974 7336
rect 25029 7327 25087 7333
rect 25029 7293 25041 7327
rect 25075 7324 25087 7327
rect 25670 7324 25676 7336
rect 25075 7296 25676 7324
rect 25075 7293 25087 7296
rect 25029 7287 25087 7293
rect 25670 7284 25676 7296
rect 25728 7284 25734 7336
rect 17485 7191 17543 7197
rect 17485 7188 17497 7191
rect 17172 7160 17497 7188
rect 17172 7148 17178 7160
rect 17485 7157 17497 7160
rect 17531 7157 17543 7191
rect 17485 7151 17543 7157
rect 17666 7148 17672 7200
rect 17724 7188 17730 7200
rect 17761 7191 17819 7197
rect 17761 7188 17773 7191
rect 17724 7160 17773 7188
rect 17724 7148 17730 7160
rect 17761 7157 17773 7160
rect 17807 7157 17819 7191
rect 18126 7188 18132 7200
rect 18039 7160 18132 7188
rect 17761 7151 17819 7157
rect 18126 7148 18132 7160
rect 18184 7188 18190 7200
rect 18862 7188 18868 7200
rect 18184 7160 18868 7188
rect 18184 7148 18190 7160
rect 18862 7148 18868 7160
rect 18920 7148 18926 7200
rect 21254 7188 21260 7200
rect 21215 7160 21260 7188
rect 21254 7148 21260 7160
rect 21312 7148 21318 7200
rect 21349 7191 21407 7197
rect 21349 7157 21361 7191
rect 21395 7188 21407 7191
rect 21530 7188 21536 7200
rect 21395 7160 21536 7188
rect 21395 7157 21407 7160
rect 21349 7151 21407 7157
rect 21530 7148 21536 7160
rect 21588 7188 21594 7200
rect 22174 7188 22180 7200
rect 21588 7160 22180 7188
rect 21588 7148 21594 7160
rect 22174 7148 22180 7160
rect 22232 7148 22238 7200
rect 23462 7188 23468 7200
rect 23423 7160 23468 7188
rect 23462 7148 23468 7160
rect 23520 7148 23526 7200
rect 23830 7188 23836 7200
rect 23791 7160 23836 7188
rect 23830 7148 23836 7160
rect 23888 7148 23894 7200
rect 23922 7148 23928 7200
rect 23980 7188 23986 7200
rect 25210 7188 25216 7200
rect 23980 7160 24025 7188
rect 25171 7160 25216 7188
rect 23980 7148 23986 7160
rect 25210 7148 25216 7160
rect 25268 7148 25274 7200
rect 816 7098 26576 7120
rect 816 7046 10027 7098
rect 10079 7046 10091 7098
rect 10143 7046 10155 7098
rect 10207 7046 10219 7098
rect 10271 7046 19360 7098
rect 19412 7046 19424 7098
rect 19476 7046 19488 7098
rect 19540 7046 19552 7098
rect 19604 7046 26576 7098
rect 816 7024 26576 7046
rect 9754 6984 9760 6996
rect 9715 6956 9760 6984
rect 9754 6944 9760 6956
rect 9812 6944 9818 6996
rect 11137 6987 11195 6993
rect 11137 6953 11149 6987
rect 11183 6984 11195 6987
rect 12793 6987 12851 6993
rect 11183 6956 11217 6984
rect 11183 6953 11195 6956
rect 11137 6947 11195 6953
rect 12793 6953 12805 6987
rect 12839 6984 12851 6987
rect 12974 6984 12980 6996
rect 12839 6956 12980 6984
rect 12839 6953 12851 6956
rect 12793 6947 12851 6953
rect 7822 6916 7828 6928
rect 6828 6888 7828 6916
rect 6828 6857 6856 6888
rect 7822 6876 7828 6888
rect 7880 6876 7886 6928
rect 10674 6876 10680 6928
rect 10732 6916 10738 6928
rect 11045 6919 11103 6925
rect 11045 6916 11057 6919
rect 10732 6888 11057 6916
rect 10732 6876 10738 6888
rect 11045 6885 11057 6888
rect 11091 6916 11103 6919
rect 11152 6916 11180 6947
rect 12974 6944 12980 6956
rect 13032 6984 13038 6996
rect 13345 6987 13403 6993
rect 13345 6984 13357 6987
rect 13032 6956 13357 6984
rect 13032 6944 13038 6956
rect 13345 6953 13357 6956
rect 13391 6953 13403 6987
rect 13345 6947 13403 6953
rect 14262 6944 14268 6996
rect 14320 6984 14326 6996
rect 15550 6984 15556 6996
rect 14320 6956 15556 6984
rect 14320 6944 14326 6956
rect 15550 6944 15556 6956
rect 15608 6984 15614 6996
rect 16013 6987 16071 6993
rect 16013 6984 16025 6987
rect 15608 6956 16025 6984
rect 15608 6944 15614 6956
rect 16013 6953 16025 6956
rect 16059 6953 16071 6987
rect 16013 6947 16071 6953
rect 17758 6944 17764 6996
rect 17816 6984 17822 6996
rect 18313 6987 18371 6993
rect 18313 6984 18325 6987
rect 17816 6956 18325 6984
rect 17816 6944 17822 6956
rect 18313 6953 18325 6956
rect 18359 6953 18371 6987
rect 19230 6984 19236 6996
rect 19191 6956 19236 6984
rect 18313 6947 18371 6953
rect 19230 6944 19236 6956
rect 19288 6944 19294 6996
rect 19969 6987 20027 6993
rect 19969 6953 19981 6987
rect 20015 6984 20027 6987
rect 20150 6984 20156 6996
rect 20015 6956 20156 6984
rect 20015 6953 20027 6956
rect 19969 6947 20027 6953
rect 20150 6944 20156 6956
rect 20208 6944 20214 6996
rect 20613 6987 20671 6993
rect 20613 6953 20625 6987
rect 20659 6984 20671 6987
rect 21254 6984 21260 6996
rect 20659 6956 21260 6984
rect 20659 6953 20671 6956
rect 20613 6947 20671 6953
rect 21254 6944 21260 6956
rect 21312 6944 21318 6996
rect 23830 6944 23836 6996
rect 23888 6984 23894 6996
rect 24569 6987 24627 6993
rect 24569 6984 24581 6987
rect 23888 6956 24581 6984
rect 23888 6944 23894 6956
rect 24569 6953 24581 6956
rect 24615 6953 24627 6987
rect 24569 6947 24627 6953
rect 12054 6916 12060 6928
rect 11091 6888 12060 6916
rect 11091 6885 11103 6888
rect 11045 6879 11103 6885
rect 11428 6860 11456 6888
rect 12054 6876 12060 6888
rect 12112 6876 12118 6928
rect 15921 6919 15979 6925
rect 15921 6885 15933 6919
rect 15967 6916 15979 6919
rect 16102 6916 16108 6928
rect 15967 6888 16108 6916
rect 15967 6885 15979 6888
rect 15921 6879 15979 6885
rect 16102 6876 16108 6888
rect 16160 6876 16166 6928
rect 18862 6876 18868 6928
rect 18920 6916 18926 6928
rect 21806 6916 21812 6928
rect 18920 6888 21812 6916
rect 18920 6876 18926 6888
rect 21806 6876 21812 6888
rect 21864 6876 21870 6928
rect 6813 6851 6871 6857
rect 6813 6817 6825 6851
rect 6859 6817 6871 6851
rect 6813 6811 6871 6817
rect 6902 6808 6908 6860
rect 6960 6848 6966 6860
rect 7069 6851 7127 6857
rect 7069 6848 7081 6851
rect 6960 6820 7081 6848
rect 6960 6808 6966 6820
rect 7069 6817 7081 6820
rect 7115 6817 7127 6851
rect 7069 6811 7127 6817
rect 8190 6808 8196 6860
rect 8248 6848 8254 6860
rect 10493 6851 10551 6857
rect 10493 6848 10505 6851
rect 8248 6820 10505 6848
rect 8248 6808 8254 6820
rect 10493 6817 10505 6820
rect 10539 6848 10551 6851
rect 10766 6848 10772 6860
rect 10539 6820 10772 6848
rect 10539 6817 10551 6820
rect 10493 6811 10551 6817
rect 10766 6808 10772 6820
rect 10824 6808 10830 6860
rect 11318 6848 11324 6860
rect 11279 6820 11324 6848
rect 11318 6808 11324 6820
rect 11376 6808 11382 6860
rect 11410 6808 11416 6860
rect 11468 6848 11474 6860
rect 11686 6857 11692 6860
rect 11680 6848 11692 6857
rect 11468 6820 11561 6848
rect 11647 6820 11692 6848
rect 11468 6808 11474 6820
rect 11680 6811 11692 6820
rect 11686 6808 11692 6811
rect 11744 6808 11750 6860
rect 15185 6851 15243 6857
rect 15185 6817 15197 6851
rect 15231 6848 15243 6851
rect 15826 6848 15832 6860
rect 15231 6820 15832 6848
rect 15231 6817 15243 6820
rect 15185 6811 15243 6817
rect 15826 6808 15832 6820
rect 15884 6808 15890 6860
rect 16470 6808 16476 6860
rect 16528 6848 16534 6860
rect 16637 6851 16695 6857
rect 16637 6848 16649 6851
rect 16528 6820 16649 6848
rect 16528 6808 16534 6820
rect 16637 6817 16649 6820
rect 16683 6817 16695 6851
rect 20978 6848 20984 6860
rect 20939 6820 20984 6848
rect 16637 6811 16695 6817
rect 20978 6808 20984 6820
rect 21036 6808 21042 6860
rect 21898 6808 21904 6860
rect 21956 6848 21962 6860
rect 22542 6857 22548 6860
rect 22525 6851 22548 6857
rect 22525 6848 22537 6851
rect 21956 6820 22537 6848
rect 21956 6808 21962 6820
rect 22525 6817 22537 6820
rect 22600 6848 22606 6860
rect 22600 6820 22673 6848
rect 22525 6811 22548 6817
rect 22542 6808 22548 6811
rect 22600 6808 22606 6820
rect 24566 6808 24572 6860
rect 24624 6848 24630 6860
rect 24753 6851 24811 6857
rect 24753 6848 24765 6851
rect 24624 6820 24765 6848
rect 24624 6808 24630 6820
rect 24753 6817 24765 6820
rect 24799 6817 24811 6851
rect 24753 6811 24811 6817
rect 9662 6740 9668 6792
rect 9720 6780 9726 6792
rect 9849 6783 9907 6789
rect 9849 6780 9861 6783
rect 9720 6752 9861 6780
rect 9720 6740 9726 6752
rect 9849 6749 9861 6752
rect 9895 6749 9907 6783
rect 9849 6743 9907 6749
rect 9941 6783 9999 6789
rect 9941 6749 9953 6783
rect 9987 6749 9999 6783
rect 13894 6780 13900 6792
rect 13855 6752 13900 6780
rect 9941 6743 9999 6749
rect 9386 6712 9392 6724
rect 9347 6684 9392 6712
rect 9386 6672 9392 6684
rect 9444 6672 9450 6724
rect 9570 6672 9576 6724
rect 9628 6712 9634 6724
rect 9956 6712 9984 6743
rect 13894 6740 13900 6752
rect 13952 6740 13958 6792
rect 14538 6740 14544 6792
rect 14596 6780 14602 6792
rect 16105 6783 16163 6789
rect 14596 6752 15964 6780
rect 14596 6740 14602 6752
rect 15366 6712 15372 6724
rect 9628 6684 9984 6712
rect 15327 6684 15372 6712
rect 9628 6672 9634 6684
rect 15366 6672 15372 6684
rect 15424 6672 15430 6724
rect 15458 6672 15464 6724
rect 15516 6712 15522 6724
rect 15553 6715 15611 6721
rect 15553 6712 15565 6715
rect 15516 6684 15565 6712
rect 15516 6672 15522 6684
rect 15553 6681 15565 6684
rect 15599 6681 15611 6715
rect 15936 6712 15964 6752
rect 16105 6749 16117 6783
rect 16151 6749 16163 6783
rect 16105 6743 16163 6749
rect 16381 6783 16439 6789
rect 16381 6749 16393 6783
rect 16427 6749 16439 6783
rect 16381 6743 16439 6749
rect 16120 6712 16148 6743
rect 15936 6684 16148 6712
rect 15553 6675 15611 6681
rect 8193 6647 8251 6653
rect 8193 6613 8205 6647
rect 8239 6644 8251 6647
rect 9588 6644 9616 6672
rect 8239 6616 9616 6644
rect 8239 6613 8251 6616
rect 8193 6607 8251 6613
rect 13618 6604 13624 6656
rect 13676 6644 13682 6656
rect 13713 6647 13771 6653
rect 13713 6644 13725 6647
rect 13676 6616 13725 6644
rect 13676 6604 13682 6616
rect 13713 6613 13725 6616
rect 13759 6613 13771 6647
rect 13713 6607 13771 6613
rect 13802 6604 13808 6656
rect 13860 6644 13866 6656
rect 14357 6647 14415 6653
rect 14357 6644 14369 6647
rect 13860 6616 14369 6644
rect 13860 6604 13866 6616
rect 14357 6613 14369 6616
rect 14403 6613 14415 6647
rect 14357 6607 14415 6613
rect 14817 6647 14875 6653
rect 14817 6613 14829 6647
rect 14863 6644 14875 6647
rect 16396 6644 16424 6743
rect 18310 6740 18316 6792
rect 18368 6780 18374 6792
rect 18586 6780 18592 6792
rect 18368 6752 18592 6780
rect 18368 6740 18374 6752
rect 18586 6740 18592 6752
rect 18644 6740 18650 6792
rect 19325 6783 19383 6789
rect 19325 6749 19337 6783
rect 19371 6749 19383 6783
rect 19325 6743 19383 6749
rect 17761 6715 17819 6721
rect 17761 6681 17773 6715
rect 17807 6712 17819 6715
rect 17850 6712 17856 6724
rect 17807 6684 17856 6712
rect 17807 6681 17819 6684
rect 17761 6675 17819 6681
rect 17850 6672 17856 6684
rect 17908 6672 17914 6724
rect 18770 6672 18776 6724
rect 18828 6712 18834 6724
rect 18865 6715 18923 6721
rect 18865 6712 18877 6715
rect 18828 6684 18877 6712
rect 18828 6672 18834 6684
rect 18865 6681 18877 6684
rect 18911 6681 18923 6715
rect 18865 6675 18923 6681
rect 17114 6644 17120 6656
rect 14863 6616 17120 6644
rect 14863 6613 14875 6616
rect 14817 6607 14875 6613
rect 17114 6604 17120 6616
rect 17172 6604 17178 6656
rect 18678 6644 18684 6656
rect 18639 6616 18684 6644
rect 18678 6604 18684 6616
rect 18736 6644 18742 6656
rect 19340 6644 19368 6743
rect 19414 6740 19420 6792
rect 19472 6780 19478 6792
rect 19472 6752 19517 6780
rect 19472 6740 19478 6752
rect 20886 6740 20892 6792
rect 20944 6780 20950 6792
rect 21073 6783 21131 6789
rect 21073 6780 21085 6783
rect 20944 6752 21085 6780
rect 20944 6740 20950 6752
rect 21073 6749 21085 6752
rect 21119 6749 21131 6783
rect 21073 6743 21131 6749
rect 21165 6783 21223 6789
rect 21165 6749 21177 6783
rect 21211 6749 21223 6783
rect 21165 6743 21223 6749
rect 20334 6672 20340 6724
rect 20392 6712 20398 6724
rect 20429 6715 20487 6721
rect 20429 6712 20441 6715
rect 20392 6684 20441 6712
rect 20392 6672 20398 6684
rect 20429 6681 20441 6684
rect 20475 6712 20487 6715
rect 21180 6712 21208 6743
rect 22082 6740 22088 6792
rect 22140 6780 22146 6792
rect 22269 6783 22327 6789
rect 22269 6780 22281 6783
rect 22140 6752 22281 6780
rect 22140 6740 22146 6752
rect 22269 6749 22281 6752
rect 22315 6749 22327 6783
rect 22269 6743 22327 6749
rect 20475 6684 21208 6712
rect 20475 6681 20487 6684
rect 20429 6675 20487 6681
rect 23370 6672 23376 6724
rect 23428 6712 23434 6724
rect 24014 6712 24020 6724
rect 23428 6684 24020 6712
rect 23428 6672 23434 6684
rect 24014 6672 24020 6684
rect 24072 6712 24078 6724
rect 24201 6715 24259 6721
rect 24201 6712 24213 6715
rect 24072 6684 24213 6712
rect 24072 6672 24078 6684
rect 24201 6681 24213 6684
rect 24247 6712 24259 6715
rect 24842 6712 24848 6724
rect 24247 6684 24848 6712
rect 24247 6681 24259 6684
rect 24201 6675 24259 6681
rect 24842 6672 24848 6684
rect 24900 6672 24906 6724
rect 21806 6644 21812 6656
rect 18736 6616 19368 6644
rect 21767 6616 21812 6644
rect 18736 6604 18742 6616
rect 21806 6604 21812 6616
rect 21864 6604 21870 6656
rect 22174 6644 22180 6656
rect 22135 6616 22180 6644
rect 22174 6604 22180 6616
rect 22232 6604 22238 6656
rect 23646 6644 23652 6656
rect 23607 6616 23652 6644
rect 23646 6604 23652 6616
rect 23704 6604 23710 6656
rect 24934 6644 24940 6656
rect 24895 6616 24940 6644
rect 24934 6604 24940 6616
rect 24992 6604 24998 6656
rect 816 6554 26576 6576
rect 816 6502 5360 6554
rect 5412 6502 5424 6554
rect 5476 6502 5488 6554
rect 5540 6502 5552 6554
rect 5604 6502 14694 6554
rect 14746 6502 14758 6554
rect 14810 6502 14822 6554
rect 14874 6502 14886 6554
rect 14938 6502 24027 6554
rect 24079 6502 24091 6554
rect 24143 6502 24155 6554
rect 24207 6502 24219 6554
rect 24271 6502 26576 6554
rect 816 6480 26576 6502
rect 6902 6440 6908 6452
rect 6863 6412 6908 6440
rect 6902 6400 6908 6412
rect 6960 6400 6966 6452
rect 9754 6400 9760 6452
rect 9812 6440 9818 6452
rect 10033 6443 10091 6449
rect 10033 6440 10045 6443
rect 9812 6412 10045 6440
rect 9812 6400 9818 6412
rect 10033 6409 10045 6412
rect 10079 6409 10091 6443
rect 12238 6440 12244 6452
rect 12199 6412 12244 6440
rect 10033 6403 10091 6409
rect 12238 6400 12244 6412
rect 12296 6400 12302 6452
rect 13345 6443 13403 6449
rect 13345 6409 13357 6443
rect 13391 6440 13403 6443
rect 15185 6443 15243 6449
rect 15185 6440 15197 6443
rect 13391 6412 15197 6440
rect 13391 6409 13403 6412
rect 13345 6403 13403 6409
rect 15185 6409 15197 6412
rect 15231 6409 15243 6443
rect 15185 6403 15243 6409
rect 17209 6443 17267 6449
rect 17209 6409 17221 6443
rect 17255 6440 17267 6443
rect 17298 6440 17304 6452
rect 17255 6412 17304 6440
rect 17255 6409 17267 6412
rect 17209 6403 17267 6409
rect 12882 6304 12888 6316
rect 12795 6276 12888 6304
rect 12882 6264 12888 6276
rect 12940 6304 12946 6316
rect 13360 6304 13388 6403
rect 12940 6276 13388 6304
rect 12940 6264 12946 6276
rect 7273 6239 7331 6245
rect 7273 6205 7285 6239
rect 7319 6236 7331 6239
rect 7641 6239 7699 6245
rect 7641 6236 7653 6239
rect 7319 6208 7653 6236
rect 7319 6205 7331 6208
rect 7273 6199 7331 6205
rect 7641 6205 7653 6208
rect 7687 6236 7699 6239
rect 7822 6236 7828 6248
rect 7687 6208 7828 6236
rect 7687 6205 7699 6208
rect 7641 6199 7699 6205
rect 7822 6196 7828 6208
rect 7880 6236 7886 6248
rect 8098 6236 8104 6248
rect 7880 6208 8104 6236
rect 7880 6196 7886 6208
rect 8098 6196 8104 6208
rect 8156 6236 8162 6248
rect 9202 6236 9208 6248
rect 8156 6208 9208 6236
rect 8156 6196 8162 6208
rect 9202 6196 9208 6208
rect 9260 6196 9266 6248
rect 13802 6236 13808 6248
rect 13763 6208 13808 6236
rect 13802 6196 13808 6208
rect 13860 6196 13866 6248
rect 15826 6236 15832 6248
rect 15787 6208 15832 6236
rect 15826 6196 15832 6208
rect 15884 6196 15890 6248
rect 16565 6239 16623 6245
rect 16565 6205 16577 6239
rect 16611 6236 16623 6239
rect 17224 6236 17252 6403
rect 17298 6400 17304 6412
rect 17356 6400 17362 6452
rect 18494 6440 18500 6452
rect 18455 6412 18500 6440
rect 18494 6400 18500 6412
rect 18552 6400 18558 6452
rect 20334 6440 20340 6452
rect 20295 6412 20340 6440
rect 20334 6400 20340 6412
rect 20392 6400 20398 6452
rect 20886 6440 20892 6452
rect 20847 6412 20892 6440
rect 20886 6400 20892 6412
rect 20944 6400 20950 6452
rect 21530 6440 21536 6452
rect 21491 6412 21536 6440
rect 21530 6400 21536 6412
rect 21588 6400 21594 6452
rect 21714 6440 21720 6452
rect 21675 6412 21720 6440
rect 21714 6400 21720 6412
rect 21772 6400 21778 6452
rect 22542 6400 22548 6452
rect 22600 6440 22606 6452
rect 22729 6443 22787 6449
rect 22729 6440 22741 6443
rect 22600 6412 22741 6440
rect 22600 6400 22606 6412
rect 22729 6409 22741 6412
rect 22775 6409 22787 6443
rect 22729 6403 22787 6409
rect 24566 6400 24572 6452
rect 24624 6440 24630 6452
rect 25397 6443 25455 6449
rect 25397 6440 25409 6443
rect 24624 6412 25409 6440
rect 24624 6400 24630 6412
rect 25397 6409 25409 6412
rect 25443 6409 25455 6443
rect 25397 6403 25455 6409
rect 24842 6372 24848 6384
rect 24803 6344 24848 6372
rect 24842 6332 24848 6344
rect 24900 6332 24906 6384
rect 22174 6264 22180 6316
rect 22232 6304 22238 6316
rect 22361 6307 22419 6313
rect 22361 6304 22373 6307
rect 22232 6276 22373 6304
rect 22232 6264 22238 6276
rect 22361 6273 22373 6276
rect 22407 6304 22419 6307
rect 22407 6276 23140 6304
rect 22407 6273 22419 6276
rect 22361 6267 22419 6273
rect 16611 6208 17252 6236
rect 17853 6239 17911 6245
rect 16611 6205 16623 6208
rect 16565 6199 16623 6205
rect 17853 6205 17865 6239
rect 17899 6236 17911 6239
rect 18494 6236 18500 6248
rect 17899 6208 18500 6236
rect 17899 6205 17911 6208
rect 17853 6199 17911 6205
rect 18494 6196 18500 6208
rect 18552 6196 18558 6248
rect 18954 6236 18960 6248
rect 18788 6208 18960 6236
rect 8009 6171 8067 6177
rect 8009 6137 8021 6171
rect 8055 6168 8067 6171
rect 8346 6171 8404 6177
rect 8346 6168 8358 6171
rect 8055 6140 8358 6168
rect 8055 6137 8067 6140
rect 8009 6131 8067 6137
rect 8346 6137 8358 6140
rect 8392 6168 8404 6171
rect 9294 6168 9300 6180
rect 8392 6140 9300 6168
rect 8392 6137 8404 6140
rect 8346 6131 8404 6137
rect 9294 6128 9300 6140
rect 9352 6128 9358 6180
rect 9386 6128 9392 6180
rect 9444 6168 9450 6180
rect 9662 6168 9668 6180
rect 9444 6140 9668 6168
rect 9444 6128 9450 6140
rect 9662 6128 9668 6140
rect 9720 6168 9726 6180
rect 10401 6171 10459 6177
rect 10401 6168 10413 6171
rect 9720 6140 10413 6168
rect 9720 6128 9726 6140
rect 10401 6137 10413 6140
rect 10447 6137 10459 6171
rect 10401 6131 10459 6137
rect 10953 6171 11011 6177
rect 10953 6137 10965 6171
rect 10999 6168 11011 6171
rect 14050 6171 14108 6177
rect 14050 6168 14062 6171
rect 10999 6140 12744 6168
rect 10999 6137 11011 6140
rect 10953 6131 11011 6137
rect 12716 6112 12744 6140
rect 13636 6140 14062 6168
rect 13636 6112 13664 6140
rect 14050 6137 14062 6140
rect 14096 6137 14108 6171
rect 14050 6131 14108 6137
rect 16654 6128 16660 6180
rect 16712 6168 16718 6180
rect 17482 6168 17488 6180
rect 16712 6140 17488 6168
rect 16712 6128 16718 6140
rect 17482 6128 17488 6140
rect 17540 6128 17546 6180
rect 18788 6168 18816 6208
rect 18954 6196 18960 6208
rect 19012 6196 19018 6248
rect 17868 6140 18816 6168
rect 18865 6171 18923 6177
rect 9478 6100 9484 6112
rect 9439 6072 9484 6100
rect 9478 6060 9484 6072
rect 9536 6060 9542 6112
rect 11042 6100 11048 6112
rect 11003 6072 11048 6100
rect 11042 6060 11048 6072
rect 11100 6060 11106 6112
rect 11502 6100 11508 6112
rect 11463 6072 11508 6100
rect 11502 6060 11508 6072
rect 11560 6060 11566 6112
rect 11965 6103 12023 6109
rect 11965 6069 11977 6103
rect 12011 6100 12023 6103
rect 12606 6100 12612 6112
rect 12011 6072 12612 6100
rect 12011 6069 12023 6072
rect 11965 6063 12023 6069
rect 12606 6060 12612 6072
rect 12664 6060 12670 6112
rect 12698 6060 12704 6112
rect 12756 6100 12762 6112
rect 13618 6100 13624 6112
rect 12756 6072 12801 6100
rect 13579 6072 13624 6100
rect 12756 6060 12762 6072
rect 13618 6060 13624 6072
rect 13676 6060 13682 6112
rect 16102 6100 16108 6112
rect 16063 6072 16108 6100
rect 16102 6060 16108 6072
rect 16160 6060 16166 6112
rect 16746 6100 16752 6112
rect 16707 6072 16752 6100
rect 16746 6060 16752 6072
rect 16804 6060 16810 6112
rect 17114 6060 17120 6112
rect 17172 6100 17178 6112
rect 17868 6100 17896 6140
rect 18865 6137 18877 6171
rect 18911 6168 18923 6171
rect 19046 6168 19052 6180
rect 18911 6140 19052 6168
rect 18911 6137 18923 6140
rect 18865 6131 18923 6137
rect 19046 6128 19052 6140
rect 19104 6168 19110 6180
rect 19224 6171 19282 6177
rect 19224 6168 19236 6171
rect 19104 6140 19236 6168
rect 19104 6128 19110 6140
rect 19224 6137 19236 6140
rect 19270 6168 19282 6171
rect 19414 6168 19420 6180
rect 19270 6140 19420 6168
rect 19270 6137 19282 6140
rect 19224 6131 19282 6137
rect 19414 6128 19420 6140
rect 19472 6128 19478 6180
rect 21806 6128 21812 6180
rect 21864 6168 21870 6180
rect 22085 6171 22143 6177
rect 22085 6168 22097 6171
rect 21864 6140 22097 6168
rect 21864 6128 21870 6140
rect 22085 6137 22097 6140
rect 22131 6168 22143 6171
rect 22266 6168 22272 6180
rect 22131 6140 22272 6168
rect 22131 6137 22143 6140
rect 22085 6131 22143 6137
rect 22266 6128 22272 6140
rect 22324 6128 22330 6180
rect 23112 6168 23140 6276
rect 23278 6196 23284 6248
rect 23336 6236 23342 6248
rect 23465 6239 23523 6245
rect 23465 6236 23477 6239
rect 23336 6208 23477 6236
rect 23336 6196 23342 6208
rect 23465 6205 23477 6208
rect 23511 6205 23523 6239
rect 23465 6199 23523 6205
rect 23646 6168 23652 6180
rect 23112 6140 23652 6168
rect 23112 6112 23140 6140
rect 23646 6128 23652 6140
rect 23704 6177 23710 6180
rect 23704 6171 23768 6177
rect 23704 6137 23722 6171
rect 23756 6137 23768 6171
rect 23704 6131 23768 6137
rect 23704 6128 23710 6131
rect 18034 6100 18040 6112
rect 17172 6072 17896 6100
rect 17995 6072 18040 6100
rect 17172 6060 17178 6072
rect 18034 6060 18040 6072
rect 18092 6060 18098 6112
rect 21530 6060 21536 6112
rect 21588 6100 21594 6112
rect 22174 6100 22180 6112
rect 21588 6072 22180 6100
rect 21588 6060 21594 6072
rect 22174 6060 22180 6072
rect 22232 6060 22238 6112
rect 23094 6100 23100 6112
rect 23055 6072 23100 6100
rect 23094 6060 23100 6072
rect 23152 6060 23158 6112
rect 25857 6103 25915 6109
rect 25857 6069 25869 6103
rect 25903 6100 25915 6103
rect 25946 6100 25952 6112
rect 25903 6072 25952 6100
rect 25903 6069 25915 6072
rect 25857 6063 25915 6069
rect 25946 6060 25952 6072
rect 26004 6100 26010 6112
rect 26133 6103 26191 6109
rect 26133 6100 26145 6103
rect 26004 6072 26145 6100
rect 26004 6060 26010 6072
rect 26133 6069 26145 6072
rect 26179 6069 26191 6103
rect 26133 6063 26191 6069
rect 816 6010 26576 6032
rect 816 5958 10027 6010
rect 10079 5958 10091 6010
rect 10143 5958 10155 6010
rect 10207 5958 10219 6010
rect 10271 5958 19360 6010
rect 19412 5958 19424 6010
rect 19476 5958 19488 6010
rect 19540 5958 19552 6010
rect 19604 5958 26576 6010
rect 816 5936 26576 5958
rect 6902 5856 6908 5908
rect 6960 5896 6966 5908
rect 8745 5899 8803 5905
rect 8745 5896 8757 5899
rect 6960 5868 8757 5896
rect 6960 5856 6966 5868
rect 8745 5865 8757 5868
rect 8791 5896 8803 5899
rect 9110 5896 9116 5908
rect 8791 5868 9116 5896
rect 8791 5865 8803 5868
rect 8745 5859 8803 5865
rect 9110 5856 9116 5868
rect 9168 5896 9174 5908
rect 9478 5896 9484 5908
rect 9168 5868 9484 5896
rect 9168 5856 9174 5868
rect 9478 5856 9484 5868
rect 9536 5856 9542 5908
rect 9570 5856 9576 5908
rect 9628 5896 9634 5908
rect 9846 5896 9852 5908
rect 9628 5868 9673 5896
rect 9807 5868 9852 5896
rect 9628 5856 9634 5868
rect 9846 5856 9852 5868
rect 9904 5856 9910 5908
rect 10217 5899 10275 5905
rect 10217 5865 10229 5899
rect 10263 5896 10275 5899
rect 11042 5896 11048 5908
rect 10263 5868 11048 5896
rect 10263 5865 10275 5868
rect 10217 5859 10275 5865
rect 9662 5788 9668 5840
rect 9720 5828 9726 5840
rect 10232 5828 10260 5859
rect 11042 5856 11048 5868
rect 11100 5856 11106 5908
rect 12606 5856 12612 5908
rect 12664 5896 12670 5908
rect 13897 5899 13955 5905
rect 13897 5896 13909 5899
rect 12664 5868 13909 5896
rect 12664 5856 12670 5868
rect 13897 5865 13909 5868
rect 13943 5865 13955 5899
rect 13897 5859 13955 5865
rect 14538 5856 14544 5908
rect 14596 5896 14602 5908
rect 14725 5899 14783 5905
rect 14725 5896 14737 5899
rect 14596 5868 14737 5896
rect 14596 5856 14602 5868
rect 14725 5865 14737 5868
rect 14771 5865 14783 5899
rect 15550 5896 15556 5908
rect 15511 5868 15556 5896
rect 14725 5859 14783 5865
rect 15550 5856 15556 5868
rect 15608 5856 15614 5908
rect 17117 5899 17175 5905
rect 17117 5865 17129 5899
rect 17163 5896 17175 5899
rect 17574 5896 17580 5908
rect 17163 5868 17580 5896
rect 17163 5865 17175 5868
rect 17117 5859 17175 5865
rect 17574 5856 17580 5868
rect 17632 5856 17638 5908
rect 18957 5899 19015 5905
rect 18957 5865 18969 5899
rect 19003 5896 19015 5899
rect 19046 5896 19052 5908
rect 19003 5868 19052 5896
rect 19003 5865 19015 5868
rect 18957 5859 19015 5865
rect 19046 5856 19052 5868
rect 19104 5896 19110 5908
rect 19509 5899 19567 5905
rect 19509 5896 19521 5899
rect 19104 5868 19521 5896
rect 19104 5856 19110 5868
rect 19509 5865 19521 5868
rect 19555 5865 19567 5899
rect 19874 5896 19880 5908
rect 19835 5868 19880 5896
rect 19509 5859 19567 5865
rect 19874 5856 19880 5868
rect 19932 5856 19938 5908
rect 21438 5856 21444 5908
rect 21496 5896 21502 5908
rect 21993 5899 22051 5905
rect 21993 5896 22005 5899
rect 21496 5868 22005 5896
rect 21496 5856 21502 5868
rect 21993 5865 22005 5868
rect 22039 5865 22051 5899
rect 21993 5859 22051 5865
rect 23370 5856 23376 5908
rect 23428 5896 23434 5908
rect 23428 5868 23692 5896
rect 23428 5856 23434 5868
rect 23664 5840 23692 5868
rect 11318 5828 11324 5840
rect 9720 5800 10260 5828
rect 11231 5800 11324 5828
rect 9720 5788 9726 5800
rect 11318 5788 11324 5800
rect 11376 5828 11382 5840
rect 12054 5828 12060 5840
rect 11376 5800 12060 5828
rect 11376 5788 11382 5800
rect 12054 5788 12060 5800
rect 12112 5788 12118 5840
rect 17850 5837 17856 5840
rect 17844 5828 17856 5837
rect 17811 5800 17856 5828
rect 17844 5791 17856 5800
rect 17850 5788 17856 5791
rect 17908 5788 17914 5840
rect 20334 5788 20340 5840
rect 20392 5828 20398 5840
rect 20858 5831 20916 5837
rect 20858 5828 20870 5831
rect 20392 5800 20870 5828
rect 20392 5788 20398 5800
rect 20858 5797 20870 5800
rect 20904 5797 20916 5831
rect 20858 5791 20916 5797
rect 23646 5788 23652 5840
rect 23704 5837 23710 5840
rect 23704 5831 23768 5837
rect 23704 5797 23722 5831
rect 23756 5797 23768 5831
rect 23704 5791 23768 5797
rect 23704 5788 23710 5791
rect 8006 5720 8012 5772
rect 8064 5760 8070 5772
rect 8101 5763 8159 5769
rect 8101 5760 8113 5763
rect 8064 5732 8113 5760
rect 8064 5720 8070 5732
rect 8101 5729 8113 5732
rect 8147 5729 8159 5763
rect 8101 5723 8159 5729
rect 9294 5720 9300 5772
rect 9352 5760 9358 5772
rect 9846 5760 9852 5772
rect 9352 5732 9852 5760
rect 9352 5720 9358 5732
rect 9846 5720 9852 5732
rect 9904 5760 9910 5772
rect 9904 5732 10444 5760
rect 9904 5720 9910 5732
rect 7914 5652 7920 5704
rect 7972 5692 7978 5704
rect 8190 5692 8196 5704
rect 7972 5664 8196 5692
rect 7972 5652 7978 5664
rect 8190 5652 8196 5664
rect 8248 5652 8254 5704
rect 8285 5695 8343 5701
rect 8285 5661 8297 5695
rect 8331 5661 8343 5695
rect 8285 5655 8343 5661
rect 9205 5695 9263 5701
rect 9205 5661 9217 5695
rect 9251 5692 9263 5695
rect 10306 5692 10312 5704
rect 9251 5664 10312 5692
rect 9251 5661 9263 5664
rect 9205 5655 9263 5661
rect 7730 5624 7736 5636
rect 7691 5596 7736 5624
rect 7730 5584 7736 5596
rect 7788 5584 7794 5636
rect 7822 5584 7828 5636
rect 7880 5624 7886 5636
rect 8300 5624 8328 5655
rect 10306 5652 10312 5664
rect 10364 5652 10370 5704
rect 10416 5701 10444 5732
rect 11042 5720 11048 5772
rect 11100 5760 11106 5772
rect 11669 5763 11727 5769
rect 11669 5760 11681 5763
rect 11100 5732 11681 5760
rect 11100 5720 11106 5732
rect 11669 5729 11681 5732
rect 11715 5729 11727 5763
rect 14998 5760 15004 5772
rect 14959 5732 15004 5760
rect 11669 5723 11727 5729
rect 14998 5720 15004 5732
rect 15056 5720 15062 5772
rect 16378 5760 16384 5772
rect 16291 5732 16384 5760
rect 16378 5720 16384 5732
rect 16436 5760 16442 5772
rect 17298 5760 17304 5772
rect 16436 5732 17304 5760
rect 16436 5720 16442 5732
rect 17298 5720 17304 5732
rect 17356 5720 17362 5772
rect 22082 5760 22088 5772
rect 20628 5732 22088 5760
rect 20628 5704 20656 5732
rect 22082 5720 22088 5732
rect 22140 5760 22146 5772
rect 22140 5732 23324 5760
rect 22140 5720 22146 5732
rect 23296 5704 23324 5732
rect 10401 5695 10459 5701
rect 10401 5661 10413 5695
rect 10447 5661 10459 5695
rect 11410 5692 11416 5704
rect 11371 5664 11416 5692
rect 10401 5655 10459 5661
rect 7880 5596 8328 5624
rect 10416 5624 10444 5655
rect 11410 5652 11416 5664
rect 11468 5652 11474 5704
rect 16470 5692 16476 5704
rect 16431 5664 16476 5692
rect 16470 5652 16476 5664
rect 16528 5652 16534 5704
rect 16562 5652 16568 5704
rect 16620 5692 16626 5704
rect 16620 5664 16665 5692
rect 16620 5652 16626 5664
rect 17114 5652 17120 5704
rect 17172 5692 17178 5704
rect 17577 5695 17635 5701
rect 17577 5692 17589 5695
rect 17172 5664 17589 5692
rect 17172 5652 17178 5664
rect 17577 5661 17589 5664
rect 17623 5661 17635 5695
rect 20610 5692 20616 5704
rect 20571 5664 20616 5692
rect 17577 5655 17635 5661
rect 20610 5652 20616 5664
rect 20668 5652 20674 5704
rect 22542 5692 22548 5704
rect 22503 5664 22548 5692
rect 22542 5652 22548 5664
rect 22600 5652 22606 5704
rect 23278 5692 23284 5704
rect 23191 5664 23284 5692
rect 23278 5652 23284 5664
rect 23336 5692 23342 5704
rect 23465 5695 23523 5701
rect 23465 5692 23477 5695
rect 23336 5664 23477 5692
rect 23336 5652 23342 5664
rect 23465 5661 23477 5664
rect 23511 5661 23523 5695
rect 23465 5655 23523 5661
rect 10416 5596 11364 5624
rect 7880 5584 7886 5596
rect 10953 5559 11011 5565
rect 10953 5525 10965 5559
rect 10999 5556 11011 5559
rect 11042 5556 11048 5568
rect 10999 5528 11048 5556
rect 10999 5525 11011 5528
rect 10953 5519 11011 5525
rect 11042 5516 11048 5528
rect 11100 5516 11106 5568
rect 11336 5556 11364 5596
rect 12606 5584 12612 5636
rect 12664 5624 12670 5636
rect 13345 5627 13403 5633
rect 13345 5624 13357 5627
rect 12664 5596 13357 5624
rect 12664 5584 12670 5596
rect 13345 5593 13357 5596
rect 13391 5624 13403 5627
rect 13713 5627 13771 5633
rect 13713 5624 13725 5627
rect 13391 5596 13725 5624
rect 13391 5593 13403 5596
rect 13345 5587 13403 5593
rect 13713 5593 13725 5596
rect 13759 5624 13771 5627
rect 13802 5624 13808 5636
rect 13759 5596 13808 5624
rect 13759 5593 13771 5596
rect 13713 5587 13771 5593
rect 13802 5584 13808 5596
rect 13860 5624 13866 5636
rect 14170 5624 14176 5636
rect 13860 5596 14176 5624
rect 13860 5584 13866 5596
rect 14170 5584 14176 5596
rect 14228 5624 14234 5636
rect 14357 5627 14415 5633
rect 14357 5624 14369 5627
rect 14228 5596 14369 5624
rect 14228 5584 14234 5596
rect 14357 5593 14369 5596
rect 14403 5593 14415 5627
rect 14357 5587 14415 5593
rect 16013 5627 16071 5633
rect 16013 5593 16025 5627
rect 16059 5624 16071 5627
rect 17393 5627 17451 5633
rect 17393 5624 17405 5627
rect 16059 5596 17405 5624
rect 16059 5593 16071 5596
rect 16013 5587 16071 5593
rect 17393 5593 17405 5596
rect 17439 5593 17451 5627
rect 17393 5587 17451 5593
rect 12793 5559 12851 5565
rect 12793 5556 12805 5559
rect 11336 5528 12805 5556
rect 12793 5525 12805 5528
rect 12839 5525 12851 5559
rect 17408 5556 17436 5587
rect 17758 5556 17764 5568
rect 17408 5528 17764 5556
rect 12793 5519 12851 5525
rect 17758 5516 17764 5528
rect 17816 5516 17822 5568
rect 20429 5559 20487 5565
rect 20429 5525 20441 5559
rect 20475 5556 20487 5559
rect 20978 5556 20984 5568
rect 20475 5528 20984 5556
rect 20475 5525 20487 5528
rect 20429 5519 20487 5525
rect 20978 5516 20984 5528
rect 21036 5556 21042 5568
rect 21530 5556 21536 5568
rect 21036 5528 21536 5556
rect 21036 5516 21042 5528
rect 21530 5516 21536 5528
rect 21588 5516 21594 5568
rect 22910 5556 22916 5568
rect 22871 5528 22916 5556
rect 22910 5516 22916 5528
rect 22968 5556 22974 5568
rect 23296 5565 23324 5652
rect 23281 5559 23339 5565
rect 23281 5556 23293 5559
rect 22968 5528 23293 5556
rect 22968 5516 22974 5528
rect 23281 5525 23293 5528
rect 23327 5525 23339 5559
rect 23281 5519 23339 5525
rect 24474 5516 24480 5568
rect 24532 5556 24538 5568
rect 24845 5559 24903 5565
rect 24845 5556 24857 5559
rect 24532 5528 24857 5556
rect 24532 5516 24538 5528
rect 24845 5525 24857 5528
rect 24891 5525 24903 5559
rect 24845 5519 24903 5525
rect 816 5466 26576 5488
rect 816 5414 5360 5466
rect 5412 5414 5424 5466
rect 5476 5414 5488 5466
rect 5540 5414 5552 5466
rect 5604 5414 14694 5466
rect 14746 5414 14758 5466
rect 14810 5414 14822 5466
rect 14874 5414 14886 5466
rect 14938 5414 24027 5466
rect 24079 5414 24091 5466
rect 24143 5414 24155 5466
rect 24207 5414 24219 5466
rect 24271 5414 26576 5466
rect 816 5392 26576 5414
rect 7457 5355 7515 5361
rect 7457 5321 7469 5355
rect 7503 5352 7515 5355
rect 7914 5352 7920 5364
rect 7503 5324 7920 5352
rect 7503 5321 7515 5324
rect 7457 5315 7515 5321
rect 7914 5312 7920 5324
rect 7972 5312 7978 5364
rect 8561 5355 8619 5361
rect 8561 5321 8573 5355
rect 8607 5352 8619 5355
rect 9386 5352 9392 5364
rect 8607 5324 9392 5352
rect 8607 5321 8619 5324
rect 8561 5315 8619 5321
rect 9386 5312 9392 5324
rect 9444 5312 9450 5364
rect 9662 5352 9668 5364
rect 9623 5324 9668 5352
rect 9662 5312 9668 5324
rect 9720 5312 9726 5364
rect 10306 5312 10312 5364
rect 10364 5352 10370 5364
rect 10493 5355 10551 5361
rect 10493 5352 10505 5355
rect 10364 5324 10505 5352
rect 10364 5312 10370 5324
rect 10493 5321 10505 5324
rect 10539 5321 10551 5355
rect 13529 5355 13587 5361
rect 13529 5352 13541 5355
rect 10493 5315 10551 5321
rect 11520 5324 13541 5352
rect 7549 5219 7607 5225
rect 7549 5185 7561 5219
rect 7595 5216 7607 5219
rect 7638 5216 7644 5228
rect 7595 5188 7644 5216
rect 7595 5185 7607 5188
rect 7549 5179 7607 5185
rect 7638 5176 7644 5188
rect 7696 5176 7702 5228
rect 9110 5216 9116 5228
rect 9071 5188 9116 5216
rect 9110 5176 9116 5188
rect 9168 5176 9174 5228
rect 11042 5216 11048 5228
rect 11003 5188 11048 5216
rect 11042 5176 11048 5188
rect 11100 5216 11106 5228
rect 11520 5225 11548 5324
rect 13529 5321 13541 5324
rect 13575 5321 13587 5355
rect 14170 5352 14176 5364
rect 14131 5324 14176 5352
rect 13529 5315 13587 5321
rect 14170 5312 14176 5324
rect 14228 5312 14234 5364
rect 17209 5355 17267 5361
rect 17209 5321 17221 5355
rect 17255 5352 17267 5355
rect 17298 5352 17304 5364
rect 17255 5324 17304 5352
rect 17255 5321 17267 5324
rect 17209 5315 17267 5321
rect 17298 5312 17304 5324
rect 17356 5312 17362 5364
rect 17482 5352 17488 5364
rect 17443 5324 17488 5352
rect 17482 5312 17488 5324
rect 17540 5312 17546 5364
rect 17761 5355 17819 5361
rect 17761 5321 17773 5355
rect 17807 5352 17819 5355
rect 18678 5352 18684 5364
rect 17807 5324 18684 5352
rect 17807 5321 17819 5324
rect 17761 5315 17819 5321
rect 18678 5312 18684 5324
rect 18736 5312 18742 5364
rect 19046 5312 19052 5364
rect 19104 5352 19110 5364
rect 19325 5355 19383 5361
rect 19325 5352 19337 5355
rect 19104 5324 19337 5352
rect 19104 5312 19110 5324
rect 19325 5321 19337 5324
rect 19371 5321 19383 5355
rect 19325 5315 19383 5321
rect 17850 5244 17856 5296
rect 17908 5284 17914 5296
rect 18773 5287 18831 5293
rect 18773 5284 18785 5287
rect 17908 5256 18785 5284
rect 17908 5244 17914 5256
rect 18328 5228 18356 5256
rect 18773 5253 18785 5256
rect 18819 5253 18831 5287
rect 18773 5247 18831 5253
rect 11505 5219 11563 5225
rect 11505 5216 11517 5219
rect 11100 5188 11517 5216
rect 11100 5176 11106 5188
rect 11505 5185 11517 5188
rect 11551 5185 11563 5219
rect 11505 5179 11563 5185
rect 11965 5219 12023 5225
rect 11965 5185 11977 5219
rect 12011 5216 12023 5219
rect 12011 5188 12284 5216
rect 12011 5185 12023 5188
rect 11965 5179 12023 5185
rect 11318 5108 11324 5160
rect 11376 5148 11382 5160
rect 12149 5151 12207 5157
rect 12149 5148 12161 5151
rect 11376 5120 12161 5148
rect 11376 5108 11382 5120
rect 12149 5117 12161 5120
rect 12195 5117 12207 5151
rect 12256 5148 12284 5188
rect 14170 5176 14176 5228
rect 14228 5216 14234 5228
rect 15185 5219 15243 5225
rect 15185 5216 15197 5219
rect 14228 5188 15197 5216
rect 14228 5176 14234 5188
rect 15185 5185 15197 5188
rect 15231 5185 15243 5219
rect 15185 5179 15243 5185
rect 17758 5176 17764 5228
rect 17816 5216 17822 5228
rect 18221 5219 18279 5225
rect 18221 5216 18233 5219
rect 17816 5188 18233 5216
rect 17816 5176 17822 5188
rect 18221 5185 18233 5188
rect 18267 5185 18279 5219
rect 18221 5179 18279 5185
rect 18310 5176 18316 5228
rect 18368 5216 18374 5228
rect 19340 5216 19368 5315
rect 20334 5312 20340 5364
rect 20392 5352 20398 5364
rect 20613 5355 20671 5361
rect 20613 5352 20625 5355
rect 20392 5324 20625 5352
rect 20392 5312 20398 5324
rect 20613 5321 20625 5324
rect 20659 5321 20671 5355
rect 20613 5315 20671 5321
rect 22177 5355 22235 5361
rect 22177 5321 22189 5355
rect 22223 5352 22235 5355
rect 22450 5352 22456 5364
rect 22223 5324 22456 5352
rect 22223 5321 22235 5324
rect 22177 5315 22235 5321
rect 22450 5312 22456 5324
rect 22508 5312 22514 5364
rect 23554 5352 23560 5364
rect 23515 5324 23560 5352
rect 23554 5312 23560 5324
rect 23612 5312 23618 5364
rect 24382 5312 24388 5364
rect 24440 5352 24446 5364
rect 25673 5355 25731 5361
rect 25673 5352 25685 5355
rect 24440 5324 25685 5352
rect 24440 5312 24446 5324
rect 24569 5287 24627 5293
rect 24569 5284 24581 5287
rect 24032 5256 24581 5284
rect 20242 5216 20248 5228
rect 18368 5188 18461 5216
rect 19340 5188 20248 5216
rect 18368 5176 18374 5188
rect 20242 5176 20248 5188
rect 20300 5216 20306 5228
rect 20610 5216 20616 5228
rect 20300 5188 20616 5216
rect 20300 5176 20306 5188
rect 20610 5176 20616 5188
rect 20668 5216 20674 5228
rect 20797 5219 20855 5225
rect 20797 5216 20809 5219
rect 20668 5188 20809 5216
rect 20668 5176 20674 5188
rect 20797 5185 20809 5188
rect 20843 5185 20855 5219
rect 20797 5179 20855 5185
rect 23189 5219 23247 5225
rect 23189 5185 23201 5219
rect 23235 5185 23247 5219
rect 23189 5179 23247 5185
rect 12416 5151 12474 5157
rect 12416 5148 12428 5151
rect 12256 5120 12428 5148
rect 12149 5111 12207 5117
rect 12416 5117 12428 5120
rect 12462 5148 12474 5151
rect 12882 5148 12888 5160
rect 12462 5120 12888 5148
rect 12462 5117 12474 5120
rect 12416 5111 12474 5117
rect 10033 5083 10091 5089
rect 10033 5049 10045 5083
rect 10079 5080 10091 5083
rect 10950 5080 10956 5092
rect 10079 5052 10956 5080
rect 10079 5049 10091 5052
rect 10033 5043 10091 5049
rect 10950 5040 10956 5052
rect 11008 5040 11014 5092
rect 12164 5080 12192 5111
rect 12882 5108 12888 5120
rect 12940 5108 12946 5160
rect 14354 5108 14360 5160
rect 14412 5148 14418 5160
rect 14541 5151 14599 5157
rect 14541 5148 14553 5151
rect 14412 5120 14553 5148
rect 14412 5108 14418 5120
rect 14541 5117 14553 5120
rect 14587 5148 14599 5151
rect 14817 5151 14875 5157
rect 14817 5148 14829 5151
rect 14587 5120 14829 5148
rect 14587 5117 14599 5120
rect 14541 5111 14599 5117
rect 14817 5117 14829 5120
rect 14863 5117 14875 5151
rect 14817 5111 14875 5117
rect 17666 5108 17672 5160
rect 17724 5148 17730 5160
rect 18129 5151 18187 5157
rect 18129 5148 18141 5151
rect 17724 5120 18141 5148
rect 17724 5108 17730 5120
rect 18129 5117 18141 5120
rect 18175 5117 18187 5151
rect 19506 5148 19512 5160
rect 19467 5120 19512 5148
rect 18129 5111 18187 5117
rect 19506 5108 19512 5120
rect 19564 5108 19570 5160
rect 19693 5151 19751 5157
rect 19693 5117 19705 5151
rect 19739 5148 19751 5151
rect 19874 5148 19880 5160
rect 19739 5120 19880 5148
rect 19739 5117 19751 5120
rect 19693 5111 19751 5117
rect 19874 5108 19880 5120
rect 19932 5108 19938 5160
rect 20337 5151 20395 5157
rect 20337 5117 20349 5151
rect 20383 5148 20395 5151
rect 21053 5151 21111 5157
rect 21053 5148 21065 5151
rect 20383 5120 21065 5148
rect 20383 5117 20395 5120
rect 20337 5111 20395 5117
rect 21053 5117 21065 5120
rect 21099 5148 21111 5151
rect 21438 5148 21444 5160
rect 21099 5120 21444 5148
rect 21099 5117 21111 5120
rect 21053 5111 21111 5117
rect 21438 5108 21444 5120
rect 21496 5108 21502 5160
rect 23204 5148 23232 5179
rect 23462 5176 23468 5228
rect 23520 5216 23526 5228
rect 24032 5225 24060 5256
rect 24569 5253 24581 5256
rect 24615 5253 24627 5287
rect 24569 5247 24627 5253
rect 24017 5219 24075 5225
rect 24017 5216 24029 5219
rect 23520 5188 24029 5216
rect 23520 5176 23526 5188
rect 24017 5185 24029 5188
rect 24063 5185 24075 5219
rect 24017 5179 24075 5185
rect 24201 5219 24259 5225
rect 24201 5185 24213 5219
rect 24247 5216 24259 5219
rect 24474 5216 24480 5228
rect 24247 5188 24480 5216
rect 24247 5185 24259 5188
rect 24201 5179 24259 5185
rect 23554 5148 23560 5160
rect 23204 5120 23560 5148
rect 23554 5108 23560 5120
rect 23612 5148 23618 5160
rect 24216 5148 24244 5179
rect 24474 5176 24480 5188
rect 24532 5176 24538 5228
rect 25136 5157 25164 5324
rect 25673 5321 25685 5324
rect 25719 5321 25731 5355
rect 25673 5315 25731 5321
rect 23612 5120 24244 5148
rect 25121 5151 25179 5157
rect 23612 5108 23618 5120
rect 25121 5117 25133 5151
rect 25167 5117 25179 5151
rect 25121 5111 25179 5117
rect 12606 5080 12612 5092
rect 12164 5052 12612 5080
rect 12606 5040 12612 5052
rect 12664 5040 12670 5092
rect 15274 5040 15280 5092
rect 15332 5080 15338 5092
rect 15430 5083 15488 5089
rect 15430 5080 15442 5083
rect 15332 5052 15442 5080
rect 15332 5040 15338 5052
rect 15430 5049 15442 5052
rect 15476 5049 15488 5083
rect 15430 5043 15488 5049
rect 16654 5040 16660 5092
rect 16712 5080 16718 5092
rect 16838 5080 16844 5092
rect 16712 5052 16844 5080
rect 16712 5040 16718 5052
rect 16838 5040 16844 5052
rect 16896 5040 16902 5092
rect 19138 5040 19144 5092
rect 19196 5080 19202 5092
rect 20058 5080 20064 5092
rect 19196 5052 20064 5080
rect 19196 5040 19202 5052
rect 20058 5040 20064 5052
rect 20116 5040 20122 5092
rect 23186 5040 23192 5092
rect 23244 5080 23250 5092
rect 23925 5083 23983 5089
rect 23925 5080 23937 5083
rect 23244 5052 23937 5080
rect 23244 5040 23250 5052
rect 23925 5049 23937 5052
rect 23971 5080 23983 5083
rect 24937 5083 24995 5089
rect 24937 5080 24949 5083
rect 23971 5052 24949 5080
rect 23971 5049 23983 5052
rect 23925 5043 23983 5049
rect 24937 5049 24949 5052
rect 24983 5049 24995 5083
rect 24937 5043 24995 5049
rect 8006 5012 8012 5024
rect 7967 4984 8012 5012
rect 8006 4972 8012 4984
rect 8064 4972 8070 5024
rect 8374 5012 8380 5024
rect 8335 4984 8380 5012
rect 8374 4972 8380 4984
rect 8432 5012 8438 5024
rect 8929 5015 8987 5021
rect 8929 5012 8941 5015
rect 8432 4984 8941 5012
rect 8432 4972 8438 4984
rect 8929 4981 8941 4984
rect 8975 4981 8987 5015
rect 8929 4975 8987 4981
rect 9021 5015 9079 5021
rect 9021 4981 9033 5015
rect 9067 5012 9079 5015
rect 9294 5012 9300 5024
rect 9067 4984 9300 5012
rect 9067 4981 9079 4984
rect 9021 4975 9079 4981
rect 9294 4972 9300 4984
rect 9352 4972 9358 5024
rect 9754 4972 9760 5024
rect 9812 5012 9818 5024
rect 10309 5015 10367 5021
rect 10309 5012 10321 5015
rect 9812 4984 10321 5012
rect 9812 4972 9818 4984
rect 10309 4981 10321 4984
rect 10355 5012 10367 5015
rect 10861 5015 10919 5021
rect 10861 5012 10873 5015
rect 10355 4984 10873 5012
rect 10355 4981 10367 4984
rect 10309 4975 10367 4981
rect 10861 4981 10873 4984
rect 10907 4981 10919 5015
rect 10861 4975 10919 4981
rect 14538 4972 14544 5024
rect 14596 5012 14602 5024
rect 14633 5015 14691 5021
rect 14633 5012 14645 5015
rect 14596 4984 14645 5012
rect 14596 4972 14602 4984
rect 14633 4981 14645 4984
rect 14679 4981 14691 5015
rect 16562 5012 16568 5024
rect 16523 4984 16568 5012
rect 14633 4975 14691 4981
rect 16562 4972 16568 4984
rect 16620 4972 16626 5024
rect 19230 5012 19236 5024
rect 19191 4984 19236 5012
rect 19230 4972 19236 4984
rect 19288 4972 19294 5024
rect 19874 5012 19880 5024
rect 19835 4984 19880 5012
rect 19874 4972 19880 4984
rect 19932 4972 19938 5024
rect 22821 5015 22879 5021
rect 22821 4981 22833 5015
rect 22867 5012 22879 5015
rect 23646 5012 23652 5024
rect 22867 4984 23652 5012
rect 22867 4981 22879 4984
rect 22821 4975 22879 4981
rect 23646 4972 23652 4984
rect 23704 4972 23710 5024
rect 25302 5012 25308 5024
rect 25263 4984 25308 5012
rect 25302 4972 25308 4984
rect 25360 4972 25366 5024
rect 25946 4972 25952 5024
rect 26004 5012 26010 5024
rect 26041 5015 26099 5021
rect 26041 5012 26053 5015
rect 26004 4984 26053 5012
rect 26004 4972 26010 4984
rect 26041 4981 26053 4984
rect 26087 4981 26099 5015
rect 26041 4975 26099 4981
rect 816 4922 26576 4944
rect 816 4870 10027 4922
rect 10079 4870 10091 4922
rect 10143 4870 10155 4922
rect 10207 4870 10219 4922
rect 10271 4870 19360 4922
rect 19412 4870 19424 4922
rect 19476 4870 19488 4922
rect 19540 4870 19552 4922
rect 19604 4870 26576 4922
rect 816 4848 26576 4870
rect 7822 4808 7828 4820
rect 7783 4780 7828 4808
rect 7822 4768 7828 4780
rect 7880 4768 7886 4820
rect 8098 4808 8104 4820
rect 8059 4780 8104 4808
rect 8098 4768 8104 4780
rect 8156 4768 8162 4820
rect 9846 4808 9852 4820
rect 9807 4780 9852 4808
rect 9846 4768 9852 4780
rect 9904 4768 9910 4820
rect 11502 4808 11508 4820
rect 11463 4780 11508 4808
rect 11502 4768 11508 4780
rect 11560 4768 11566 4820
rect 12698 4768 12704 4820
rect 12756 4808 12762 4820
rect 13345 4811 13403 4817
rect 13345 4808 13357 4811
rect 12756 4780 13357 4808
rect 12756 4768 12762 4780
rect 13345 4777 13357 4780
rect 13391 4777 13403 4811
rect 13345 4771 13403 4777
rect 14170 4768 14176 4820
rect 14228 4808 14234 4820
rect 14357 4811 14415 4817
rect 14357 4808 14369 4811
rect 14228 4780 14369 4808
rect 14228 4768 14234 4780
rect 14357 4777 14369 4780
rect 14403 4777 14415 4811
rect 15274 4808 15280 4820
rect 15235 4780 15280 4808
rect 14357 4771 14415 4777
rect 15274 4768 15280 4780
rect 15332 4768 15338 4820
rect 15642 4808 15648 4820
rect 15603 4780 15648 4808
rect 15642 4768 15648 4780
rect 15700 4768 15706 4820
rect 16105 4811 16163 4817
rect 16105 4777 16117 4811
rect 16151 4808 16163 4811
rect 16194 4808 16200 4820
rect 16151 4780 16200 4808
rect 16151 4777 16163 4780
rect 16105 4771 16163 4777
rect 14538 4740 14544 4752
rect 12900 4712 14544 4740
rect 10392 4675 10450 4681
rect 10392 4641 10404 4675
rect 10438 4672 10450 4675
rect 10674 4672 10680 4684
rect 10438 4644 10680 4672
rect 10438 4641 10450 4644
rect 10392 4635 10450 4641
rect 10674 4632 10680 4644
rect 10732 4632 10738 4684
rect 12054 4632 12060 4684
rect 12112 4672 12118 4684
rect 12900 4681 12928 4712
rect 14538 4700 14544 4712
rect 14596 4700 14602 4752
rect 14998 4700 15004 4752
rect 15056 4740 15062 4752
rect 16120 4740 16148 4771
rect 16194 4768 16200 4780
rect 16252 4768 16258 4820
rect 17206 4808 17212 4820
rect 17167 4780 17212 4808
rect 17206 4768 17212 4780
rect 17264 4768 17270 4820
rect 18310 4808 18316 4820
rect 18271 4780 18316 4808
rect 18310 4768 18316 4780
rect 18368 4768 18374 4820
rect 18954 4808 18960 4820
rect 18420 4780 18960 4808
rect 15056 4712 16148 4740
rect 17025 4743 17083 4749
rect 15056 4700 15062 4712
rect 17025 4709 17037 4743
rect 17071 4740 17083 4743
rect 17482 4740 17488 4752
rect 17071 4712 17488 4740
rect 17071 4709 17083 4712
rect 17025 4703 17083 4709
rect 17482 4700 17488 4712
rect 17540 4700 17546 4752
rect 17666 4740 17672 4752
rect 17579 4712 17672 4740
rect 17666 4700 17672 4712
rect 17724 4740 17730 4752
rect 18420 4740 18448 4780
rect 18954 4768 18960 4780
rect 19012 4808 19018 4820
rect 19141 4811 19199 4817
rect 19141 4808 19153 4811
rect 19012 4780 19153 4808
rect 19012 4768 19018 4780
rect 19141 4777 19153 4780
rect 19187 4808 19199 4811
rect 19877 4811 19935 4817
rect 19187 4780 19368 4808
rect 19187 4777 19199 4780
rect 19141 4771 19199 4777
rect 17724 4712 18448 4740
rect 17724 4700 17730 4712
rect 18586 4700 18592 4752
rect 18644 4740 18650 4752
rect 19230 4740 19236 4752
rect 18644 4712 19236 4740
rect 18644 4700 18650 4712
rect 19230 4700 19236 4712
rect 19288 4700 19294 4752
rect 19340 4740 19368 4780
rect 19877 4777 19889 4811
rect 19923 4808 19935 4811
rect 20334 4808 20340 4820
rect 19923 4780 20340 4808
rect 19923 4777 19935 4780
rect 19877 4771 19935 4777
rect 20334 4768 20340 4780
rect 20392 4768 20398 4820
rect 22082 4808 22088 4820
rect 22043 4780 22088 4808
rect 22082 4768 22088 4780
rect 22140 4768 22146 4820
rect 23186 4808 23192 4820
rect 23147 4780 23192 4808
rect 23186 4768 23192 4780
rect 23244 4768 23250 4820
rect 23370 4768 23376 4820
rect 23428 4808 23434 4820
rect 23557 4811 23615 4817
rect 23557 4808 23569 4811
rect 23428 4780 23569 4808
rect 23428 4768 23434 4780
rect 23557 4777 23569 4780
rect 23603 4777 23615 4811
rect 23557 4771 23615 4777
rect 24293 4811 24351 4817
rect 24293 4777 24305 4811
rect 24339 4808 24351 4811
rect 24658 4808 24664 4820
rect 24339 4780 24664 4808
rect 24339 4777 24351 4780
rect 24293 4771 24351 4777
rect 24658 4768 24664 4780
rect 24716 4768 24722 4820
rect 19966 4740 19972 4752
rect 19340 4712 19972 4740
rect 19966 4700 19972 4712
rect 20024 4700 20030 4752
rect 22266 4700 22272 4752
rect 22324 4740 22330 4752
rect 25026 4740 25032 4752
rect 22324 4712 25032 4740
rect 22324 4700 22330 4712
rect 25026 4700 25032 4712
rect 25084 4700 25090 4752
rect 12885 4675 12943 4681
rect 12885 4672 12897 4675
rect 12112 4644 12897 4672
rect 12112 4632 12118 4644
rect 12885 4641 12897 4644
rect 12931 4641 12943 4675
rect 12885 4635 12943 4641
rect 13526 4632 13532 4684
rect 13584 4672 13590 4684
rect 13713 4675 13771 4681
rect 13713 4672 13725 4675
rect 13584 4644 13725 4672
rect 13584 4632 13590 4644
rect 13713 4641 13725 4644
rect 13759 4641 13771 4675
rect 13713 4635 13771 4641
rect 14817 4675 14875 4681
rect 14817 4641 14829 4675
rect 14863 4672 14875 4675
rect 16013 4675 16071 4681
rect 16013 4672 16025 4675
rect 14863 4644 16025 4672
rect 14863 4641 14875 4644
rect 14817 4635 14875 4641
rect 16013 4641 16025 4644
rect 16059 4672 16071 4675
rect 16378 4672 16384 4684
rect 16059 4644 16384 4672
rect 16059 4641 16071 4644
rect 16013 4635 16071 4641
rect 16378 4632 16384 4644
rect 16436 4632 16442 4684
rect 17114 4632 17120 4684
rect 17172 4672 17178 4684
rect 17577 4675 17635 4681
rect 17577 4672 17589 4675
rect 17172 4644 17589 4672
rect 17172 4632 17178 4644
rect 17577 4641 17589 4644
rect 17623 4641 17635 4675
rect 19248 4672 19276 4700
rect 21990 4672 21996 4684
rect 19248 4644 19368 4672
rect 21951 4644 21996 4672
rect 17577 4635 17635 4641
rect 8282 4604 8288 4616
rect 8243 4576 8288 4604
rect 8282 4564 8288 4576
rect 8340 4564 8346 4616
rect 10122 4604 10128 4616
rect 10083 4576 10128 4604
rect 10122 4564 10128 4576
rect 10180 4564 10186 4616
rect 13802 4604 13808 4616
rect 13763 4576 13808 4604
rect 13802 4564 13808 4576
rect 13860 4564 13866 4616
rect 13989 4607 14047 4613
rect 13989 4573 14001 4607
rect 14035 4604 14047 4607
rect 14078 4604 14084 4616
rect 14035 4576 14084 4604
rect 14035 4573 14047 4576
rect 13989 4567 14047 4573
rect 8837 4539 8895 4545
rect 8837 4505 8849 4539
rect 8883 4536 8895 4539
rect 9294 4536 9300 4548
rect 8883 4508 9300 4536
rect 8883 4505 8895 4508
rect 8837 4499 8895 4505
rect 9294 4496 9300 4508
rect 9352 4496 9358 4548
rect 12241 4539 12299 4545
rect 12241 4505 12253 4539
rect 12287 4536 12299 4539
rect 12790 4536 12796 4548
rect 12287 4508 12796 4536
rect 12287 4505 12299 4508
rect 12241 4499 12299 4505
rect 12790 4496 12796 4508
rect 12848 4496 12854 4548
rect 13253 4539 13311 4545
rect 13253 4505 13265 4539
rect 13299 4536 13311 4539
rect 13618 4536 13624 4548
rect 13299 4508 13624 4536
rect 13299 4505 13311 4508
rect 13253 4499 13311 4505
rect 13618 4496 13624 4508
rect 13676 4536 13682 4548
rect 14004 4536 14032 4567
rect 14078 4564 14084 4576
rect 14136 4564 14142 4616
rect 16289 4607 16347 4613
rect 16289 4573 16301 4607
rect 16335 4604 16347 4607
rect 16562 4604 16568 4616
rect 16335 4576 16568 4604
rect 16335 4573 16347 4576
rect 16289 4567 16347 4573
rect 16562 4564 16568 4576
rect 16620 4564 16626 4616
rect 17482 4564 17488 4616
rect 17540 4604 17546 4616
rect 17761 4607 17819 4613
rect 17761 4604 17773 4607
rect 17540 4576 17773 4604
rect 17540 4564 17546 4576
rect 17761 4573 17773 4576
rect 17807 4573 17819 4607
rect 19138 4604 19144 4616
rect 17761 4567 17819 4573
rect 17960 4576 19144 4604
rect 13676 4508 14032 4536
rect 13676 4496 13682 4508
rect 16470 4496 16476 4548
rect 16528 4536 16534 4548
rect 16749 4539 16807 4545
rect 16749 4536 16761 4539
rect 16528 4508 16761 4536
rect 16528 4496 16534 4508
rect 16749 4505 16761 4508
rect 16795 4536 16807 4539
rect 17960 4536 17988 4576
rect 19138 4564 19144 4576
rect 19196 4604 19202 4616
rect 19340 4613 19368 4644
rect 21990 4632 21996 4644
rect 22048 4632 22054 4684
rect 24750 4672 24756 4684
rect 24711 4644 24756 4672
rect 24750 4632 24756 4644
rect 24808 4632 24814 4684
rect 19233 4607 19291 4613
rect 19233 4604 19245 4607
rect 19196 4576 19245 4604
rect 19196 4564 19202 4576
rect 19233 4573 19245 4576
rect 19279 4573 19291 4607
rect 19233 4567 19291 4573
rect 19325 4607 19383 4613
rect 19325 4573 19337 4607
rect 19371 4573 19383 4607
rect 20610 4604 20616 4616
rect 20571 4576 20616 4604
rect 19325 4567 19383 4573
rect 20610 4564 20616 4576
rect 20668 4564 20674 4616
rect 22266 4604 22272 4616
rect 22227 4576 22272 4604
rect 22266 4564 22272 4576
rect 22324 4564 22330 4616
rect 23649 4607 23707 4613
rect 23649 4573 23661 4607
rect 23695 4573 23707 4607
rect 23649 4567 23707 4573
rect 16795 4508 17988 4536
rect 16795 4505 16807 4508
rect 16749 4499 16807 4505
rect 19046 4496 19052 4548
rect 19104 4536 19110 4548
rect 20153 4539 20211 4545
rect 20153 4536 20165 4539
rect 19104 4508 20165 4536
rect 19104 4496 19110 4508
rect 20153 4505 20165 4508
rect 20199 4505 20211 4539
rect 20153 4499 20211 4505
rect 21625 4539 21683 4545
rect 21625 4505 21637 4539
rect 21671 4536 21683 4539
rect 23005 4539 23063 4545
rect 23005 4536 23017 4539
rect 21671 4508 23017 4536
rect 21671 4505 21683 4508
rect 21625 4499 21683 4505
rect 23005 4505 23017 4508
rect 23051 4536 23063 4539
rect 23664 4536 23692 4567
rect 23738 4564 23744 4616
rect 23796 4604 23802 4616
rect 23796 4576 23841 4604
rect 23796 4564 23802 4576
rect 24937 4539 24995 4545
rect 24937 4536 24949 4539
rect 23051 4508 23692 4536
rect 23725 4508 24949 4536
rect 23051 4505 23063 4508
rect 23005 4499 23063 4505
rect 9205 4471 9263 4477
rect 9205 4437 9217 4471
rect 9251 4468 9263 4471
rect 9662 4468 9668 4480
rect 9251 4440 9668 4468
rect 9251 4437 9263 4440
rect 9205 4431 9263 4437
rect 9662 4428 9668 4440
rect 9720 4428 9726 4480
rect 12606 4468 12612 4480
rect 12567 4440 12612 4468
rect 12606 4428 12612 4440
rect 12664 4428 12670 4480
rect 12698 4428 12704 4480
rect 12756 4468 12762 4480
rect 18586 4468 18592 4480
rect 12756 4440 12801 4468
rect 18547 4440 18592 4468
rect 12756 4428 12762 4440
rect 18586 4428 18592 4440
rect 18644 4428 18650 4480
rect 18770 4468 18776 4480
rect 18731 4440 18776 4468
rect 18770 4428 18776 4440
rect 18828 4428 18834 4480
rect 21257 4471 21315 4477
rect 21257 4437 21269 4471
rect 21303 4468 21315 4471
rect 21530 4468 21536 4480
rect 21303 4440 21536 4468
rect 21303 4437 21315 4440
rect 21257 4431 21315 4437
rect 21530 4428 21536 4440
rect 21588 4428 21594 4480
rect 22634 4468 22640 4480
rect 22595 4440 22640 4468
rect 22634 4428 22640 4440
rect 22692 4468 22698 4480
rect 22910 4468 22916 4480
rect 22692 4440 22916 4468
rect 22692 4428 22698 4440
rect 22910 4428 22916 4440
rect 22968 4428 22974 4480
rect 23186 4428 23192 4480
rect 23244 4468 23250 4480
rect 23725 4468 23753 4508
rect 24937 4505 24949 4508
rect 24983 4505 24995 4539
rect 24937 4499 24995 4505
rect 24658 4468 24664 4480
rect 23244 4440 23753 4468
rect 24619 4440 24664 4468
rect 23244 4428 23250 4440
rect 24658 4428 24664 4440
rect 24716 4428 24722 4480
rect 816 4378 26576 4400
rect 816 4326 5360 4378
rect 5412 4326 5424 4378
rect 5476 4326 5488 4378
rect 5540 4326 5552 4378
rect 5604 4326 14694 4378
rect 14746 4326 14758 4378
rect 14810 4326 14822 4378
rect 14874 4326 14886 4378
rect 14938 4326 24027 4378
rect 24079 4326 24091 4378
rect 24143 4326 24155 4378
rect 24207 4326 24219 4378
rect 24271 4326 26576 4378
rect 816 4304 26576 4326
rect 14078 4224 14084 4276
rect 14136 4264 14142 4276
rect 15277 4267 15335 4273
rect 15277 4264 15289 4267
rect 14136 4236 15289 4264
rect 14136 4224 14142 4236
rect 15277 4233 15289 4236
rect 15323 4233 15335 4267
rect 15277 4227 15335 4233
rect 15921 4267 15979 4273
rect 15921 4233 15933 4267
rect 15967 4264 15979 4267
rect 16562 4264 16568 4276
rect 15967 4236 16568 4264
rect 15967 4233 15979 4236
rect 15921 4227 15979 4233
rect 10125 4199 10183 4205
rect 10125 4196 10137 4199
rect 9404 4168 10137 4196
rect 7638 4088 7644 4140
rect 7696 4128 7702 4140
rect 8101 4131 8159 4137
rect 8101 4128 8113 4131
rect 7696 4100 8113 4128
rect 7696 4088 7702 4100
rect 8101 4097 8113 4100
rect 8147 4128 8159 4131
rect 9404 4128 9432 4168
rect 10125 4165 10137 4168
rect 10171 4196 10183 4199
rect 10674 4196 10680 4208
rect 10171 4168 10680 4196
rect 10171 4165 10183 4168
rect 10125 4159 10183 4165
rect 10674 4156 10680 4168
rect 10732 4156 10738 4208
rect 9662 4128 9668 4140
rect 8147 4100 9432 4128
rect 9623 4100 9668 4128
rect 8147 4097 8159 4100
rect 8101 4091 8159 4097
rect 9662 4088 9668 4100
rect 9720 4088 9726 4140
rect 11594 4128 11600 4140
rect 10968 4100 11600 4128
rect 7089 4063 7147 4069
rect 7089 4029 7101 4063
rect 7135 4060 7147 4063
rect 7135 4032 8052 4060
rect 7135 4029 7147 4032
rect 7089 4023 7147 4029
rect 8024 4001 8052 4032
rect 8926 4020 8932 4072
rect 8984 4060 8990 4072
rect 10968 4069 10996 4100
rect 11594 4088 11600 4100
rect 11652 4088 11658 4140
rect 12790 4128 12796 4140
rect 12751 4100 12796 4128
rect 12790 4088 12796 4100
rect 12848 4088 12854 4140
rect 9481 4063 9539 4069
rect 9481 4060 9493 4063
rect 8984 4032 9493 4060
rect 8984 4020 8990 4032
rect 9481 4029 9493 4032
rect 9527 4029 9539 4063
rect 9481 4023 9539 4029
rect 10953 4063 11011 4069
rect 10953 4029 10965 4063
rect 10999 4029 11011 4063
rect 11870 4060 11876 4072
rect 11831 4032 11876 4060
rect 10953 4023 11011 4029
rect 11870 4020 11876 4032
rect 11928 4060 11934 4072
rect 12517 4063 12575 4069
rect 12517 4060 12529 4063
rect 11928 4032 12529 4060
rect 11928 4020 11934 4032
rect 12517 4029 12529 4032
rect 12563 4029 12575 4063
rect 12517 4023 12575 4029
rect 12698 4020 12704 4072
rect 12756 4060 12762 4072
rect 13894 4060 13900 4072
rect 12756 4032 13900 4060
rect 12756 4020 12762 4032
rect 13894 4020 13900 4032
rect 13952 4020 13958 4072
rect 13986 4020 13992 4072
rect 14044 4060 14050 4072
rect 14164 4063 14222 4069
rect 14164 4060 14176 4063
rect 14044 4032 14176 4060
rect 14044 4020 14050 4032
rect 14164 4029 14176 4032
rect 14210 4060 14222 4063
rect 15936 4060 15964 4227
rect 16562 4224 16568 4236
rect 16620 4224 16626 4276
rect 21990 4224 21996 4276
rect 22048 4264 22054 4276
rect 22177 4267 22235 4273
rect 22177 4264 22189 4267
rect 22048 4236 22189 4264
rect 22048 4224 22054 4236
rect 22177 4233 22189 4236
rect 22223 4233 22235 4267
rect 22177 4227 22235 4233
rect 23189 4267 23247 4273
rect 23189 4233 23201 4267
rect 23235 4264 23247 4267
rect 23370 4264 23376 4276
rect 23235 4236 23376 4264
rect 23235 4233 23247 4236
rect 23189 4227 23247 4233
rect 23370 4224 23376 4236
rect 23428 4224 23434 4276
rect 23922 4264 23928 4276
rect 23883 4236 23928 4264
rect 23922 4224 23928 4236
rect 23980 4224 23986 4276
rect 24750 4224 24756 4276
rect 24808 4264 24814 4276
rect 24937 4267 24995 4273
rect 24937 4264 24949 4267
rect 24808 4236 24949 4264
rect 24808 4224 24814 4236
rect 24937 4233 24949 4236
rect 24983 4233 24995 4267
rect 24937 4227 24995 4233
rect 20334 4196 20340 4208
rect 20260 4168 20340 4196
rect 16286 4128 16292 4140
rect 16247 4100 16292 4128
rect 16286 4088 16292 4100
rect 16344 4128 16350 4140
rect 16344 4100 16424 4128
rect 16344 4088 16350 4100
rect 16396 4069 16424 4100
rect 17298 4088 17304 4140
rect 17356 4128 17362 4140
rect 18313 4131 18371 4137
rect 18313 4128 18325 4131
rect 17356 4100 18325 4128
rect 17356 4088 17362 4100
rect 18313 4097 18325 4100
rect 18359 4128 18371 4131
rect 18586 4128 18592 4140
rect 18359 4100 18592 4128
rect 18359 4097 18371 4100
rect 18313 4091 18371 4097
rect 18586 4088 18592 4100
rect 18644 4088 18650 4140
rect 18865 4131 18923 4137
rect 18865 4097 18877 4131
rect 18911 4128 18923 4131
rect 18954 4128 18960 4140
rect 18911 4100 18960 4128
rect 18911 4097 18923 4100
rect 18865 4091 18923 4097
rect 18954 4088 18960 4100
rect 19012 4088 19018 4140
rect 20260 4137 20288 4168
rect 20334 4156 20340 4168
rect 20392 4156 20398 4208
rect 22266 4156 22272 4208
rect 22324 4196 22330 4208
rect 22637 4199 22695 4205
rect 22637 4196 22649 4199
rect 22324 4168 22649 4196
rect 22324 4156 22330 4168
rect 22637 4165 22649 4168
rect 22683 4196 22695 4199
rect 23094 4196 23100 4208
rect 22683 4168 23100 4196
rect 22683 4165 22695 4168
rect 22637 4159 22695 4165
rect 23094 4156 23100 4168
rect 23152 4196 23158 4208
rect 24658 4196 24664 4208
rect 23152 4168 24664 4196
rect 23152 4156 23158 4168
rect 20245 4131 20303 4137
rect 20245 4097 20257 4131
rect 20291 4097 20303 4131
rect 20702 4128 20708 4140
rect 20615 4100 20708 4128
rect 20245 4091 20303 4097
rect 20702 4088 20708 4100
rect 20760 4128 20766 4140
rect 21717 4131 21775 4137
rect 21717 4128 21729 4131
rect 20760 4100 21729 4128
rect 20760 4088 20766 4100
rect 21717 4097 21729 4100
rect 21763 4097 21775 4131
rect 21717 4091 21775 4097
rect 23278 4088 23284 4140
rect 23336 4128 23342 4140
rect 24584 4137 24612 4168
rect 24658 4156 24664 4168
rect 24716 4156 24722 4208
rect 23741 4131 23799 4137
rect 23741 4128 23753 4131
rect 23336 4100 23753 4128
rect 23336 4088 23342 4100
rect 23741 4097 23753 4100
rect 23787 4128 23799 4131
rect 24569 4131 24627 4137
rect 23787 4100 24336 4128
rect 23787 4097 23799 4100
rect 23741 4091 23799 4097
rect 14210 4032 15964 4060
rect 16381 4063 16439 4069
rect 14210 4029 14222 4032
rect 14164 4023 14222 4029
rect 16381 4029 16393 4063
rect 16427 4029 16439 4063
rect 18221 4063 18279 4069
rect 18221 4060 18233 4063
rect 16381 4023 16439 4029
rect 17500 4032 18233 4060
rect 6537 3995 6595 4001
rect 6537 3961 6549 3995
rect 6583 3992 6595 3995
rect 7365 3995 7423 4001
rect 7365 3992 7377 3995
rect 6583 3964 7377 3992
rect 6583 3961 6595 3964
rect 6537 3955 6595 3961
rect 7365 3961 7377 3964
rect 7411 3992 7423 3995
rect 7917 3995 7975 4001
rect 7917 3992 7929 3995
rect 7411 3964 7929 3992
rect 7411 3961 7423 3964
rect 7365 3955 7423 3961
rect 7917 3961 7929 3964
rect 7963 3961 7975 3995
rect 7917 3955 7975 3961
rect 8009 3995 8067 4001
rect 8009 3961 8021 3995
rect 8055 3992 8067 3995
rect 8055 3964 9156 3992
rect 8055 3961 8067 3964
rect 8009 3955 8067 3961
rect 7546 3924 7552 3936
rect 7507 3896 7552 3924
rect 7546 3884 7552 3896
rect 7604 3884 7610 3936
rect 8650 3924 8656 3936
rect 8611 3896 8656 3924
rect 8650 3884 8656 3896
rect 8708 3884 8714 3936
rect 8926 3924 8932 3936
rect 8887 3896 8932 3924
rect 8926 3884 8932 3896
rect 8984 3884 8990 3936
rect 9128 3933 9156 3964
rect 9386 3952 9392 4004
rect 9444 3992 9450 4004
rect 10122 3992 10128 4004
rect 9444 3964 10128 3992
rect 9444 3952 9450 3964
rect 10122 3952 10128 3964
rect 10180 3992 10186 4004
rect 10769 3995 10827 4001
rect 10769 3992 10781 3995
rect 10180 3964 10781 3992
rect 10180 3952 10186 3964
rect 10769 3961 10781 3964
rect 10815 3992 10827 3995
rect 11318 3992 11324 4004
rect 10815 3964 11324 3992
rect 10815 3961 10827 3964
rect 10769 3955 10827 3961
rect 11318 3952 11324 3964
rect 11376 3952 11382 4004
rect 17500 3936 17528 4032
rect 18221 4029 18233 4032
rect 18267 4029 18279 4063
rect 18221 4023 18279 4029
rect 20886 4020 20892 4072
rect 20944 4060 20950 4072
rect 24308 4069 24336 4100
rect 24569 4097 24581 4131
rect 24615 4097 24627 4131
rect 24569 4091 24627 4097
rect 20981 4063 21039 4069
rect 20981 4060 20993 4063
rect 20944 4032 20993 4060
rect 20944 4020 20950 4032
rect 20981 4029 20993 4032
rect 21027 4029 21039 4063
rect 20981 4023 21039 4029
rect 24293 4063 24351 4069
rect 24293 4029 24305 4063
rect 24339 4060 24351 4063
rect 24474 4060 24480 4072
rect 24339 4032 24480 4060
rect 24339 4029 24351 4032
rect 24293 4023 24351 4029
rect 18126 3992 18132 4004
rect 18087 3964 18132 3992
rect 18126 3952 18132 3964
rect 18184 3952 18190 4004
rect 19230 3952 19236 4004
rect 19288 3992 19294 4004
rect 19509 3995 19567 4001
rect 19509 3992 19521 3995
rect 19288 3964 19521 3992
rect 19288 3952 19294 3964
rect 19509 3961 19521 3964
rect 19555 3992 19567 3995
rect 20996 3992 21024 4023
rect 24474 4020 24480 4032
rect 24532 4020 24538 4072
rect 21625 3995 21683 4001
rect 21625 3992 21637 3995
rect 19555 3964 20104 3992
rect 20996 3964 21637 3992
rect 19555 3961 19567 3964
rect 19509 3955 19567 3961
rect 20076 3936 20104 3964
rect 21625 3961 21637 3964
rect 21671 3992 21683 3995
rect 21714 3992 21720 4004
rect 21671 3964 21720 3992
rect 21671 3961 21683 3964
rect 21625 3955 21683 3961
rect 21714 3952 21720 3964
rect 21772 3952 21778 4004
rect 24385 3995 24443 4001
rect 24385 3961 24397 3995
rect 24431 3992 24443 3995
rect 24566 3992 24572 4004
rect 24431 3964 24572 3992
rect 24431 3961 24443 3964
rect 24385 3955 24443 3961
rect 24566 3952 24572 3964
rect 24624 3952 24630 4004
rect 9113 3927 9171 3933
rect 9113 3893 9125 3927
rect 9159 3893 9171 3927
rect 9113 3887 9171 3893
rect 9294 3884 9300 3936
rect 9352 3924 9358 3936
rect 9570 3924 9576 3936
rect 9352 3896 9576 3924
rect 9352 3884 9358 3896
rect 9570 3884 9576 3896
rect 9628 3884 9634 3936
rect 11134 3924 11140 3936
rect 11095 3896 11140 3924
rect 11134 3884 11140 3896
rect 11192 3884 11198 3936
rect 12146 3884 12152 3936
rect 12204 3924 12210 3936
rect 12606 3924 12612 3936
rect 12204 3896 12249 3924
rect 12567 3896 12612 3924
rect 12204 3884 12210 3896
rect 12606 3884 12612 3896
rect 12664 3884 12670 3936
rect 13342 3924 13348 3936
rect 13303 3896 13348 3924
rect 13342 3884 13348 3896
rect 13400 3884 13406 3936
rect 13802 3924 13808 3936
rect 13715 3896 13808 3924
rect 13802 3884 13808 3896
rect 13860 3924 13866 3936
rect 15458 3924 15464 3936
rect 13860 3896 15464 3924
rect 13860 3884 13866 3896
rect 15458 3884 15464 3896
rect 15516 3884 15522 3936
rect 16194 3884 16200 3936
rect 16252 3924 16258 3936
rect 16565 3927 16623 3933
rect 16565 3924 16577 3927
rect 16252 3896 16577 3924
rect 16252 3884 16258 3896
rect 16565 3893 16577 3896
rect 16611 3893 16623 3927
rect 17114 3924 17120 3936
rect 17075 3896 17120 3924
rect 16565 3887 16623 3893
rect 17114 3884 17120 3896
rect 17172 3884 17178 3936
rect 17482 3924 17488 3936
rect 17443 3896 17488 3924
rect 17482 3884 17488 3896
rect 17540 3884 17546 3936
rect 17758 3924 17764 3936
rect 17719 3896 17764 3924
rect 17758 3884 17764 3896
rect 17816 3884 17822 3936
rect 19601 3927 19659 3933
rect 19601 3893 19613 3927
rect 19647 3924 19659 3927
rect 19782 3924 19788 3936
rect 19647 3896 19788 3924
rect 19647 3893 19659 3896
rect 19601 3887 19659 3893
rect 19782 3884 19788 3896
rect 19840 3884 19846 3936
rect 19966 3924 19972 3936
rect 19927 3896 19972 3924
rect 19966 3884 19972 3896
rect 20024 3884 20030 3936
rect 20058 3884 20064 3936
rect 20116 3924 20122 3936
rect 21162 3924 21168 3936
rect 20116 3896 20161 3924
rect 21123 3896 21168 3924
rect 20116 3884 20122 3896
rect 21162 3884 21168 3896
rect 21220 3884 21226 3936
rect 21530 3924 21536 3936
rect 21491 3896 21536 3924
rect 21530 3884 21536 3896
rect 21588 3884 21594 3936
rect 816 3834 26576 3856
rect 816 3782 10027 3834
rect 10079 3782 10091 3834
rect 10143 3782 10155 3834
rect 10207 3782 10219 3834
rect 10271 3782 19360 3834
rect 19412 3782 19424 3834
rect 19476 3782 19488 3834
rect 19540 3782 19552 3834
rect 19604 3782 26576 3834
rect 816 3760 26576 3782
rect 7638 3720 7644 3732
rect 7599 3692 7644 3720
rect 7638 3680 7644 3692
rect 7696 3680 7702 3732
rect 10674 3680 10680 3732
rect 10732 3720 10738 3732
rect 10769 3723 10827 3729
rect 10769 3720 10781 3723
rect 10732 3692 10781 3720
rect 10732 3680 10738 3692
rect 10769 3689 10781 3692
rect 10815 3689 10827 3723
rect 11318 3720 11324 3732
rect 11279 3692 11324 3720
rect 10769 3683 10827 3689
rect 11318 3680 11324 3692
rect 11376 3680 11382 3732
rect 12790 3680 12796 3732
rect 12848 3720 12854 3732
rect 13253 3723 13311 3729
rect 13253 3720 13265 3723
rect 12848 3692 13265 3720
rect 12848 3680 12854 3692
rect 13253 3689 13265 3692
rect 13299 3689 13311 3723
rect 13986 3720 13992 3732
rect 13947 3692 13992 3720
rect 13253 3683 13311 3689
rect 13986 3680 13992 3692
rect 14044 3680 14050 3732
rect 14357 3723 14415 3729
rect 14357 3689 14369 3723
rect 14403 3720 14415 3723
rect 14538 3720 14544 3732
rect 14403 3692 14544 3720
rect 14403 3689 14415 3692
rect 14357 3683 14415 3689
rect 14538 3680 14544 3692
rect 14596 3680 14602 3732
rect 14814 3720 14820 3732
rect 14775 3692 14820 3720
rect 14814 3680 14820 3692
rect 14872 3680 14878 3732
rect 16010 3720 16016 3732
rect 15971 3692 16016 3720
rect 16010 3680 16016 3692
rect 16068 3680 16074 3732
rect 16378 3680 16384 3732
rect 16436 3720 16442 3732
rect 16565 3723 16623 3729
rect 16565 3720 16577 3723
rect 16436 3692 16577 3720
rect 16436 3680 16442 3692
rect 16565 3689 16577 3692
rect 16611 3689 16623 3723
rect 17022 3720 17028 3732
rect 16983 3692 17028 3720
rect 16565 3683 16623 3689
rect 17022 3680 17028 3692
rect 17080 3680 17086 3732
rect 17666 3720 17672 3732
rect 17627 3692 17672 3720
rect 17666 3680 17672 3692
rect 17724 3680 17730 3732
rect 18129 3723 18187 3729
rect 18129 3689 18141 3723
rect 18175 3720 18187 3723
rect 18218 3720 18224 3732
rect 18175 3692 18224 3720
rect 18175 3689 18187 3692
rect 18129 3683 18187 3689
rect 18218 3680 18224 3692
rect 18276 3680 18282 3732
rect 18589 3723 18647 3729
rect 18589 3689 18601 3723
rect 18635 3720 18647 3723
rect 18770 3720 18776 3732
rect 18635 3692 18776 3720
rect 18635 3689 18647 3692
rect 18589 3683 18647 3689
rect 18770 3680 18776 3692
rect 18828 3720 18834 3732
rect 19969 3723 20027 3729
rect 19969 3720 19981 3723
rect 18828 3692 19981 3720
rect 18828 3680 18834 3692
rect 19969 3689 19981 3692
rect 20015 3689 20027 3723
rect 19969 3683 20027 3689
rect 20429 3723 20487 3729
rect 20429 3689 20441 3723
rect 20475 3720 20487 3723
rect 21162 3720 21168 3732
rect 20475 3692 21168 3720
rect 20475 3689 20487 3692
rect 20429 3683 20487 3689
rect 21162 3680 21168 3692
rect 21220 3680 21226 3732
rect 21901 3723 21959 3729
rect 21901 3689 21913 3723
rect 21947 3720 21959 3723
rect 22082 3720 22088 3732
rect 21947 3692 22088 3720
rect 21947 3689 21959 3692
rect 21901 3683 21959 3689
rect 22082 3680 22088 3692
rect 22140 3680 22146 3732
rect 23189 3723 23247 3729
rect 23189 3689 23201 3723
rect 23235 3720 23247 3723
rect 23738 3720 23744 3732
rect 23235 3692 23744 3720
rect 23235 3689 23247 3692
rect 23189 3683 23247 3689
rect 23738 3680 23744 3692
rect 23796 3680 23802 3732
rect 9294 3612 9300 3664
rect 9352 3652 9358 3664
rect 9662 3661 9668 3664
rect 9656 3652 9668 3661
rect 9352 3624 9668 3652
rect 9352 3612 9358 3624
rect 9656 3615 9668 3624
rect 9662 3612 9668 3615
rect 9720 3612 9726 3664
rect 8193 3587 8251 3593
rect 8193 3553 8205 3587
rect 8239 3584 8251 3587
rect 8466 3584 8472 3596
rect 8239 3556 8472 3584
rect 8239 3553 8251 3556
rect 8193 3547 8251 3553
rect 8466 3544 8472 3556
rect 8524 3544 8530 3596
rect 11336 3584 11364 3680
rect 16838 3612 16844 3664
rect 16896 3652 16902 3664
rect 16933 3655 16991 3661
rect 16933 3652 16945 3655
rect 16896 3624 16945 3652
rect 16896 3612 16902 3624
rect 16933 3621 16945 3624
rect 16979 3621 16991 3655
rect 16933 3615 16991 3621
rect 17758 3612 17764 3664
rect 17816 3652 17822 3664
rect 18497 3655 18555 3661
rect 18497 3652 18509 3655
rect 17816 3624 18509 3652
rect 17816 3612 17822 3624
rect 18497 3621 18509 3624
rect 18543 3652 18555 3655
rect 18954 3652 18960 3664
rect 18543 3624 18960 3652
rect 18543 3621 18555 3624
rect 18497 3615 18555 3621
rect 18954 3612 18960 3624
rect 19012 3612 19018 3664
rect 19138 3652 19144 3664
rect 19099 3624 19144 3652
rect 19138 3612 19144 3624
rect 19196 3612 19202 3664
rect 23554 3661 23560 3664
rect 23548 3652 23560 3661
rect 23515 3624 23560 3652
rect 23548 3615 23560 3624
rect 23554 3612 23560 3615
rect 23612 3612 23618 3664
rect 11873 3587 11931 3593
rect 11873 3584 11885 3587
rect 11336 3556 11885 3584
rect 11873 3553 11885 3556
rect 11919 3584 11931 3587
rect 11962 3584 11968 3596
rect 11919 3556 11968 3584
rect 11919 3553 11931 3556
rect 11873 3547 11931 3553
rect 11962 3544 11968 3556
rect 12020 3544 12026 3596
rect 12146 3593 12152 3596
rect 12140 3547 12152 3593
rect 12204 3584 12210 3596
rect 15366 3584 15372 3596
rect 12204 3556 12240 3584
rect 15327 3556 15372 3584
rect 12146 3544 12152 3547
rect 12204 3544 12210 3556
rect 15366 3544 15372 3556
rect 15424 3544 15430 3596
rect 15458 3544 15464 3596
rect 15516 3584 15522 3596
rect 16378 3584 16384 3596
rect 15516 3556 16384 3584
rect 15516 3544 15522 3556
rect 16378 3544 16384 3556
rect 16436 3544 16442 3596
rect 18037 3587 18095 3593
rect 18037 3553 18049 3587
rect 18083 3584 18095 3587
rect 18126 3584 18132 3596
rect 18083 3556 18132 3584
rect 18083 3553 18095 3556
rect 18037 3547 18095 3553
rect 18126 3544 18132 3556
rect 18184 3544 18190 3596
rect 22269 3587 22327 3593
rect 22269 3553 22281 3587
rect 22315 3584 22327 3587
rect 22634 3584 22640 3596
rect 22315 3556 22640 3584
rect 22315 3553 22327 3556
rect 22269 3547 22327 3553
rect 22634 3544 22640 3556
rect 22692 3584 22698 3596
rect 23281 3587 23339 3593
rect 23281 3584 23293 3587
rect 22692 3556 23293 3584
rect 22692 3544 22698 3556
rect 23281 3553 23293 3556
rect 23327 3584 23339 3587
rect 24566 3584 24572 3596
rect 23327 3556 24572 3584
rect 23327 3553 23339 3556
rect 23281 3547 23339 3553
rect 24566 3544 24572 3556
rect 24624 3544 24630 3596
rect 9386 3516 9392 3528
rect 8760 3488 9392 3516
rect 8377 3383 8435 3389
rect 8377 3349 8389 3383
rect 8423 3380 8435 3383
rect 8558 3380 8564 3392
rect 8423 3352 8564 3380
rect 8423 3349 8435 3352
rect 8377 3343 8435 3349
rect 8558 3340 8564 3352
rect 8616 3340 8622 3392
rect 8650 3340 8656 3392
rect 8708 3380 8714 3392
rect 8760 3389 8788 3488
rect 9386 3476 9392 3488
rect 9444 3516 9450 3528
rect 15550 3516 15556 3528
rect 9444 3488 9537 3516
rect 15511 3488 15556 3516
rect 9444 3476 9450 3488
rect 15550 3476 15556 3488
rect 15608 3476 15614 3528
rect 17206 3516 17212 3528
rect 17167 3488 17212 3516
rect 17206 3476 17212 3488
rect 17264 3476 17270 3528
rect 18678 3516 18684 3528
rect 18639 3488 18684 3516
rect 18678 3476 18684 3488
rect 18736 3476 18742 3528
rect 21254 3516 21260 3528
rect 21215 3488 21260 3516
rect 21254 3476 21260 3488
rect 21312 3476 21318 3528
rect 21346 3476 21352 3528
rect 21404 3516 21410 3528
rect 21404 3488 21449 3516
rect 21404 3476 21410 3488
rect 8745 3383 8803 3389
rect 8745 3380 8757 3383
rect 8708 3352 8757 3380
rect 8708 3340 8714 3352
rect 8745 3349 8757 3352
rect 8791 3349 8803 3383
rect 8745 3343 8803 3349
rect 9205 3383 9263 3389
rect 9205 3349 9217 3383
rect 9251 3380 9263 3383
rect 9570 3380 9576 3392
rect 9251 3352 9576 3380
rect 9251 3349 9263 3352
rect 9205 3343 9263 3349
rect 9570 3340 9576 3352
rect 9628 3380 9634 3392
rect 10490 3380 10496 3392
rect 9628 3352 10496 3380
rect 9628 3340 9634 3352
rect 10490 3340 10496 3352
rect 10548 3340 10554 3392
rect 11781 3383 11839 3389
rect 11781 3349 11793 3383
rect 11827 3380 11839 3383
rect 12882 3380 12888 3392
rect 11827 3352 12888 3380
rect 11827 3349 11839 3352
rect 11781 3343 11839 3349
rect 12882 3340 12888 3352
rect 12940 3340 12946 3392
rect 14998 3380 15004 3392
rect 14959 3352 15004 3380
rect 14998 3340 15004 3352
rect 15056 3340 15062 3392
rect 16473 3383 16531 3389
rect 16473 3349 16485 3383
rect 16519 3380 16531 3383
rect 17298 3380 17304 3392
rect 16519 3352 17304 3380
rect 16519 3349 16531 3352
rect 16473 3343 16531 3349
rect 17298 3340 17304 3352
rect 17356 3340 17362 3392
rect 19138 3340 19144 3392
rect 19196 3380 19202 3392
rect 19601 3383 19659 3389
rect 19601 3380 19613 3383
rect 19196 3352 19613 3380
rect 19196 3340 19202 3352
rect 19601 3349 19613 3352
rect 19647 3380 19659 3383
rect 19966 3380 19972 3392
rect 19647 3352 19972 3380
rect 19647 3349 19659 3352
rect 19601 3343 19659 3349
rect 19966 3340 19972 3352
rect 20024 3340 20030 3392
rect 20794 3380 20800 3392
rect 20755 3352 20800 3380
rect 20794 3340 20800 3352
rect 20852 3340 20858 3392
rect 24658 3380 24664 3392
rect 24619 3352 24664 3380
rect 24658 3340 24664 3352
rect 24716 3340 24722 3392
rect 816 3290 26576 3312
rect 816 3238 5360 3290
rect 5412 3238 5424 3290
rect 5476 3238 5488 3290
rect 5540 3238 5552 3290
rect 5604 3238 14694 3290
rect 14746 3238 14758 3290
rect 14810 3238 14822 3290
rect 14874 3238 14886 3290
rect 14938 3238 24027 3290
rect 24079 3238 24091 3290
rect 24143 3238 24155 3290
rect 24207 3238 24219 3290
rect 24271 3238 26576 3290
rect 816 3216 26576 3238
rect 7733 3179 7791 3185
rect 7733 3145 7745 3179
rect 7779 3176 7791 3179
rect 8650 3176 8656 3188
rect 7779 3148 8656 3176
rect 7779 3145 7791 3148
rect 7733 3139 7791 3145
rect 8650 3136 8656 3148
rect 8708 3136 8714 3188
rect 8834 3176 8840 3188
rect 8795 3148 8840 3176
rect 8834 3136 8840 3148
rect 8892 3136 8898 3188
rect 9662 3136 9668 3188
rect 9720 3176 9726 3188
rect 10677 3179 10735 3185
rect 10677 3176 10689 3179
rect 9720 3148 10689 3176
rect 9720 3136 9726 3148
rect 10677 3145 10689 3148
rect 10723 3145 10735 3179
rect 12422 3176 12428 3188
rect 12383 3148 12428 3176
rect 10677 3139 10735 3145
rect 12422 3136 12428 3148
rect 12480 3136 12486 3188
rect 15369 3179 15427 3185
rect 15369 3145 15381 3179
rect 15415 3176 15427 3179
rect 15550 3176 15556 3188
rect 15415 3148 15556 3176
rect 15415 3145 15427 3148
rect 15369 3139 15427 3145
rect 15550 3136 15556 3148
rect 15608 3136 15614 3188
rect 16378 3176 16384 3188
rect 16339 3148 16384 3176
rect 16378 3136 16384 3148
rect 16436 3136 16442 3188
rect 16838 3136 16844 3188
rect 16896 3176 16902 3188
rect 17393 3179 17451 3185
rect 17393 3176 17405 3179
rect 16896 3148 17405 3176
rect 16896 3136 16902 3148
rect 17393 3145 17405 3148
rect 17439 3145 17451 3179
rect 17393 3139 17451 3145
rect 18678 3136 18684 3188
rect 18736 3176 18742 3188
rect 19141 3179 19199 3185
rect 19141 3176 19153 3179
rect 18736 3148 19153 3176
rect 18736 3136 18742 3148
rect 19141 3145 19153 3148
rect 19187 3176 19199 3179
rect 19693 3179 19751 3185
rect 19693 3176 19705 3179
rect 19187 3148 19705 3176
rect 19187 3145 19199 3148
rect 19141 3139 19199 3145
rect 19693 3145 19705 3148
rect 19739 3145 19751 3179
rect 19693 3139 19751 3145
rect 21254 3136 21260 3188
rect 21312 3176 21318 3188
rect 22085 3179 22143 3185
rect 22085 3176 22097 3179
rect 21312 3148 22097 3176
rect 21312 3136 21318 3148
rect 22085 3145 22097 3148
rect 22131 3145 22143 3179
rect 23186 3176 23192 3188
rect 23147 3148 23192 3176
rect 22085 3139 22143 3145
rect 23186 3136 23192 3148
rect 23244 3136 23250 3188
rect 8101 3111 8159 3117
rect 8101 3077 8113 3111
rect 8147 3108 8159 3111
rect 8466 3108 8472 3120
rect 8147 3080 8472 3108
rect 8147 3077 8159 3080
rect 8101 3071 8159 3077
rect 8466 3068 8472 3080
rect 8524 3068 8530 3120
rect 8668 3108 8696 3136
rect 8668 3080 9156 3108
rect 8193 2975 8251 2981
rect 8193 2941 8205 2975
rect 8239 2972 8251 2975
rect 8834 2972 8840 2984
rect 8239 2944 8840 2972
rect 8239 2941 8251 2944
rect 8193 2935 8251 2941
rect 8834 2932 8840 2944
rect 8892 2932 8898 2984
rect 9128 2972 9156 3080
rect 15090 3068 15096 3120
rect 15148 3108 15154 3120
rect 16657 3111 16715 3117
rect 16657 3108 16669 3111
rect 15148 3080 16669 3108
rect 15148 3068 15154 3080
rect 16657 3077 16669 3080
rect 16703 3077 16715 3111
rect 17022 3108 17028 3120
rect 16983 3080 17028 3108
rect 16657 3071 16715 3077
rect 17022 3068 17028 3080
rect 17080 3068 17086 3120
rect 9205 3043 9263 3049
rect 9205 3009 9217 3043
rect 9251 3040 9263 3043
rect 11597 3043 11655 3049
rect 9251 3012 9432 3040
rect 9251 3009 9263 3012
rect 9205 3003 9263 3009
rect 9297 2975 9355 2981
rect 9297 2972 9309 2975
rect 9128 2944 9309 2972
rect 9297 2941 9309 2944
rect 9343 2941 9355 2975
rect 9404 2972 9432 3012
rect 11597 3009 11609 3043
rect 11643 3040 11655 3043
rect 13066 3040 13072 3052
rect 11643 3012 13072 3040
rect 11643 3009 11655 3012
rect 11597 3003 11655 3009
rect 13066 3000 13072 3012
rect 13124 3000 13130 3052
rect 13894 3000 13900 3052
rect 13952 3040 13958 3052
rect 13989 3043 14047 3049
rect 13989 3040 14001 3043
rect 13952 3012 14001 3040
rect 13952 3000 13958 3012
rect 13989 3009 14001 3012
rect 14035 3009 14047 3043
rect 13989 3003 14047 3009
rect 15366 3000 15372 3052
rect 15424 3040 15430 3052
rect 15921 3043 15979 3049
rect 15921 3040 15933 3043
rect 15424 3012 15933 3040
rect 15424 3000 15430 3012
rect 15921 3009 15933 3012
rect 15967 3009 15979 3043
rect 20242 3040 20248 3052
rect 20203 3012 20248 3040
rect 15921 3003 15979 3009
rect 20242 3000 20248 3012
rect 20300 3000 20306 3052
rect 22821 3043 22879 3049
rect 22821 3009 22833 3043
rect 22867 3040 22879 3043
rect 23554 3040 23560 3052
rect 22867 3012 23560 3040
rect 22867 3009 22879 3012
rect 22821 3003 22879 3009
rect 23554 3000 23560 3012
rect 23612 3000 23618 3052
rect 23922 3040 23928 3052
rect 23883 3012 23928 3040
rect 23922 3000 23928 3012
rect 23980 3040 23986 3052
rect 24385 3043 24443 3049
rect 24385 3040 24397 3043
rect 23980 3012 24397 3040
rect 23980 3000 23986 3012
rect 24385 3009 24397 3012
rect 24431 3040 24443 3043
rect 24658 3040 24664 3052
rect 24431 3012 24664 3040
rect 24431 3009 24443 3012
rect 24385 3003 24443 3009
rect 24658 3000 24664 3012
rect 24716 3000 24722 3052
rect 9564 2975 9622 2981
rect 9564 2972 9576 2975
rect 9404 2944 9576 2972
rect 9297 2935 9355 2941
rect 9564 2941 9576 2944
rect 9610 2972 9622 2975
rect 10398 2972 10404 2984
rect 9610 2944 10404 2972
rect 9610 2941 9622 2944
rect 9564 2935 9622 2941
rect 10398 2932 10404 2944
rect 10456 2932 10462 2984
rect 12146 2932 12152 2984
rect 12204 2972 12210 2984
rect 13437 2975 13495 2981
rect 13437 2972 13449 2975
rect 12204 2944 13449 2972
rect 12204 2932 12210 2944
rect 13437 2941 13449 2944
rect 13483 2972 13495 2975
rect 13526 2972 13532 2984
rect 13483 2944 13532 2972
rect 13483 2941 13495 2944
rect 13437 2935 13495 2941
rect 13526 2932 13532 2944
rect 13584 2932 13590 2984
rect 16010 2932 16016 2984
rect 16068 2972 16074 2984
rect 16473 2975 16531 2981
rect 16473 2972 16485 2975
rect 16068 2944 16485 2972
rect 16068 2932 16074 2944
rect 16473 2941 16485 2944
rect 16519 2941 16531 2975
rect 17758 2972 17764 2984
rect 17671 2944 17764 2972
rect 16473 2935 16531 2941
rect 17758 2932 17764 2944
rect 17816 2972 17822 2984
rect 20260 2972 20288 3000
rect 20512 2975 20570 2981
rect 20512 2972 20524 2975
rect 17816 2944 20288 2972
rect 20352 2944 20524 2972
rect 17816 2932 17822 2944
rect 7178 2904 7184 2916
rect 7139 2876 7184 2904
rect 7178 2864 7184 2876
rect 7236 2864 7242 2916
rect 11870 2904 11876 2916
rect 11831 2876 11876 2904
rect 11870 2864 11876 2876
rect 11928 2904 11934 2916
rect 12793 2907 12851 2913
rect 12793 2904 12805 2907
rect 11928 2876 12805 2904
rect 11928 2864 11934 2876
rect 12793 2873 12805 2876
rect 12839 2873 12851 2907
rect 12793 2867 12851 2873
rect 12882 2864 12888 2916
rect 12940 2904 12946 2916
rect 13897 2907 13955 2913
rect 12940 2876 12985 2904
rect 12940 2864 12946 2876
rect 13897 2873 13909 2907
rect 13943 2904 13955 2907
rect 14234 2907 14292 2913
rect 14234 2904 14246 2907
rect 13943 2876 14246 2904
rect 13943 2873 13955 2876
rect 13897 2867 13955 2873
rect 14234 2873 14246 2876
rect 14280 2904 14292 2907
rect 14538 2904 14544 2916
rect 14280 2876 14544 2904
rect 14280 2873 14292 2876
rect 14234 2867 14292 2873
rect 14538 2864 14544 2876
rect 14596 2864 14602 2916
rect 17298 2864 17304 2916
rect 17356 2904 17362 2916
rect 18006 2907 18064 2913
rect 18006 2904 18018 2907
rect 17356 2876 18018 2904
rect 17356 2864 17362 2876
rect 18006 2873 18018 2876
rect 18052 2904 18064 2907
rect 19046 2904 19052 2916
rect 18052 2876 19052 2904
rect 18052 2873 18064 2876
rect 18006 2867 18064 2873
rect 19046 2864 19052 2876
rect 19104 2864 19110 2916
rect 20153 2907 20211 2913
rect 20153 2873 20165 2907
rect 20199 2904 20211 2907
rect 20242 2904 20248 2916
rect 20199 2876 20248 2904
rect 20199 2873 20211 2876
rect 20153 2867 20211 2873
rect 20242 2864 20248 2876
rect 20300 2904 20306 2916
rect 20352 2904 20380 2944
rect 20512 2941 20524 2944
rect 20558 2972 20570 2975
rect 21346 2972 21352 2984
rect 20558 2944 21352 2972
rect 20558 2941 20570 2944
rect 20512 2935 20570 2941
rect 21346 2932 21352 2944
rect 21404 2932 21410 2984
rect 23462 2932 23468 2984
rect 23520 2972 23526 2984
rect 23741 2975 23799 2981
rect 23741 2972 23753 2975
rect 23520 2944 23753 2972
rect 23520 2932 23526 2944
rect 23741 2941 23753 2944
rect 23787 2941 23799 2975
rect 23741 2935 23799 2941
rect 20300 2876 20380 2904
rect 20300 2864 20306 2876
rect 23186 2864 23192 2916
rect 23244 2904 23250 2916
rect 23830 2904 23836 2916
rect 23244 2876 23836 2904
rect 23244 2864 23250 2876
rect 23830 2864 23836 2876
rect 23888 2864 23894 2916
rect 24566 2864 24572 2916
rect 24624 2904 24630 2916
rect 24845 2907 24903 2913
rect 24845 2904 24857 2907
rect 24624 2876 24857 2904
rect 24624 2864 24630 2876
rect 24845 2873 24857 2876
rect 24891 2904 24903 2907
rect 24891 2876 25624 2904
rect 24891 2873 24903 2876
rect 24845 2867 24903 2873
rect 8377 2839 8435 2845
rect 8377 2805 8389 2839
rect 8423 2836 8435 2839
rect 8650 2836 8656 2848
rect 8423 2808 8656 2836
rect 8423 2805 8435 2808
rect 8377 2799 8435 2805
rect 8650 2796 8656 2808
rect 8708 2796 8714 2848
rect 10398 2796 10404 2848
rect 10456 2836 10462 2848
rect 13710 2836 13716 2848
rect 10456 2808 13716 2836
rect 10456 2796 10462 2808
rect 13710 2796 13716 2808
rect 13768 2796 13774 2848
rect 21625 2839 21683 2845
rect 21625 2805 21637 2839
rect 21671 2836 21683 2839
rect 21714 2836 21720 2848
rect 21671 2808 21720 2836
rect 21671 2805 21683 2808
rect 21625 2799 21683 2805
rect 21714 2796 21720 2808
rect 21772 2796 21778 2848
rect 22085 2839 22143 2845
rect 22085 2805 22097 2839
rect 22131 2836 22143 2839
rect 22269 2839 22327 2845
rect 22269 2836 22281 2839
rect 22131 2808 22281 2836
rect 22131 2805 22143 2808
rect 22085 2799 22143 2805
rect 22269 2805 22281 2808
rect 22315 2836 22327 2839
rect 23373 2839 23431 2845
rect 23373 2836 23385 2839
rect 22315 2808 23385 2836
rect 22315 2805 22327 2808
rect 22269 2799 22327 2805
rect 23373 2805 23385 2808
rect 23419 2805 23431 2839
rect 25118 2836 25124 2848
rect 25079 2808 25124 2836
rect 23373 2799 23431 2805
rect 25118 2796 25124 2808
rect 25176 2796 25182 2848
rect 25596 2845 25624 2876
rect 25581 2839 25639 2845
rect 25581 2805 25593 2839
rect 25627 2836 25639 2839
rect 25762 2836 25768 2848
rect 25627 2808 25768 2836
rect 25627 2805 25639 2808
rect 25581 2799 25639 2805
rect 25762 2796 25768 2808
rect 25820 2836 25826 2848
rect 25857 2839 25915 2845
rect 25857 2836 25869 2839
rect 25820 2808 25869 2836
rect 25820 2796 25826 2808
rect 25857 2805 25869 2808
rect 25903 2805 25915 2839
rect 25857 2799 25915 2805
rect 816 2746 26576 2768
rect 816 2694 10027 2746
rect 10079 2694 10091 2746
rect 10143 2694 10155 2746
rect 10207 2694 10219 2746
rect 10271 2694 19360 2746
rect 19412 2694 19424 2746
rect 19476 2694 19488 2746
rect 19540 2694 19552 2746
rect 19604 2694 26576 2746
rect 816 2672 26576 2694
rect 9294 2632 9300 2644
rect 9255 2604 9300 2632
rect 9294 2592 9300 2604
rect 9352 2592 9358 2644
rect 10674 2632 10680 2644
rect 10635 2604 10680 2632
rect 10674 2592 10680 2604
rect 10732 2592 10738 2644
rect 11781 2635 11839 2641
rect 11781 2601 11793 2635
rect 11827 2632 11839 2635
rect 12054 2632 12060 2644
rect 11827 2604 12060 2632
rect 11827 2601 11839 2604
rect 11781 2595 11839 2601
rect 6997 2567 7055 2573
rect 6997 2533 7009 2567
rect 7043 2564 7055 2567
rect 10217 2567 10275 2573
rect 7043 2536 8512 2564
rect 7043 2533 7055 2536
rect 6997 2527 7055 2533
rect 7365 2499 7423 2505
rect 7365 2465 7377 2499
rect 7411 2496 7423 2499
rect 8190 2496 8196 2508
rect 7411 2468 8196 2496
rect 7411 2465 7423 2468
rect 7365 2459 7423 2465
rect 8190 2456 8196 2468
rect 8248 2456 8254 2508
rect 8484 2440 8512 2536
rect 10217 2533 10229 2567
rect 10263 2564 10275 2567
rect 10950 2564 10956 2576
rect 10263 2536 10956 2564
rect 10263 2533 10275 2536
rect 10217 2527 10275 2533
rect 10950 2524 10956 2536
rect 11008 2564 11014 2576
rect 11137 2567 11195 2573
rect 11137 2564 11149 2567
rect 11008 2536 11149 2564
rect 11008 2524 11014 2536
rect 11137 2533 11149 2536
rect 11183 2533 11195 2567
rect 11137 2527 11195 2533
rect 8929 2499 8987 2505
rect 8929 2465 8941 2499
rect 8975 2496 8987 2499
rect 9573 2499 9631 2505
rect 9573 2496 9585 2499
rect 8975 2468 9585 2496
rect 8975 2465 8987 2468
rect 8929 2459 8987 2465
rect 9573 2465 9585 2468
rect 9619 2496 9631 2499
rect 10398 2496 10404 2508
rect 9619 2468 10404 2496
rect 9619 2465 9631 2468
rect 9573 2459 9631 2465
rect 10398 2456 10404 2468
rect 10456 2456 10462 2508
rect 10490 2456 10496 2508
rect 10548 2496 10554 2508
rect 11045 2499 11103 2505
rect 11045 2496 11057 2499
rect 10548 2468 11057 2496
rect 10548 2456 10554 2468
rect 11045 2465 11057 2468
rect 11091 2465 11103 2499
rect 11045 2459 11103 2465
rect 7733 2431 7791 2437
rect 7733 2397 7745 2431
rect 7779 2428 7791 2431
rect 8282 2428 8288 2440
rect 7779 2400 8288 2428
rect 7779 2397 7791 2400
rect 7733 2391 7791 2397
rect 8282 2388 8288 2400
rect 8340 2388 8346 2440
rect 8466 2428 8472 2440
rect 8427 2400 8472 2428
rect 8466 2388 8472 2400
rect 8524 2388 8530 2440
rect 11321 2431 11379 2437
rect 11321 2397 11333 2431
rect 11367 2428 11379 2431
rect 11796 2428 11824 2595
rect 12054 2592 12060 2604
rect 12112 2592 12118 2644
rect 13526 2592 13532 2644
rect 13584 2632 13590 2644
rect 13713 2635 13771 2641
rect 13713 2632 13725 2635
rect 13584 2604 13725 2632
rect 13584 2592 13590 2604
rect 13713 2601 13725 2604
rect 13759 2601 13771 2635
rect 16562 2632 16568 2644
rect 16523 2604 16568 2632
rect 13713 2595 13771 2601
rect 16562 2592 16568 2604
rect 16620 2592 16626 2644
rect 17206 2632 17212 2644
rect 17167 2604 17212 2632
rect 17206 2592 17212 2604
rect 17264 2592 17270 2644
rect 19046 2592 19052 2644
rect 19104 2632 19110 2644
rect 19417 2635 19475 2641
rect 19417 2632 19429 2635
rect 19104 2604 19429 2632
rect 19104 2592 19110 2604
rect 19417 2601 19429 2604
rect 19463 2601 19475 2635
rect 20702 2632 20708 2644
rect 20663 2604 20708 2632
rect 19417 2595 19475 2601
rect 20702 2592 20708 2604
rect 20760 2592 20766 2644
rect 21346 2592 21352 2644
rect 21404 2632 21410 2644
rect 22269 2635 22327 2641
rect 22269 2632 22281 2635
rect 21404 2604 22281 2632
rect 21404 2592 21410 2604
rect 22269 2601 22281 2604
rect 22315 2601 22327 2635
rect 22269 2595 22327 2601
rect 23002 2592 23008 2644
rect 23060 2632 23066 2644
rect 23741 2635 23799 2641
rect 23741 2632 23753 2635
rect 23060 2604 23753 2632
rect 23060 2592 23066 2604
rect 23741 2601 23753 2604
rect 23787 2601 23799 2635
rect 24198 2632 24204 2644
rect 24159 2604 24204 2632
rect 23741 2595 23799 2601
rect 24198 2592 24204 2604
rect 24256 2632 24262 2644
rect 24753 2635 24811 2641
rect 24753 2632 24765 2635
rect 24256 2604 24765 2632
rect 24256 2592 24262 2604
rect 24753 2601 24765 2604
rect 24799 2601 24811 2635
rect 25762 2632 25768 2644
rect 25723 2604 25768 2632
rect 24753 2595 24811 2601
rect 25762 2592 25768 2604
rect 25820 2592 25826 2644
rect 12149 2567 12207 2573
rect 12149 2533 12161 2567
rect 12195 2564 12207 2567
rect 12600 2567 12658 2573
rect 12600 2564 12612 2567
rect 12195 2536 12612 2564
rect 12195 2533 12207 2536
rect 12149 2527 12207 2533
rect 12600 2533 12612 2536
rect 12646 2564 12658 2567
rect 13066 2564 13072 2576
rect 12646 2536 13072 2564
rect 12646 2533 12658 2536
rect 12600 2527 12658 2533
rect 13066 2524 13072 2536
rect 13124 2524 13130 2576
rect 14633 2567 14691 2573
rect 14633 2533 14645 2567
rect 14679 2564 14691 2567
rect 15001 2567 15059 2573
rect 15001 2564 15013 2567
rect 14679 2536 15013 2564
rect 14679 2533 14691 2536
rect 14633 2527 14691 2533
rect 15001 2533 15013 2536
rect 15047 2564 15059 2567
rect 15452 2567 15510 2573
rect 15452 2564 15464 2567
rect 15047 2536 15464 2564
rect 15047 2533 15059 2536
rect 15001 2527 15059 2533
rect 15452 2533 15464 2536
rect 15498 2564 15510 2567
rect 15550 2564 15556 2576
rect 15498 2536 15556 2564
rect 15498 2533 15510 2536
rect 15452 2527 15510 2533
rect 15550 2524 15556 2536
rect 15608 2524 15614 2576
rect 20720 2564 20748 2592
rect 21134 2567 21192 2573
rect 21134 2564 21146 2567
rect 20720 2536 21146 2564
rect 21134 2533 21146 2536
rect 21180 2533 21192 2567
rect 21134 2527 21192 2533
rect 11962 2456 11968 2508
rect 12020 2496 12026 2508
rect 12333 2499 12391 2505
rect 12333 2496 12345 2499
rect 12020 2468 12345 2496
rect 12020 2456 12026 2468
rect 12333 2465 12345 2468
rect 12379 2465 12391 2499
rect 12333 2459 12391 2465
rect 13894 2456 13900 2508
rect 13952 2496 13958 2508
rect 18310 2505 18316 2508
rect 15185 2499 15243 2505
rect 15185 2496 15197 2499
rect 13952 2468 15197 2496
rect 13952 2456 13958 2468
rect 15185 2465 15197 2468
rect 15231 2465 15243 2499
rect 15185 2459 15243 2465
rect 17853 2499 17911 2505
rect 17853 2465 17865 2499
rect 17899 2496 17911 2499
rect 18304 2496 18316 2505
rect 17899 2468 18316 2496
rect 17899 2465 17911 2468
rect 17853 2459 17911 2465
rect 18304 2459 18316 2468
rect 18310 2456 18316 2459
rect 18368 2456 18374 2508
rect 20426 2456 20432 2508
rect 20484 2496 20490 2508
rect 20889 2499 20947 2505
rect 20889 2496 20901 2499
rect 20484 2468 20901 2496
rect 20484 2456 20490 2468
rect 20889 2465 20901 2468
rect 20935 2465 20947 2499
rect 20889 2459 20947 2465
rect 21714 2456 21720 2508
rect 21772 2496 21778 2508
rect 23005 2499 23063 2505
rect 23005 2496 23017 2499
rect 21772 2468 23017 2496
rect 21772 2456 21778 2468
rect 23005 2465 23017 2468
rect 23051 2465 23063 2499
rect 24106 2496 24112 2508
rect 24067 2468 24112 2496
rect 23005 2459 23063 2465
rect 11367 2400 11824 2428
rect 11367 2397 11379 2400
rect 11321 2391 11379 2397
rect 17758 2388 17764 2440
rect 17816 2428 17822 2440
rect 18037 2431 18095 2437
rect 18037 2428 18049 2431
rect 17816 2400 18049 2428
rect 17816 2388 17822 2400
rect 18037 2397 18049 2400
rect 18083 2397 18095 2431
rect 18037 2391 18095 2397
rect 7822 2360 7828 2372
rect 7783 2332 7828 2360
rect 7822 2320 7828 2332
rect 7880 2320 7886 2372
rect 23020 2360 23048 2459
rect 24106 2456 24112 2468
rect 24164 2496 24170 2508
rect 25121 2499 25179 2505
rect 25121 2496 25133 2499
rect 24164 2468 25133 2496
rect 24164 2456 24170 2468
rect 25121 2465 25133 2468
rect 25167 2465 25179 2499
rect 25121 2459 25179 2465
rect 24293 2431 24351 2437
rect 24293 2397 24305 2431
rect 24339 2397 24351 2431
rect 24293 2391 24351 2397
rect 24308 2360 24336 2391
rect 24566 2388 24572 2440
rect 24624 2428 24630 2440
rect 25305 2431 25363 2437
rect 25305 2428 25317 2431
rect 24624 2400 25317 2428
rect 24624 2388 24630 2400
rect 25305 2397 25317 2400
rect 25351 2397 25363 2431
rect 25305 2391 25363 2397
rect 23020 2332 24336 2360
rect 9757 2295 9815 2301
rect 9757 2261 9769 2295
rect 9803 2292 9815 2295
rect 10398 2292 10404 2304
rect 9803 2264 10404 2292
rect 9803 2261 9815 2264
rect 9757 2255 9815 2261
rect 10398 2252 10404 2264
rect 10456 2252 10462 2304
rect 10490 2252 10496 2304
rect 10548 2292 10554 2304
rect 20242 2292 20248 2304
rect 10548 2264 10593 2292
rect 20203 2264 20248 2292
rect 10548 2252 10554 2264
rect 20242 2252 20248 2264
rect 20300 2252 20306 2304
rect 23462 2292 23468 2304
rect 23423 2264 23468 2292
rect 23462 2252 23468 2264
rect 23520 2252 23526 2304
rect 816 2202 26576 2224
rect 816 2150 5360 2202
rect 5412 2150 5424 2202
rect 5476 2150 5488 2202
rect 5540 2150 5552 2202
rect 5604 2150 14694 2202
rect 14746 2150 14758 2202
rect 14810 2150 14822 2202
rect 14874 2150 14886 2202
rect 14938 2150 24027 2202
rect 24079 2150 24091 2202
rect 24143 2150 24155 2202
rect 24207 2150 24219 2202
rect 24271 2150 26576 2202
rect 816 2128 26576 2150
rect 21622 1980 21628 2032
rect 21680 2020 21686 2032
rect 24014 2020 24020 2032
rect 21680 1992 24020 2020
rect 21680 1980 21686 1992
rect 24014 1980 24020 1992
rect 24072 1980 24078 2032
rect 17482 552 17488 604
rect 17540 592 17546 604
rect 18034 592 18040 604
rect 17540 564 18040 592
rect 17540 552 17546 564
rect 18034 552 18040 564
rect 18092 552 18098 604
rect 18126 552 18132 604
rect 18184 592 18190 604
rect 18586 592 18592 604
rect 18184 564 18592 592
rect 18184 552 18190 564
rect 18586 552 18592 564
rect 18644 552 18650 604
rect 22082 552 22088 604
rect 22140 592 22146 604
rect 25210 592 25216 604
rect 22140 564 25216 592
rect 22140 552 22146 564
rect 25210 552 25216 564
rect 25268 552 25274 604
rect 25946 552 25952 604
rect 26004 592 26010 604
rect 26314 592 26320 604
rect 26004 564 26320 592
rect 26004 552 26010 564
rect 26314 552 26320 564
rect 26372 552 26378 604
<< via1 >>
rect 10027 25542 10079 25594
rect 10091 25542 10143 25594
rect 10155 25542 10207 25594
rect 10219 25542 10271 25594
rect 19360 25542 19412 25594
rect 19424 25542 19476 25594
rect 19488 25542 19540 25594
rect 19552 25542 19604 25594
rect 5360 24998 5412 25050
rect 5424 24998 5476 25050
rect 5488 24998 5540 25050
rect 5552 24998 5604 25050
rect 14694 24998 14746 25050
rect 14758 24998 14810 25050
rect 14822 24998 14874 25050
rect 14886 24998 14938 25050
rect 24027 24998 24079 25050
rect 24091 24998 24143 25050
rect 24155 24998 24207 25050
rect 24219 24998 24271 25050
rect 10027 24454 10079 24506
rect 10091 24454 10143 24506
rect 10155 24454 10207 24506
rect 10219 24454 10271 24506
rect 19360 24454 19412 24506
rect 19424 24454 19476 24506
rect 19488 24454 19540 24506
rect 19552 24454 19604 24506
rect 24848 24352 24900 24404
rect 5360 23910 5412 23962
rect 5424 23910 5476 23962
rect 5488 23910 5540 23962
rect 5552 23910 5604 23962
rect 14694 23910 14746 23962
rect 14758 23910 14810 23962
rect 14822 23910 14874 23962
rect 14886 23910 14938 23962
rect 24027 23910 24079 23962
rect 24091 23910 24143 23962
rect 24155 23910 24207 23962
rect 24219 23910 24271 23962
rect 24480 23851 24532 23860
rect 24480 23817 24489 23851
rect 24489 23817 24523 23851
rect 24523 23817 24532 23851
rect 24480 23808 24532 23817
rect 23652 23604 23704 23656
rect 2492 23468 2544 23520
rect 3780 23468 3832 23520
rect 10027 23366 10079 23418
rect 10091 23366 10143 23418
rect 10155 23366 10207 23418
rect 10219 23366 10271 23418
rect 19360 23366 19412 23418
rect 19424 23366 19476 23418
rect 19488 23366 19540 23418
rect 19552 23366 19604 23418
rect 10680 23307 10732 23316
rect 10680 23273 10689 23307
rect 10689 23273 10723 23307
rect 10723 23273 10732 23307
rect 10680 23264 10732 23273
rect 24480 23307 24532 23316
rect 24480 23273 24489 23307
rect 24489 23273 24523 23307
rect 24523 23273 24532 23307
rect 24480 23264 24532 23273
rect 10496 23171 10548 23180
rect 10496 23137 10505 23171
rect 10505 23137 10539 23171
rect 10539 23137 10548 23171
rect 10496 23128 10548 23137
rect 23836 23128 23888 23180
rect 5360 22822 5412 22874
rect 5424 22822 5476 22874
rect 5488 22822 5540 22874
rect 5552 22822 5604 22874
rect 14694 22822 14746 22874
rect 14758 22822 14810 22874
rect 14822 22822 14874 22874
rect 14886 22822 14938 22874
rect 24027 22822 24079 22874
rect 24091 22822 24143 22874
rect 24155 22822 24207 22874
rect 24219 22822 24271 22874
rect 24572 22720 24624 22772
rect 23652 22627 23704 22636
rect 23652 22593 23661 22627
rect 23661 22593 23695 22627
rect 23695 22593 23704 22627
rect 23652 22584 23704 22593
rect 24664 22559 24716 22568
rect 24664 22525 24673 22559
rect 24673 22525 24707 22559
rect 24707 22525 24716 22559
rect 24664 22516 24716 22525
rect 23192 22491 23244 22500
rect 23192 22457 23201 22491
rect 23201 22457 23235 22491
rect 23235 22457 23244 22491
rect 23192 22448 23244 22457
rect 9760 22380 9812 22432
rect 10496 22423 10548 22432
rect 10496 22389 10505 22423
rect 10505 22389 10539 22423
rect 10539 22389 10548 22423
rect 10496 22380 10548 22389
rect 23836 22380 23888 22432
rect 24388 22423 24440 22432
rect 24388 22389 24397 22423
rect 24397 22389 24431 22423
rect 24431 22389 24440 22423
rect 24388 22380 24440 22389
rect 10027 22278 10079 22330
rect 10091 22278 10143 22330
rect 10155 22278 10207 22330
rect 10219 22278 10271 22330
rect 19360 22278 19412 22330
rect 19424 22278 19476 22330
rect 19488 22278 19540 22330
rect 19552 22278 19604 22330
rect 9760 22151 9812 22160
rect 9760 22117 9769 22151
rect 9769 22117 9803 22151
rect 9803 22117 9812 22151
rect 9760 22108 9812 22117
rect 9392 22040 9444 22092
rect 12336 22040 12388 22092
rect 24388 22040 24440 22092
rect 12428 22015 12480 22024
rect 12428 21981 12437 22015
rect 12437 21981 12471 22015
rect 12471 21981 12480 22015
rect 12428 21972 12480 21981
rect 23744 21904 23796 21956
rect 5360 21734 5412 21786
rect 5424 21734 5476 21786
rect 5488 21734 5540 21786
rect 5552 21734 5604 21786
rect 14694 21734 14746 21786
rect 14758 21734 14810 21786
rect 14822 21734 14874 21786
rect 14886 21734 14938 21786
rect 24027 21734 24079 21786
rect 24091 21734 24143 21786
rect 24155 21734 24207 21786
rect 24219 21734 24271 21786
rect 24480 21675 24532 21684
rect 24480 21641 24489 21675
rect 24489 21641 24523 21675
rect 24523 21641 24532 21675
rect 24480 21632 24532 21641
rect 24388 21496 24440 21548
rect 14728 21471 14780 21480
rect 14728 21437 14737 21471
rect 14737 21437 14771 21471
rect 14771 21437 14780 21471
rect 14728 21428 14780 21437
rect 24112 21471 24164 21480
rect 24112 21437 24121 21471
rect 24121 21437 24155 21471
rect 24155 21437 24164 21471
rect 24112 21428 24164 21437
rect 24296 21471 24348 21480
rect 24296 21437 24305 21471
rect 24305 21437 24339 21471
rect 24339 21437 24348 21471
rect 24296 21428 24348 21437
rect 15004 21403 15056 21412
rect 15004 21369 15013 21403
rect 15013 21369 15047 21403
rect 15047 21369 15056 21403
rect 15004 21360 15056 21369
rect 9392 21292 9444 21344
rect 12336 21335 12388 21344
rect 12336 21301 12345 21335
rect 12345 21301 12379 21335
rect 12379 21301 12388 21335
rect 12336 21292 12388 21301
rect 10027 21190 10079 21242
rect 10091 21190 10143 21242
rect 10155 21190 10207 21242
rect 10219 21190 10271 21242
rect 19360 21190 19412 21242
rect 19424 21190 19476 21242
rect 19488 21190 19540 21242
rect 19552 21190 19604 21242
rect 24756 21131 24808 21140
rect 24756 21097 24765 21131
rect 24765 21097 24799 21131
rect 24799 21097 24808 21131
rect 24756 21088 24808 21097
rect 24296 21020 24348 21072
rect 23192 20952 23244 21004
rect 24572 20995 24624 21004
rect 24572 20961 24581 20995
rect 24581 20961 24615 20995
rect 24615 20961 24624 20995
rect 24572 20952 24624 20961
rect 5360 20646 5412 20698
rect 5424 20646 5476 20698
rect 5488 20646 5540 20698
rect 5552 20646 5604 20698
rect 14694 20646 14746 20698
rect 14758 20646 14810 20698
rect 14822 20646 14874 20698
rect 14886 20646 14938 20698
rect 24027 20646 24079 20698
rect 24091 20646 24143 20698
rect 24155 20646 24207 20698
rect 24219 20646 24271 20698
rect 23560 20587 23612 20596
rect 23560 20553 23569 20587
rect 23569 20553 23603 20587
rect 23603 20553 23612 20587
rect 23560 20544 23612 20553
rect 23192 20383 23244 20392
rect 23192 20349 23201 20383
rect 23201 20349 23235 20383
rect 23235 20349 23244 20383
rect 23192 20340 23244 20349
rect 23376 20383 23428 20392
rect 23376 20349 23385 20383
rect 23385 20349 23419 20383
rect 23419 20349 23428 20383
rect 23376 20340 23428 20349
rect 24572 20247 24624 20256
rect 24572 20213 24581 20247
rect 24581 20213 24615 20247
rect 24615 20213 24624 20247
rect 24572 20204 24624 20213
rect 10027 20102 10079 20154
rect 10091 20102 10143 20154
rect 10155 20102 10207 20154
rect 10219 20102 10271 20154
rect 19360 20102 19412 20154
rect 19424 20102 19476 20154
rect 19488 20102 19540 20154
rect 19552 20102 19604 20154
rect 24388 20000 24440 20052
rect 21444 19975 21496 19984
rect 21444 19941 21453 19975
rect 21453 19941 21487 19975
rect 21487 19941 21496 19975
rect 21444 19932 21496 19941
rect 23376 19932 23428 19984
rect 21168 19907 21220 19916
rect 21168 19873 21177 19907
rect 21177 19873 21211 19907
rect 21211 19873 21220 19907
rect 21168 19864 21220 19873
rect 22456 19907 22508 19916
rect 22456 19873 22465 19907
rect 22465 19873 22499 19907
rect 22499 19873 22508 19907
rect 22456 19864 22508 19873
rect 24388 19864 24440 19916
rect 5360 19558 5412 19610
rect 5424 19558 5476 19610
rect 5488 19558 5540 19610
rect 5552 19558 5604 19610
rect 14694 19558 14746 19610
rect 14758 19558 14810 19610
rect 14822 19558 14874 19610
rect 14886 19558 14938 19610
rect 24027 19558 24079 19610
rect 24091 19558 24143 19610
rect 24155 19558 24207 19610
rect 24219 19558 24271 19610
rect 23652 19252 23704 19304
rect 20616 19116 20668 19168
rect 21168 19159 21220 19168
rect 21168 19125 21177 19159
rect 21177 19125 21211 19159
rect 21211 19125 21220 19159
rect 21168 19116 21220 19125
rect 22456 19159 22508 19168
rect 22456 19125 22465 19159
rect 22465 19125 22499 19159
rect 22499 19125 22508 19159
rect 22456 19116 22508 19125
rect 24112 19159 24164 19168
rect 24112 19125 24121 19159
rect 24121 19125 24155 19159
rect 24155 19125 24164 19159
rect 24112 19116 24164 19125
rect 24388 19116 24440 19168
rect 24480 19159 24532 19168
rect 24480 19125 24489 19159
rect 24489 19125 24523 19159
rect 24523 19125 24532 19159
rect 24480 19116 24532 19125
rect 10027 19014 10079 19066
rect 10091 19014 10143 19066
rect 10155 19014 10207 19066
rect 10219 19014 10271 19066
rect 19360 19014 19412 19066
rect 19424 19014 19476 19066
rect 19488 19014 19540 19066
rect 19552 19014 19604 19066
rect 11140 18955 11192 18964
rect 11140 18921 11149 18955
rect 11149 18921 11183 18955
rect 11183 18921 11192 18955
rect 11140 18912 11192 18921
rect 10772 18776 10824 18828
rect 15372 18776 15424 18828
rect 15740 18819 15792 18828
rect 15740 18785 15749 18819
rect 15749 18785 15783 18819
rect 15783 18785 15792 18819
rect 15740 18776 15792 18785
rect 5360 18470 5412 18522
rect 5424 18470 5476 18522
rect 5488 18470 5540 18522
rect 5552 18470 5604 18522
rect 14694 18470 14746 18522
rect 14758 18470 14810 18522
rect 14822 18470 14874 18522
rect 14886 18470 14938 18522
rect 24027 18470 24079 18522
rect 24091 18470 24143 18522
rect 24155 18470 24207 18522
rect 24219 18470 24271 18522
rect 24848 18411 24900 18420
rect 24848 18377 24857 18411
rect 24857 18377 24891 18411
rect 24891 18377 24900 18411
rect 24848 18368 24900 18377
rect 23652 18275 23704 18284
rect 23652 18241 23661 18275
rect 23661 18241 23695 18275
rect 23695 18241 23704 18275
rect 23652 18232 23704 18241
rect 23192 18164 23244 18216
rect 24664 18207 24716 18216
rect 24664 18173 24673 18207
rect 24673 18173 24707 18207
rect 24707 18173 24716 18207
rect 24664 18164 24716 18173
rect 10772 18028 10824 18080
rect 15372 18028 15424 18080
rect 10027 17926 10079 17978
rect 10091 17926 10143 17978
rect 10155 17926 10207 17978
rect 10219 17926 10271 17978
rect 19360 17926 19412 17978
rect 19424 17926 19476 17978
rect 19488 17926 19540 17978
rect 19552 17926 19604 17978
rect 10680 17756 10732 17808
rect 9852 17688 9904 17740
rect 15832 17731 15884 17740
rect 15832 17697 15841 17731
rect 15841 17697 15875 17731
rect 15875 17697 15884 17731
rect 15832 17688 15884 17697
rect 16016 17595 16068 17604
rect 16016 17561 16025 17595
rect 16025 17561 16059 17595
rect 16059 17561 16068 17595
rect 16016 17552 16068 17561
rect 5360 17382 5412 17434
rect 5424 17382 5476 17434
rect 5488 17382 5540 17434
rect 5552 17382 5604 17434
rect 14694 17382 14746 17434
rect 14758 17382 14810 17434
rect 14822 17382 14874 17434
rect 14886 17382 14938 17434
rect 24027 17382 24079 17434
rect 24091 17382 24143 17434
rect 24155 17382 24207 17434
rect 24219 17382 24271 17434
rect 24388 17280 24440 17332
rect 12152 17076 12204 17128
rect 24296 17119 24348 17128
rect 24296 17085 24305 17119
rect 24305 17085 24339 17119
rect 24339 17085 24348 17119
rect 24296 17076 24348 17085
rect 12888 17051 12940 17060
rect 12888 17017 12897 17051
rect 12897 17017 12931 17051
rect 12931 17017 12940 17051
rect 12888 17008 12940 17017
rect 9852 16940 9904 16992
rect 15832 16983 15884 16992
rect 15832 16949 15841 16983
rect 15841 16949 15875 16983
rect 15875 16949 15884 16983
rect 15832 16940 15884 16949
rect 10027 16838 10079 16890
rect 10091 16838 10143 16890
rect 10155 16838 10207 16890
rect 10219 16838 10271 16890
rect 19360 16838 19412 16890
rect 19424 16838 19476 16890
rect 19488 16838 19540 16890
rect 19552 16838 19604 16890
rect 24480 16779 24532 16788
rect 24480 16745 24489 16779
rect 24489 16745 24523 16779
rect 24523 16745 24532 16779
rect 24480 16736 24532 16745
rect 15832 16668 15884 16720
rect 15004 16643 15056 16652
rect 15004 16609 15013 16643
rect 15013 16609 15047 16643
rect 15047 16609 15056 16643
rect 15004 16600 15056 16609
rect 24388 16600 24440 16652
rect 5360 16294 5412 16346
rect 5424 16294 5476 16346
rect 5488 16294 5540 16346
rect 5552 16294 5604 16346
rect 14694 16294 14746 16346
rect 14758 16294 14810 16346
rect 14822 16294 14874 16346
rect 14886 16294 14938 16346
rect 24027 16294 24079 16346
rect 24091 16294 24143 16346
rect 24155 16294 24207 16346
rect 24219 16294 24271 16346
rect 23836 16192 23888 16244
rect 18224 16099 18276 16108
rect 18224 16065 18233 16099
rect 18233 16065 18267 16099
rect 18267 16065 18276 16099
rect 18224 16056 18276 16065
rect 15004 15895 15056 15904
rect 15004 15861 15013 15895
rect 15013 15861 15047 15895
rect 15047 15861 15056 15895
rect 15004 15852 15056 15861
rect 23836 15988 23888 16040
rect 18868 15852 18920 15904
rect 24112 15895 24164 15904
rect 24112 15861 24121 15895
rect 24121 15861 24155 15895
rect 24155 15861 24164 15895
rect 24112 15852 24164 15861
rect 24388 15852 24440 15904
rect 10027 15750 10079 15802
rect 10091 15750 10143 15802
rect 10155 15750 10207 15802
rect 10219 15750 10271 15802
rect 19360 15750 19412 15802
rect 19424 15750 19476 15802
rect 19488 15750 19540 15802
rect 19552 15750 19604 15802
rect 24112 15580 24164 15632
rect 22732 15512 22784 15564
rect 24388 15555 24440 15564
rect 24388 15521 24397 15555
rect 24397 15521 24431 15555
rect 24431 15521 24440 15555
rect 24388 15512 24440 15521
rect 26320 15308 26372 15360
rect 5360 15206 5412 15258
rect 5424 15206 5476 15258
rect 5488 15206 5540 15258
rect 5552 15206 5604 15258
rect 14694 15206 14746 15258
rect 14758 15206 14810 15258
rect 14822 15206 14874 15258
rect 14886 15206 14938 15258
rect 24027 15206 24079 15258
rect 24091 15206 24143 15258
rect 24155 15206 24207 15258
rect 24219 15206 24271 15258
rect 24388 15147 24440 15156
rect 24388 15113 24397 15147
rect 24397 15113 24431 15147
rect 24431 15113 24440 15147
rect 24388 15104 24440 15113
rect 24572 15104 24624 15156
rect 23836 15011 23888 15020
rect 23836 14977 23845 15011
rect 23845 14977 23879 15011
rect 23879 14977 23888 15011
rect 23836 14968 23888 14977
rect 23560 14943 23612 14952
rect 23560 14909 23569 14943
rect 23569 14909 23603 14943
rect 23603 14909 23612 14943
rect 23560 14900 23612 14909
rect 24848 14943 24900 14952
rect 24848 14909 24857 14943
rect 24857 14909 24891 14943
rect 24891 14909 24900 14943
rect 24848 14900 24900 14909
rect 22732 14807 22784 14816
rect 22732 14773 22741 14807
rect 22741 14773 22775 14807
rect 22775 14773 22784 14807
rect 22732 14764 22784 14773
rect 10027 14662 10079 14714
rect 10091 14662 10143 14714
rect 10155 14662 10207 14714
rect 10219 14662 10271 14714
rect 19360 14662 19412 14714
rect 19424 14662 19476 14714
rect 19488 14662 19540 14714
rect 19552 14662 19604 14714
rect 24664 14560 24716 14612
rect 24848 14492 24900 14544
rect 23100 14467 23152 14476
rect 23100 14433 23109 14467
rect 23109 14433 23143 14467
rect 23143 14433 23152 14467
rect 23100 14424 23152 14433
rect 24388 14467 24440 14476
rect 24388 14433 24397 14467
rect 24397 14433 24431 14467
rect 24431 14433 24440 14467
rect 24388 14424 24440 14433
rect 20984 14356 21036 14408
rect 5360 14118 5412 14170
rect 5424 14118 5476 14170
rect 5488 14118 5540 14170
rect 5552 14118 5604 14170
rect 14694 14118 14746 14170
rect 14758 14118 14810 14170
rect 14822 14118 14874 14170
rect 14886 14118 14938 14170
rect 24027 14118 24079 14170
rect 24091 14118 24143 14170
rect 24155 14118 24207 14170
rect 24219 14118 24271 14170
rect 23468 14016 23520 14068
rect 24848 13991 24900 14000
rect 24848 13957 24857 13991
rect 24857 13957 24891 13991
rect 24891 13957 24900 13991
rect 24848 13948 24900 13957
rect 18592 13923 18644 13932
rect 18592 13889 18601 13923
rect 18601 13889 18635 13923
rect 18635 13889 18644 13923
rect 18592 13880 18644 13889
rect 18776 13812 18828 13864
rect 21812 13812 21864 13864
rect 23100 13855 23152 13864
rect 23100 13821 23109 13855
rect 23109 13821 23143 13855
rect 23143 13821 23152 13855
rect 23100 13812 23152 13821
rect 20432 13676 20484 13728
rect 21904 13719 21956 13728
rect 21904 13685 21913 13719
rect 21913 13685 21947 13719
rect 21947 13685 21956 13719
rect 21904 13676 21956 13685
rect 23652 13676 23704 13728
rect 10027 13574 10079 13626
rect 10091 13574 10143 13626
rect 10155 13574 10207 13626
rect 10219 13574 10271 13626
rect 19360 13574 19412 13626
rect 19424 13574 19476 13626
rect 19488 13574 19540 13626
rect 19552 13574 19604 13626
rect 20616 13515 20668 13524
rect 20616 13481 20625 13515
rect 20625 13481 20659 13515
rect 20659 13481 20668 13515
rect 20616 13472 20668 13481
rect 20984 13515 21036 13524
rect 20984 13481 20993 13515
rect 20993 13481 21027 13515
rect 21027 13481 21036 13515
rect 20984 13472 21036 13481
rect 23192 13472 23244 13524
rect 23284 13472 23336 13524
rect 22916 13336 22968 13388
rect 24388 13336 24440 13388
rect 19236 13311 19288 13320
rect 19236 13277 19245 13311
rect 19245 13277 19279 13311
rect 19279 13277 19288 13311
rect 19236 13268 19288 13277
rect 19420 13132 19472 13184
rect 20524 13132 20576 13184
rect 21352 13268 21404 13320
rect 23100 13311 23152 13320
rect 23100 13277 23109 13311
rect 23109 13277 23143 13311
rect 23143 13277 23152 13311
rect 23100 13268 23152 13277
rect 22180 13132 22232 13184
rect 23376 13132 23428 13184
rect 5360 13030 5412 13082
rect 5424 13030 5476 13082
rect 5488 13030 5540 13082
rect 5552 13030 5604 13082
rect 14694 13030 14746 13082
rect 14758 13030 14810 13082
rect 14822 13030 14874 13082
rect 14886 13030 14938 13082
rect 24027 13030 24079 13082
rect 24091 13030 24143 13082
rect 24155 13030 24207 13082
rect 24219 13030 24271 13082
rect 18960 12971 19012 12980
rect 18960 12937 18969 12971
rect 18969 12937 19003 12971
rect 19003 12937 19012 12971
rect 18960 12928 19012 12937
rect 20984 12928 21036 12980
rect 22916 12928 22968 12980
rect 23192 12971 23244 12980
rect 23192 12937 23201 12971
rect 23201 12937 23235 12971
rect 23235 12937 23244 12971
rect 23192 12928 23244 12937
rect 24848 12971 24900 12980
rect 24848 12937 24857 12971
rect 24857 12937 24891 12971
rect 24891 12937 24900 12971
rect 24848 12928 24900 12937
rect 25308 12971 25360 12980
rect 25308 12937 25317 12971
rect 25317 12937 25351 12971
rect 25351 12937 25360 12971
rect 25308 12928 25360 12937
rect 24296 12903 24348 12912
rect 24296 12869 24305 12903
rect 24305 12869 24339 12903
rect 24339 12869 24348 12903
rect 24296 12860 24348 12869
rect 19144 12792 19196 12844
rect 19420 12835 19472 12844
rect 19420 12801 19429 12835
rect 19429 12801 19463 12835
rect 19463 12801 19472 12835
rect 19420 12792 19472 12801
rect 21168 12835 21220 12844
rect 21168 12801 21177 12835
rect 21177 12801 21211 12835
rect 21211 12801 21220 12835
rect 21168 12792 21220 12801
rect 23652 12835 23704 12844
rect 23652 12801 23661 12835
rect 23661 12801 23695 12835
rect 23695 12801 23704 12835
rect 23652 12792 23704 12801
rect 19788 12724 19840 12776
rect 21076 12724 21128 12776
rect 23376 12767 23428 12776
rect 23376 12733 23385 12767
rect 23385 12733 23419 12767
rect 23419 12733 23428 12767
rect 23376 12724 23428 12733
rect 25308 12724 25360 12776
rect 18592 12656 18644 12708
rect 16476 12588 16528 12640
rect 20524 12631 20576 12640
rect 20524 12597 20533 12631
rect 20533 12597 20567 12631
rect 20567 12597 20576 12631
rect 20524 12588 20576 12597
rect 21812 12588 21864 12640
rect 10027 12486 10079 12538
rect 10091 12486 10143 12538
rect 10155 12486 10207 12538
rect 10219 12486 10271 12538
rect 19360 12486 19412 12538
rect 19424 12486 19476 12538
rect 19488 12486 19540 12538
rect 19552 12486 19604 12538
rect 18500 12384 18552 12436
rect 18868 12384 18920 12436
rect 21352 12384 21404 12436
rect 22640 12427 22692 12436
rect 22640 12393 22649 12427
rect 22649 12393 22683 12427
rect 22683 12393 22692 12427
rect 22640 12384 22692 12393
rect 23100 12384 23152 12436
rect 16660 12359 16712 12368
rect 16660 12325 16669 12359
rect 16669 12325 16703 12359
rect 16703 12325 16712 12359
rect 16660 12316 16712 12325
rect 17856 12316 17908 12368
rect 16384 12291 16436 12300
rect 16384 12257 16393 12291
rect 16393 12257 16427 12291
rect 16427 12257 16436 12291
rect 16384 12248 16436 12257
rect 18684 12248 18736 12300
rect 21168 12248 21220 12300
rect 18868 12044 18920 12096
rect 19604 12044 19656 12096
rect 24756 12248 24808 12300
rect 21996 12155 22048 12164
rect 21996 12121 22005 12155
rect 22005 12121 22039 12155
rect 22039 12121 22048 12155
rect 21996 12112 22048 12121
rect 22088 12044 22140 12096
rect 5360 11942 5412 11994
rect 5424 11942 5476 11994
rect 5488 11942 5540 11994
rect 5552 11942 5604 11994
rect 14694 11942 14746 11994
rect 14758 11942 14810 11994
rect 14822 11942 14874 11994
rect 14886 11942 14938 11994
rect 24027 11942 24079 11994
rect 24091 11942 24143 11994
rect 24155 11942 24207 11994
rect 24219 11942 24271 11994
rect 21168 11840 21220 11892
rect 22824 11883 22876 11892
rect 22824 11849 22833 11883
rect 22833 11849 22867 11883
rect 22867 11849 22876 11883
rect 22824 11840 22876 11849
rect 24480 11883 24532 11892
rect 16384 11772 16436 11824
rect 15924 11747 15976 11756
rect 15924 11713 15933 11747
rect 15933 11713 15967 11747
rect 15967 11713 15976 11747
rect 15924 11704 15976 11713
rect 17856 11704 17908 11756
rect 19604 11747 19656 11756
rect 19604 11713 19613 11747
rect 19613 11713 19647 11747
rect 19647 11713 19656 11747
rect 19604 11704 19656 11713
rect 24480 11849 24489 11883
rect 24489 11849 24523 11883
rect 24523 11849 24532 11883
rect 24480 11840 24532 11849
rect 24756 11883 24808 11892
rect 24756 11849 24765 11883
rect 24765 11849 24799 11883
rect 24799 11849 24808 11883
rect 24756 11840 24808 11849
rect 25124 11883 25176 11892
rect 25124 11849 25133 11883
rect 25133 11849 25167 11883
rect 25167 11849 25176 11883
rect 25124 11840 25176 11849
rect 23928 11747 23980 11756
rect 23928 11713 23937 11747
rect 23937 11713 23971 11747
rect 23971 11713 23980 11747
rect 23928 11704 23980 11713
rect 18684 11636 18736 11688
rect 22824 11636 22876 11688
rect 24940 11679 24992 11688
rect 24940 11645 24949 11679
rect 24949 11645 24983 11679
rect 24983 11645 24992 11679
rect 24940 11636 24992 11645
rect 16016 11568 16068 11620
rect 22916 11568 22968 11620
rect 17856 11500 17908 11552
rect 18316 11500 18368 11552
rect 19696 11500 19748 11552
rect 22088 11500 22140 11552
rect 22364 11543 22416 11552
rect 22364 11509 22373 11543
rect 22373 11509 22407 11543
rect 22407 11509 22416 11543
rect 22364 11500 22416 11509
rect 23192 11543 23244 11552
rect 23192 11509 23201 11543
rect 23201 11509 23235 11543
rect 23235 11509 23244 11543
rect 23192 11500 23244 11509
rect 23376 11543 23428 11552
rect 23376 11509 23385 11543
rect 23385 11509 23419 11543
rect 23419 11509 23428 11543
rect 23376 11500 23428 11509
rect 10027 11398 10079 11450
rect 10091 11398 10143 11450
rect 10155 11398 10207 11450
rect 10219 11398 10271 11450
rect 19360 11398 19412 11450
rect 19424 11398 19476 11450
rect 19488 11398 19540 11450
rect 19552 11398 19604 11450
rect 17856 11339 17908 11348
rect 17856 11305 17865 11339
rect 17865 11305 17899 11339
rect 17899 11305 17908 11339
rect 17856 11296 17908 11305
rect 18960 11339 19012 11348
rect 18960 11305 18969 11339
rect 18969 11305 19003 11339
rect 19003 11305 19012 11339
rect 18960 11296 19012 11305
rect 19052 11296 19104 11348
rect 19236 11296 19288 11348
rect 20432 11296 20484 11348
rect 13624 11203 13676 11212
rect 13624 11169 13633 11203
rect 13633 11169 13667 11203
rect 13667 11169 13676 11203
rect 13624 11160 13676 11169
rect 15004 11203 15056 11212
rect 15004 11169 15013 11203
rect 15013 11169 15047 11203
rect 15047 11169 15056 11203
rect 15004 11160 15056 11169
rect 15280 11203 15332 11212
rect 15280 11169 15289 11203
rect 15289 11169 15323 11203
rect 15323 11169 15332 11203
rect 15280 11160 15332 11169
rect 15832 11203 15884 11212
rect 15832 11169 15841 11203
rect 15841 11169 15875 11203
rect 15875 11169 15884 11203
rect 17396 11228 17448 11280
rect 18868 11271 18920 11280
rect 18868 11237 18877 11271
rect 18877 11237 18911 11271
rect 18911 11237 18920 11271
rect 18868 11228 18920 11237
rect 20524 11228 20576 11280
rect 22640 11228 22692 11280
rect 15832 11160 15884 11169
rect 16568 11160 16620 11212
rect 19880 11160 19932 11212
rect 25400 11160 25452 11212
rect 13716 11092 13768 11144
rect 19512 11135 19564 11144
rect 19512 11101 19521 11135
rect 19521 11101 19555 11135
rect 19555 11101 19564 11135
rect 19512 11092 19564 11101
rect 21168 11092 21220 11144
rect 21996 11092 22048 11144
rect 22088 11092 22140 11144
rect 18316 11024 18368 11076
rect 20616 11067 20668 11076
rect 20616 11033 20625 11067
rect 20625 11033 20659 11067
rect 20659 11033 20668 11067
rect 20616 11024 20668 11033
rect 24940 11067 24992 11076
rect 24940 11033 24949 11067
rect 24949 11033 24983 11067
rect 24983 11033 24992 11067
rect 24940 11024 24992 11033
rect 16660 10956 16712 11008
rect 22272 10956 22324 11008
rect 23928 10956 23980 11008
rect 24756 10956 24808 11008
rect 5360 10854 5412 10906
rect 5424 10854 5476 10906
rect 5488 10854 5540 10906
rect 5552 10854 5604 10906
rect 14694 10854 14746 10906
rect 14758 10854 14810 10906
rect 14822 10854 14874 10906
rect 14886 10854 14938 10906
rect 24027 10854 24079 10906
rect 24091 10854 24143 10906
rect 24155 10854 24207 10906
rect 24219 10854 24271 10906
rect 13440 10752 13492 10804
rect 16108 10795 16160 10804
rect 16108 10761 16117 10795
rect 16117 10761 16151 10795
rect 16151 10761 16160 10795
rect 16108 10752 16160 10761
rect 18960 10752 19012 10804
rect 20432 10752 20484 10804
rect 21168 10795 21220 10804
rect 21168 10761 21177 10795
rect 21177 10761 21211 10795
rect 21211 10761 21220 10795
rect 21168 10752 21220 10761
rect 21904 10752 21956 10804
rect 22640 10752 22692 10804
rect 25400 10795 25452 10804
rect 25400 10761 25409 10795
rect 25409 10761 25443 10795
rect 25443 10761 25452 10795
rect 25400 10752 25452 10761
rect 15004 10684 15056 10736
rect 21720 10727 21772 10736
rect 21720 10693 21729 10727
rect 21729 10693 21763 10727
rect 21763 10693 21772 10727
rect 21720 10684 21772 10693
rect 14728 10659 14780 10668
rect 14728 10625 14737 10659
rect 14737 10625 14771 10659
rect 14771 10625 14780 10659
rect 14728 10616 14780 10625
rect 16660 10659 16712 10668
rect 16660 10625 16669 10659
rect 16669 10625 16703 10659
rect 16703 10625 16712 10659
rect 16660 10616 16712 10625
rect 17672 10616 17724 10668
rect 18684 10616 18736 10668
rect 22272 10659 22324 10668
rect 22272 10625 22281 10659
rect 22281 10625 22315 10659
rect 22315 10625 22324 10659
rect 22272 10616 22324 10625
rect 16476 10591 16528 10600
rect 16476 10557 16485 10591
rect 16485 10557 16519 10591
rect 16519 10557 16528 10591
rect 16476 10548 16528 10557
rect 16568 10548 16620 10600
rect 17396 10548 17448 10600
rect 18868 10548 18920 10600
rect 22180 10591 22232 10600
rect 22180 10557 22189 10591
rect 22189 10557 22223 10591
rect 22223 10557 22232 10591
rect 22180 10548 22232 10557
rect 23284 10548 23336 10600
rect 13900 10480 13952 10532
rect 14360 10412 14412 10464
rect 19512 10480 19564 10532
rect 16660 10412 16712 10464
rect 17764 10455 17816 10464
rect 17764 10421 17773 10455
rect 17773 10421 17807 10455
rect 17807 10421 17816 10455
rect 17764 10412 17816 10421
rect 21904 10480 21956 10532
rect 24756 10455 24808 10464
rect 24756 10421 24765 10455
rect 24765 10421 24799 10455
rect 24799 10421 24808 10455
rect 24756 10412 24808 10421
rect 10027 10310 10079 10362
rect 10091 10310 10143 10362
rect 10155 10310 10207 10362
rect 10219 10310 10271 10362
rect 19360 10310 19412 10362
rect 19424 10310 19476 10362
rect 19488 10310 19540 10362
rect 19552 10310 19604 10362
rect 13900 10251 13952 10260
rect 13900 10217 13909 10251
rect 13909 10217 13943 10251
rect 13943 10217 13952 10251
rect 13900 10208 13952 10217
rect 17396 10251 17448 10260
rect 17396 10217 17405 10251
rect 17405 10217 17439 10251
rect 17439 10217 17448 10251
rect 17396 10208 17448 10217
rect 19880 10251 19932 10260
rect 19880 10217 19889 10251
rect 19889 10217 19923 10251
rect 19923 10217 19932 10251
rect 19880 10208 19932 10217
rect 20524 10208 20576 10260
rect 21628 10208 21680 10260
rect 22180 10208 22232 10260
rect 23376 10208 23428 10260
rect 14728 10140 14780 10192
rect 15004 10140 15056 10192
rect 19144 10140 19196 10192
rect 24756 10140 24808 10192
rect 15096 10115 15148 10124
rect 15096 10081 15105 10115
rect 15105 10081 15139 10115
rect 15139 10081 15148 10115
rect 15096 10072 15148 10081
rect 15832 10072 15884 10124
rect 18868 10072 18920 10124
rect 19052 10072 19104 10124
rect 21168 10115 21220 10124
rect 21168 10081 21177 10115
rect 21177 10081 21211 10115
rect 21211 10081 21220 10115
rect 21168 10072 21220 10081
rect 17856 10047 17908 10056
rect 17856 10013 17865 10047
rect 17865 10013 17899 10047
rect 17899 10013 17908 10047
rect 17856 10004 17908 10013
rect 17580 9936 17632 9988
rect 21260 10047 21312 10056
rect 21260 10013 21269 10047
rect 21269 10013 21303 10047
rect 21303 10013 21312 10047
rect 21260 10004 21312 10013
rect 21720 10004 21772 10056
rect 23284 10047 23336 10056
rect 13624 9911 13676 9920
rect 13624 9877 13633 9911
rect 13633 9877 13667 9911
rect 13667 9877 13676 9911
rect 13624 9868 13676 9877
rect 14360 9911 14412 9920
rect 14360 9877 14369 9911
rect 14369 9877 14403 9911
rect 14403 9877 14412 9911
rect 14360 9868 14412 9877
rect 16568 9868 16620 9920
rect 18316 9911 18368 9920
rect 18316 9877 18325 9911
rect 18325 9877 18359 9911
rect 18359 9877 18368 9911
rect 18316 9868 18368 9877
rect 18960 9868 19012 9920
rect 22272 9911 22324 9920
rect 22272 9877 22281 9911
rect 22281 9877 22315 9911
rect 22315 9877 22324 9911
rect 23284 10013 23293 10047
rect 23293 10013 23327 10047
rect 23327 10013 23336 10047
rect 23284 10004 23336 10013
rect 22272 9868 22324 9877
rect 24480 9868 24532 9920
rect 5360 9766 5412 9818
rect 5424 9766 5476 9818
rect 5488 9766 5540 9818
rect 5552 9766 5604 9818
rect 14694 9766 14746 9818
rect 14758 9766 14810 9818
rect 14822 9766 14874 9818
rect 14886 9766 14938 9818
rect 24027 9766 24079 9818
rect 24091 9766 24143 9818
rect 24155 9766 24207 9818
rect 24219 9766 24271 9818
rect 15004 9707 15056 9716
rect 15004 9673 15013 9707
rect 15013 9673 15047 9707
rect 15047 9673 15056 9707
rect 15004 9664 15056 9673
rect 16660 9664 16712 9716
rect 24756 9707 24808 9716
rect 16200 9596 16252 9648
rect 24756 9673 24765 9707
rect 24765 9673 24799 9707
rect 24799 9673 24808 9707
rect 24756 9664 24808 9673
rect 18316 9596 18368 9648
rect 21352 9596 21404 9648
rect 22824 9639 22876 9648
rect 22824 9605 22833 9639
rect 22833 9605 22867 9639
rect 22867 9605 22876 9639
rect 22824 9596 22876 9605
rect 23376 9596 23428 9648
rect 24480 9639 24532 9648
rect 13624 9571 13676 9580
rect 13624 9537 13633 9571
rect 13633 9537 13667 9571
rect 13667 9537 13676 9571
rect 13624 9528 13676 9537
rect 16568 9528 16620 9580
rect 17948 9528 18000 9580
rect 18960 9460 19012 9512
rect 19604 9460 19656 9512
rect 13532 9435 13584 9444
rect 13532 9401 13541 9435
rect 13541 9401 13575 9435
rect 13575 9401 13584 9435
rect 13532 9392 13584 9401
rect 17488 9435 17540 9444
rect 17488 9401 17497 9435
rect 17497 9401 17531 9435
rect 17531 9401 17540 9435
rect 17488 9392 17540 9401
rect 18592 9392 18644 9444
rect 19788 9460 19840 9512
rect 23192 9571 23244 9580
rect 23192 9537 23201 9571
rect 23201 9537 23235 9571
rect 23235 9537 23244 9571
rect 23192 9528 23244 9537
rect 23744 9528 23796 9580
rect 24480 9605 24489 9639
rect 24489 9605 24523 9639
rect 24523 9605 24532 9639
rect 24480 9596 24532 9605
rect 24020 9571 24072 9580
rect 24020 9537 24029 9571
rect 24029 9537 24063 9571
rect 24063 9537 24072 9571
rect 24020 9528 24072 9537
rect 10956 9324 11008 9376
rect 12612 9367 12664 9376
rect 12612 9333 12621 9367
rect 12621 9333 12655 9367
rect 12655 9333 12664 9367
rect 12612 9324 12664 9333
rect 15924 9367 15976 9376
rect 15924 9333 15933 9367
rect 15933 9333 15967 9367
rect 15967 9333 15976 9367
rect 15924 9324 15976 9333
rect 16660 9324 16712 9376
rect 18224 9367 18276 9376
rect 18224 9333 18233 9367
rect 18233 9333 18267 9367
rect 18267 9333 18276 9367
rect 18224 9324 18276 9333
rect 18316 9324 18368 9376
rect 18500 9324 18552 9376
rect 18868 9367 18920 9376
rect 18868 9333 18877 9367
rect 18877 9333 18911 9367
rect 18911 9333 18920 9367
rect 18868 9324 18920 9333
rect 20340 9392 20392 9444
rect 21260 9392 21312 9444
rect 21720 9367 21772 9376
rect 21720 9333 21729 9367
rect 21729 9333 21763 9367
rect 21763 9333 21772 9367
rect 21720 9324 21772 9333
rect 22364 9367 22416 9376
rect 22364 9333 22373 9367
rect 22373 9333 22407 9367
rect 22407 9333 22416 9367
rect 22364 9324 22416 9333
rect 23744 9435 23796 9444
rect 23744 9401 23753 9435
rect 23753 9401 23787 9435
rect 23787 9401 23796 9435
rect 23744 9392 23796 9401
rect 23468 9324 23520 9376
rect 10027 9222 10079 9274
rect 10091 9222 10143 9274
rect 10155 9222 10207 9274
rect 10219 9222 10271 9274
rect 19360 9222 19412 9274
rect 19424 9222 19476 9274
rect 19488 9222 19540 9274
rect 19552 9222 19604 9274
rect 10588 9163 10640 9172
rect 10588 9129 10597 9163
rect 10597 9129 10631 9163
rect 10631 9129 10640 9163
rect 10588 9120 10640 9129
rect 13532 9163 13584 9172
rect 10956 9027 11008 9036
rect 10956 8993 10965 9027
rect 10965 8993 10999 9027
rect 10999 8993 11008 9027
rect 10956 8984 11008 8993
rect 10496 8823 10548 8832
rect 10496 8789 10505 8823
rect 10505 8789 10539 8823
rect 10539 8789 10548 8823
rect 11784 8916 11836 8968
rect 12060 8916 12112 8968
rect 12336 9052 12388 9104
rect 13532 9129 13541 9163
rect 13541 9129 13575 9163
rect 13575 9129 13584 9163
rect 14084 9163 14136 9172
rect 13532 9120 13584 9129
rect 14084 9129 14093 9163
rect 14093 9129 14127 9163
rect 14127 9129 14136 9163
rect 14084 9120 14136 9129
rect 15372 9120 15424 9172
rect 16568 9163 16620 9172
rect 16568 9129 16577 9163
rect 16577 9129 16611 9163
rect 16611 9129 16620 9163
rect 16568 9120 16620 9129
rect 17488 9120 17540 9172
rect 17672 9120 17724 9172
rect 18500 9120 18552 9172
rect 19788 9163 19840 9172
rect 19788 9129 19797 9163
rect 19797 9129 19831 9163
rect 19831 9129 19840 9163
rect 19788 9120 19840 9129
rect 21168 9120 21220 9172
rect 21812 9163 21864 9172
rect 21812 9129 21821 9163
rect 21821 9129 21855 9163
rect 21855 9129 21864 9163
rect 21812 9120 21864 9129
rect 13624 9052 13676 9104
rect 16660 9052 16712 9104
rect 17396 9052 17448 9104
rect 17948 9052 18000 9104
rect 23192 9052 23244 9104
rect 24020 9052 24072 9104
rect 15372 9027 15424 9036
rect 15372 8993 15381 9027
rect 15381 8993 15415 9027
rect 15415 8993 15424 9027
rect 15372 8984 15424 8993
rect 15464 9027 15516 9036
rect 15464 8993 15473 9027
rect 15473 8993 15507 9027
rect 15507 8993 15516 9027
rect 15464 8984 15516 8993
rect 16752 8984 16804 9036
rect 20984 9027 21036 9036
rect 20984 8993 20993 9027
rect 20993 8993 21027 9027
rect 21027 8993 21036 9027
rect 20984 8984 21036 8993
rect 15556 8959 15608 8968
rect 15556 8925 15565 8959
rect 15565 8925 15599 8959
rect 15599 8925 15608 8959
rect 15556 8916 15608 8925
rect 17212 8848 17264 8900
rect 20616 8916 20668 8968
rect 20800 8848 20852 8900
rect 21628 8848 21680 8900
rect 22272 8848 22324 8900
rect 10496 8780 10548 8789
rect 19144 8780 19196 8832
rect 20892 8780 20944 8832
rect 22180 8823 22232 8832
rect 22180 8789 22189 8823
rect 22189 8789 22223 8823
rect 22223 8789 22232 8823
rect 22180 8780 22232 8789
rect 23376 8780 23428 8832
rect 23744 8780 23796 8832
rect 24664 8780 24716 8832
rect 5360 8678 5412 8730
rect 5424 8678 5476 8730
rect 5488 8678 5540 8730
rect 5552 8678 5604 8730
rect 14694 8678 14746 8730
rect 14758 8678 14810 8730
rect 14822 8678 14874 8730
rect 14886 8678 14938 8730
rect 24027 8678 24079 8730
rect 24091 8678 24143 8730
rect 24155 8678 24207 8730
rect 24219 8678 24271 8730
rect 10956 8576 11008 8628
rect 11784 8619 11836 8628
rect 11784 8585 11793 8619
rect 11793 8585 11827 8619
rect 11827 8585 11836 8619
rect 11784 8576 11836 8585
rect 12336 8576 12388 8628
rect 14360 8576 14412 8628
rect 15372 8576 15424 8628
rect 17396 8619 17448 8628
rect 17396 8585 17405 8619
rect 17405 8585 17439 8619
rect 17439 8585 17448 8619
rect 17396 8576 17448 8585
rect 18500 8619 18552 8628
rect 18500 8585 18509 8619
rect 18509 8585 18543 8619
rect 18543 8585 18552 8619
rect 18500 8576 18552 8585
rect 19788 8576 19840 8628
rect 20616 8619 20668 8628
rect 20616 8585 20625 8619
rect 20625 8585 20659 8619
rect 20659 8585 20668 8619
rect 20616 8576 20668 8585
rect 21536 8576 21588 8628
rect 20340 8508 20392 8560
rect 14084 8483 14136 8492
rect 14084 8449 14093 8483
rect 14093 8449 14127 8483
rect 14127 8449 14136 8483
rect 14084 8440 14136 8449
rect 15096 8440 15148 8492
rect 18592 8483 18644 8492
rect 18592 8449 18601 8483
rect 18601 8449 18635 8483
rect 18635 8449 18644 8483
rect 18592 8440 18644 8449
rect 22180 8483 22232 8492
rect 22180 8449 22189 8483
rect 22189 8449 22223 8483
rect 22223 8449 22232 8483
rect 22180 8440 22232 8449
rect 23192 8551 23244 8560
rect 23192 8517 23201 8551
rect 23201 8517 23235 8551
rect 23235 8517 23244 8551
rect 23192 8508 23244 8517
rect 10680 8372 10732 8424
rect 14268 8372 14320 8424
rect 18500 8372 18552 8424
rect 21904 8372 21956 8424
rect 23192 8372 23244 8424
rect 23376 8415 23428 8424
rect 23376 8381 23385 8415
rect 23385 8381 23419 8415
rect 23419 8381 23428 8415
rect 23376 8372 23428 8381
rect 24664 8372 24716 8424
rect 9576 8304 9628 8356
rect 13348 8347 13400 8356
rect 13348 8313 13357 8347
rect 13357 8313 13391 8347
rect 13391 8313 13400 8347
rect 13348 8304 13400 8313
rect 14820 8304 14872 8356
rect 15556 8304 15608 8356
rect 10956 8236 11008 8288
rect 12520 8236 12572 8288
rect 16752 8304 16804 8356
rect 20984 8347 21036 8356
rect 20984 8313 20993 8347
rect 20993 8313 21027 8347
rect 21027 8313 21036 8347
rect 20984 8304 21036 8313
rect 22456 8304 22508 8356
rect 23744 8304 23796 8356
rect 16384 8236 16436 8288
rect 10027 8134 10079 8186
rect 10091 8134 10143 8186
rect 10155 8134 10207 8186
rect 10219 8134 10271 8186
rect 19360 8134 19412 8186
rect 19424 8134 19476 8186
rect 19488 8134 19540 8186
rect 19552 8134 19604 8186
rect 11784 8032 11836 8084
rect 13164 8075 13216 8084
rect 13164 8041 13173 8075
rect 13173 8041 13207 8075
rect 13207 8041 13216 8075
rect 13164 8032 13216 8041
rect 14820 8075 14872 8084
rect 14820 8041 14829 8075
rect 14829 8041 14863 8075
rect 14863 8041 14872 8075
rect 14820 8032 14872 8041
rect 16384 8075 16436 8084
rect 16384 8041 16393 8075
rect 16393 8041 16427 8075
rect 16427 8041 16436 8075
rect 16384 8032 16436 8041
rect 17764 8032 17816 8084
rect 10956 7939 11008 7948
rect 10956 7905 10990 7939
rect 10990 7905 11008 7939
rect 10956 7896 11008 7905
rect 12520 7896 12572 7948
rect 14544 7896 14596 7948
rect 17856 7896 17908 7948
rect 9760 7828 9812 7880
rect 10680 7871 10732 7880
rect 10680 7837 10689 7871
rect 10689 7837 10723 7871
rect 10723 7837 10732 7871
rect 10680 7828 10732 7837
rect 13624 7871 13676 7880
rect 13624 7837 13633 7871
rect 13633 7837 13667 7871
rect 13667 7837 13676 7871
rect 13624 7828 13676 7837
rect 15004 7871 15056 7880
rect 12980 7760 13032 7812
rect 15004 7837 15013 7871
rect 15013 7837 15047 7871
rect 15047 7837 15056 7871
rect 15004 7828 15056 7837
rect 20340 8032 20392 8084
rect 23192 8075 23244 8084
rect 23192 8041 23201 8075
rect 23201 8041 23235 8075
rect 23235 8041 23244 8075
rect 23192 8032 23244 8041
rect 23652 8075 23704 8084
rect 23652 8041 23661 8075
rect 23661 8041 23695 8075
rect 23695 8041 23704 8075
rect 23652 8032 23704 8041
rect 24664 8075 24716 8084
rect 24664 8041 24673 8075
rect 24673 8041 24707 8075
rect 24707 8041 24716 8075
rect 24664 8032 24716 8041
rect 20432 7964 20484 8016
rect 21628 7964 21680 8016
rect 21352 7896 21404 7948
rect 23100 7896 23152 7948
rect 24572 7896 24624 7948
rect 18316 7828 18368 7880
rect 18592 7828 18644 7880
rect 19880 7828 19932 7880
rect 23744 7871 23796 7880
rect 23744 7837 23753 7871
rect 23753 7837 23787 7871
rect 23787 7837 23796 7871
rect 23744 7828 23796 7837
rect 23928 7828 23980 7880
rect 24664 7828 24716 7880
rect 19236 7760 19288 7812
rect 24940 7803 24992 7812
rect 7828 7735 7880 7744
rect 7828 7701 7837 7735
rect 7837 7701 7871 7735
rect 7871 7701 7880 7735
rect 7828 7692 7880 7701
rect 17212 7692 17264 7744
rect 18316 7692 18368 7744
rect 20800 7692 20852 7744
rect 20892 7692 20944 7744
rect 24940 7769 24949 7803
rect 24949 7769 24983 7803
rect 24983 7769 24992 7803
rect 24940 7760 24992 7769
rect 21996 7735 22048 7744
rect 21996 7701 22005 7735
rect 22005 7701 22039 7735
rect 22039 7701 22048 7735
rect 21996 7692 22048 7701
rect 22180 7692 22232 7744
rect 22916 7735 22968 7744
rect 22916 7701 22925 7735
rect 22925 7701 22959 7735
rect 22959 7701 22968 7735
rect 22916 7692 22968 7701
rect 23928 7692 23980 7744
rect 5360 7590 5412 7642
rect 5424 7590 5476 7642
rect 5488 7590 5540 7642
rect 5552 7590 5604 7642
rect 14694 7590 14746 7642
rect 14758 7590 14810 7642
rect 14822 7590 14874 7642
rect 14886 7590 14938 7642
rect 24027 7590 24079 7642
rect 24091 7590 24143 7642
rect 24155 7590 24207 7642
rect 24219 7590 24271 7642
rect 3872 7488 3924 7540
rect 5160 7488 5212 7540
rect 8012 7488 8064 7540
rect 10496 7531 10548 7540
rect 10496 7497 10505 7531
rect 10505 7497 10539 7531
rect 10539 7497 10548 7531
rect 10496 7488 10548 7497
rect 12520 7531 12572 7540
rect 12520 7497 12529 7531
rect 12529 7497 12563 7531
rect 12563 7497 12572 7531
rect 12520 7488 12572 7497
rect 15188 7488 15240 7540
rect 20800 7531 20852 7540
rect 20800 7497 20809 7531
rect 20809 7497 20843 7531
rect 20843 7497 20852 7531
rect 20800 7488 20852 7497
rect 21260 7488 21312 7540
rect 21352 7488 21404 7540
rect 22456 7531 22508 7540
rect 22456 7497 22465 7531
rect 22465 7497 22499 7531
rect 22499 7497 22508 7531
rect 22456 7488 22508 7497
rect 23652 7488 23704 7540
rect 24572 7488 24624 7540
rect 25676 7531 25728 7540
rect 25676 7497 25685 7531
rect 25685 7497 25719 7531
rect 25719 7497 25728 7531
rect 25676 7488 25728 7497
rect 25952 7488 26004 7540
rect 26596 7488 26648 7540
rect 9208 7463 9260 7472
rect 9208 7429 9217 7463
rect 9217 7429 9251 7463
rect 9251 7429 9260 7463
rect 9208 7420 9260 7429
rect 14360 7420 14412 7472
rect 16752 7420 16804 7472
rect 19144 7420 19196 7472
rect 10956 7352 11008 7404
rect 12060 7352 12112 7404
rect 18316 7395 18368 7404
rect 18316 7361 18325 7395
rect 18325 7361 18359 7395
rect 18359 7361 18368 7395
rect 18316 7352 18368 7361
rect 19972 7395 20024 7404
rect 19972 7361 19981 7395
rect 19981 7361 20015 7395
rect 20015 7361 20024 7395
rect 19972 7352 20024 7361
rect 20156 7352 20208 7404
rect 23100 7463 23152 7472
rect 23100 7429 23109 7463
rect 23109 7429 23143 7463
rect 23143 7429 23152 7463
rect 23100 7420 23152 7429
rect 21444 7395 21496 7404
rect 21444 7361 21453 7395
rect 21453 7361 21487 7395
rect 21487 7361 21496 7395
rect 21444 7352 21496 7361
rect 24020 7395 24072 7404
rect 24020 7361 24029 7395
rect 24029 7361 24063 7395
rect 24063 7361 24072 7395
rect 24020 7352 24072 7361
rect 7828 7327 7880 7336
rect 7828 7293 7837 7327
rect 7837 7293 7871 7327
rect 7871 7293 7880 7327
rect 7828 7284 7880 7293
rect 12980 7327 13032 7336
rect 12980 7293 13014 7327
rect 13014 7293 13032 7327
rect 12980 7284 13032 7293
rect 15188 7327 15240 7336
rect 15188 7293 15197 7327
rect 15197 7293 15231 7327
rect 15231 7293 15240 7327
rect 15188 7284 15240 7293
rect 20064 7284 20116 7336
rect 20892 7284 20944 7336
rect 8012 7216 8064 7268
rect 10312 7259 10364 7268
rect 10312 7225 10321 7259
rect 10321 7225 10355 7259
rect 10355 7225 10364 7259
rect 10312 7216 10364 7225
rect 9208 7148 9260 7200
rect 10680 7148 10732 7200
rect 10772 7148 10824 7200
rect 14544 7148 14596 7200
rect 17120 7148 17172 7200
rect 19972 7216 20024 7268
rect 22916 7284 22968 7336
rect 25676 7284 25728 7336
rect 17672 7148 17724 7200
rect 18132 7191 18184 7200
rect 18132 7157 18141 7191
rect 18141 7157 18175 7191
rect 18175 7157 18184 7191
rect 18868 7191 18920 7200
rect 18132 7148 18184 7157
rect 18868 7157 18877 7191
rect 18877 7157 18911 7191
rect 18911 7157 18920 7191
rect 18868 7148 18920 7157
rect 21260 7191 21312 7200
rect 21260 7157 21269 7191
rect 21269 7157 21303 7191
rect 21303 7157 21312 7191
rect 21260 7148 21312 7157
rect 21536 7148 21588 7200
rect 22180 7148 22232 7200
rect 23468 7191 23520 7200
rect 23468 7157 23477 7191
rect 23477 7157 23511 7191
rect 23511 7157 23520 7191
rect 23468 7148 23520 7157
rect 23836 7191 23888 7200
rect 23836 7157 23845 7191
rect 23845 7157 23879 7191
rect 23879 7157 23888 7191
rect 23836 7148 23888 7157
rect 23928 7191 23980 7200
rect 23928 7157 23937 7191
rect 23937 7157 23971 7191
rect 23971 7157 23980 7191
rect 25216 7191 25268 7200
rect 23928 7148 23980 7157
rect 25216 7157 25225 7191
rect 25225 7157 25259 7191
rect 25259 7157 25268 7191
rect 25216 7148 25268 7157
rect 10027 7046 10079 7098
rect 10091 7046 10143 7098
rect 10155 7046 10207 7098
rect 10219 7046 10271 7098
rect 19360 7046 19412 7098
rect 19424 7046 19476 7098
rect 19488 7046 19540 7098
rect 19552 7046 19604 7098
rect 9760 6987 9812 6996
rect 9760 6953 9769 6987
rect 9769 6953 9803 6987
rect 9803 6953 9812 6987
rect 9760 6944 9812 6953
rect 7828 6876 7880 6928
rect 10680 6876 10732 6928
rect 12980 6944 13032 6996
rect 14268 6944 14320 6996
rect 15556 6944 15608 6996
rect 17764 6944 17816 6996
rect 19236 6987 19288 6996
rect 19236 6953 19245 6987
rect 19245 6953 19279 6987
rect 19279 6953 19288 6987
rect 19236 6944 19288 6953
rect 20156 6944 20208 6996
rect 21260 6944 21312 6996
rect 23836 6944 23888 6996
rect 12060 6876 12112 6928
rect 16108 6876 16160 6928
rect 18868 6876 18920 6928
rect 21812 6876 21864 6928
rect 6908 6808 6960 6860
rect 8196 6808 8248 6860
rect 10772 6808 10824 6860
rect 11324 6851 11376 6860
rect 11324 6817 11333 6851
rect 11333 6817 11367 6851
rect 11367 6817 11376 6851
rect 11324 6808 11376 6817
rect 11416 6851 11468 6860
rect 11416 6817 11425 6851
rect 11425 6817 11459 6851
rect 11459 6817 11468 6851
rect 11692 6851 11744 6860
rect 11416 6808 11468 6817
rect 11692 6817 11726 6851
rect 11726 6817 11744 6851
rect 11692 6808 11744 6817
rect 15832 6808 15884 6860
rect 16476 6808 16528 6860
rect 20984 6851 21036 6860
rect 20984 6817 20993 6851
rect 20993 6817 21027 6851
rect 21027 6817 21036 6851
rect 20984 6808 21036 6817
rect 21904 6808 21956 6860
rect 22548 6851 22600 6860
rect 22548 6817 22571 6851
rect 22571 6817 22600 6851
rect 22548 6808 22600 6817
rect 24572 6808 24624 6860
rect 9668 6740 9720 6792
rect 13900 6783 13952 6792
rect 9392 6715 9444 6724
rect 9392 6681 9401 6715
rect 9401 6681 9435 6715
rect 9435 6681 9444 6715
rect 9392 6672 9444 6681
rect 9576 6672 9628 6724
rect 13900 6749 13909 6783
rect 13909 6749 13943 6783
rect 13943 6749 13952 6783
rect 13900 6740 13952 6749
rect 14544 6740 14596 6792
rect 15372 6715 15424 6724
rect 15372 6681 15381 6715
rect 15381 6681 15415 6715
rect 15415 6681 15424 6715
rect 15372 6672 15424 6681
rect 15464 6672 15516 6724
rect 13624 6604 13676 6656
rect 13808 6604 13860 6656
rect 18316 6740 18368 6792
rect 18592 6740 18644 6792
rect 17856 6672 17908 6724
rect 18776 6672 18828 6724
rect 17120 6604 17172 6656
rect 18684 6647 18736 6656
rect 18684 6613 18693 6647
rect 18693 6613 18727 6647
rect 18727 6613 18736 6647
rect 19420 6783 19472 6792
rect 19420 6749 19429 6783
rect 19429 6749 19463 6783
rect 19463 6749 19472 6783
rect 19420 6740 19472 6749
rect 20892 6740 20944 6792
rect 20340 6672 20392 6724
rect 22088 6740 22140 6792
rect 23376 6672 23428 6724
rect 24020 6672 24072 6724
rect 24848 6672 24900 6724
rect 21812 6647 21864 6656
rect 18684 6604 18736 6613
rect 21812 6613 21821 6647
rect 21821 6613 21855 6647
rect 21855 6613 21864 6647
rect 21812 6604 21864 6613
rect 22180 6647 22232 6656
rect 22180 6613 22189 6647
rect 22189 6613 22223 6647
rect 22223 6613 22232 6647
rect 22180 6604 22232 6613
rect 23652 6647 23704 6656
rect 23652 6613 23661 6647
rect 23661 6613 23695 6647
rect 23695 6613 23704 6647
rect 23652 6604 23704 6613
rect 24940 6647 24992 6656
rect 24940 6613 24949 6647
rect 24949 6613 24983 6647
rect 24983 6613 24992 6647
rect 24940 6604 24992 6613
rect 5360 6502 5412 6554
rect 5424 6502 5476 6554
rect 5488 6502 5540 6554
rect 5552 6502 5604 6554
rect 14694 6502 14746 6554
rect 14758 6502 14810 6554
rect 14822 6502 14874 6554
rect 14886 6502 14938 6554
rect 24027 6502 24079 6554
rect 24091 6502 24143 6554
rect 24155 6502 24207 6554
rect 24219 6502 24271 6554
rect 6908 6443 6960 6452
rect 6908 6409 6917 6443
rect 6917 6409 6951 6443
rect 6951 6409 6960 6443
rect 6908 6400 6960 6409
rect 9760 6400 9812 6452
rect 12244 6443 12296 6452
rect 12244 6409 12253 6443
rect 12253 6409 12287 6443
rect 12287 6409 12296 6443
rect 12244 6400 12296 6409
rect 12888 6307 12940 6316
rect 12888 6273 12897 6307
rect 12897 6273 12931 6307
rect 12931 6273 12940 6307
rect 12888 6264 12940 6273
rect 7828 6196 7880 6248
rect 8104 6239 8156 6248
rect 8104 6205 8113 6239
rect 8113 6205 8147 6239
rect 8147 6205 8156 6239
rect 8104 6196 8156 6205
rect 9208 6196 9260 6248
rect 13808 6239 13860 6248
rect 13808 6205 13817 6239
rect 13817 6205 13851 6239
rect 13851 6205 13860 6239
rect 13808 6196 13860 6205
rect 15832 6239 15884 6248
rect 15832 6205 15841 6239
rect 15841 6205 15875 6239
rect 15875 6205 15884 6239
rect 15832 6196 15884 6205
rect 17304 6400 17356 6452
rect 18500 6443 18552 6452
rect 18500 6409 18509 6443
rect 18509 6409 18543 6443
rect 18543 6409 18552 6443
rect 18500 6400 18552 6409
rect 20340 6443 20392 6452
rect 20340 6409 20349 6443
rect 20349 6409 20383 6443
rect 20383 6409 20392 6443
rect 20340 6400 20392 6409
rect 20892 6443 20944 6452
rect 20892 6409 20901 6443
rect 20901 6409 20935 6443
rect 20935 6409 20944 6443
rect 20892 6400 20944 6409
rect 21536 6443 21588 6452
rect 21536 6409 21545 6443
rect 21545 6409 21579 6443
rect 21579 6409 21588 6443
rect 21536 6400 21588 6409
rect 21720 6443 21772 6452
rect 21720 6409 21729 6443
rect 21729 6409 21763 6443
rect 21763 6409 21772 6443
rect 21720 6400 21772 6409
rect 22548 6400 22600 6452
rect 24572 6400 24624 6452
rect 24848 6375 24900 6384
rect 24848 6341 24857 6375
rect 24857 6341 24891 6375
rect 24891 6341 24900 6375
rect 24848 6332 24900 6341
rect 22180 6264 22232 6316
rect 18500 6196 18552 6248
rect 18960 6239 19012 6248
rect 9300 6128 9352 6180
rect 9392 6128 9444 6180
rect 9668 6128 9720 6180
rect 16660 6128 16712 6180
rect 17488 6171 17540 6180
rect 17488 6137 17497 6171
rect 17497 6137 17531 6171
rect 17531 6137 17540 6171
rect 17488 6128 17540 6137
rect 18960 6205 18969 6239
rect 18969 6205 19003 6239
rect 19003 6205 19012 6239
rect 18960 6196 19012 6205
rect 9484 6103 9536 6112
rect 9484 6069 9493 6103
rect 9493 6069 9527 6103
rect 9527 6069 9536 6103
rect 9484 6060 9536 6069
rect 11048 6103 11100 6112
rect 11048 6069 11057 6103
rect 11057 6069 11091 6103
rect 11091 6069 11100 6103
rect 11048 6060 11100 6069
rect 11508 6103 11560 6112
rect 11508 6069 11517 6103
rect 11517 6069 11551 6103
rect 11551 6069 11560 6103
rect 11508 6060 11560 6069
rect 12612 6103 12664 6112
rect 12612 6069 12621 6103
rect 12621 6069 12655 6103
rect 12655 6069 12664 6103
rect 12612 6060 12664 6069
rect 12704 6103 12756 6112
rect 12704 6069 12713 6103
rect 12713 6069 12747 6103
rect 12747 6069 12756 6103
rect 13624 6103 13676 6112
rect 12704 6060 12756 6069
rect 13624 6069 13633 6103
rect 13633 6069 13667 6103
rect 13667 6069 13676 6103
rect 13624 6060 13676 6069
rect 16108 6103 16160 6112
rect 16108 6069 16117 6103
rect 16117 6069 16151 6103
rect 16151 6069 16160 6103
rect 16108 6060 16160 6069
rect 16752 6103 16804 6112
rect 16752 6069 16761 6103
rect 16761 6069 16795 6103
rect 16795 6069 16804 6103
rect 16752 6060 16804 6069
rect 17120 6060 17172 6112
rect 19052 6128 19104 6180
rect 19420 6128 19472 6180
rect 21812 6128 21864 6180
rect 22272 6128 22324 6180
rect 23284 6196 23336 6248
rect 23652 6128 23704 6180
rect 18040 6103 18092 6112
rect 18040 6069 18049 6103
rect 18049 6069 18083 6103
rect 18083 6069 18092 6103
rect 18040 6060 18092 6069
rect 21536 6060 21588 6112
rect 22180 6103 22232 6112
rect 22180 6069 22189 6103
rect 22189 6069 22223 6103
rect 22223 6069 22232 6103
rect 22180 6060 22232 6069
rect 23100 6103 23152 6112
rect 23100 6069 23109 6103
rect 23109 6069 23143 6103
rect 23143 6069 23152 6103
rect 23100 6060 23152 6069
rect 25952 6060 26004 6112
rect 10027 5958 10079 6010
rect 10091 5958 10143 6010
rect 10155 5958 10207 6010
rect 10219 5958 10271 6010
rect 19360 5958 19412 6010
rect 19424 5958 19476 6010
rect 19488 5958 19540 6010
rect 19552 5958 19604 6010
rect 6908 5856 6960 5908
rect 9116 5856 9168 5908
rect 9484 5856 9536 5908
rect 9576 5899 9628 5908
rect 9576 5865 9585 5899
rect 9585 5865 9619 5899
rect 9619 5865 9628 5899
rect 9852 5899 9904 5908
rect 9576 5856 9628 5865
rect 9852 5865 9861 5899
rect 9861 5865 9895 5899
rect 9895 5865 9904 5899
rect 9852 5856 9904 5865
rect 9668 5788 9720 5840
rect 11048 5856 11100 5908
rect 12612 5856 12664 5908
rect 14544 5856 14596 5908
rect 15556 5899 15608 5908
rect 15556 5865 15565 5899
rect 15565 5865 15599 5899
rect 15599 5865 15608 5899
rect 15556 5856 15608 5865
rect 17580 5856 17632 5908
rect 19052 5856 19104 5908
rect 19880 5899 19932 5908
rect 19880 5865 19889 5899
rect 19889 5865 19923 5899
rect 19923 5865 19932 5899
rect 19880 5856 19932 5865
rect 21444 5856 21496 5908
rect 23376 5856 23428 5908
rect 11324 5831 11376 5840
rect 11324 5797 11333 5831
rect 11333 5797 11367 5831
rect 11367 5797 11376 5831
rect 11324 5788 11376 5797
rect 12060 5788 12112 5840
rect 17856 5831 17908 5840
rect 17856 5797 17890 5831
rect 17890 5797 17908 5831
rect 17856 5788 17908 5797
rect 20340 5788 20392 5840
rect 23652 5788 23704 5840
rect 8012 5720 8064 5772
rect 9300 5720 9352 5772
rect 9852 5720 9904 5772
rect 7920 5652 7972 5704
rect 8196 5695 8248 5704
rect 8196 5661 8205 5695
rect 8205 5661 8239 5695
rect 8239 5661 8248 5695
rect 8196 5652 8248 5661
rect 10312 5695 10364 5704
rect 7736 5627 7788 5636
rect 7736 5593 7745 5627
rect 7745 5593 7779 5627
rect 7779 5593 7788 5627
rect 7736 5584 7788 5593
rect 7828 5584 7880 5636
rect 10312 5661 10321 5695
rect 10321 5661 10355 5695
rect 10355 5661 10364 5695
rect 10312 5652 10364 5661
rect 11048 5720 11100 5772
rect 15004 5763 15056 5772
rect 15004 5729 15013 5763
rect 15013 5729 15047 5763
rect 15047 5729 15056 5763
rect 15004 5720 15056 5729
rect 16384 5763 16436 5772
rect 16384 5729 16393 5763
rect 16393 5729 16427 5763
rect 16427 5729 16436 5763
rect 16384 5720 16436 5729
rect 17304 5720 17356 5772
rect 22088 5720 22140 5772
rect 11416 5695 11468 5704
rect 11416 5661 11425 5695
rect 11425 5661 11459 5695
rect 11459 5661 11468 5695
rect 11416 5652 11468 5661
rect 16476 5695 16528 5704
rect 16476 5661 16485 5695
rect 16485 5661 16519 5695
rect 16519 5661 16528 5695
rect 16476 5652 16528 5661
rect 16568 5695 16620 5704
rect 16568 5661 16577 5695
rect 16577 5661 16611 5695
rect 16611 5661 16620 5695
rect 16568 5652 16620 5661
rect 17120 5652 17172 5704
rect 20616 5695 20668 5704
rect 20616 5661 20625 5695
rect 20625 5661 20659 5695
rect 20659 5661 20668 5695
rect 20616 5652 20668 5661
rect 22548 5695 22600 5704
rect 22548 5661 22557 5695
rect 22557 5661 22591 5695
rect 22591 5661 22600 5695
rect 22548 5652 22600 5661
rect 23284 5652 23336 5704
rect 11048 5516 11100 5568
rect 12612 5584 12664 5636
rect 13808 5584 13860 5636
rect 14176 5584 14228 5636
rect 17764 5516 17816 5568
rect 20984 5516 21036 5568
rect 21536 5516 21588 5568
rect 22916 5559 22968 5568
rect 22916 5525 22925 5559
rect 22925 5525 22959 5559
rect 22959 5525 22968 5559
rect 22916 5516 22968 5525
rect 24480 5516 24532 5568
rect 5360 5414 5412 5466
rect 5424 5414 5476 5466
rect 5488 5414 5540 5466
rect 5552 5414 5604 5466
rect 14694 5414 14746 5466
rect 14758 5414 14810 5466
rect 14822 5414 14874 5466
rect 14886 5414 14938 5466
rect 24027 5414 24079 5466
rect 24091 5414 24143 5466
rect 24155 5414 24207 5466
rect 24219 5414 24271 5466
rect 7920 5312 7972 5364
rect 9392 5312 9444 5364
rect 9668 5355 9720 5364
rect 9668 5321 9677 5355
rect 9677 5321 9711 5355
rect 9711 5321 9720 5355
rect 9668 5312 9720 5321
rect 10312 5312 10364 5364
rect 7644 5176 7696 5228
rect 9116 5219 9168 5228
rect 9116 5185 9125 5219
rect 9125 5185 9159 5219
rect 9159 5185 9168 5219
rect 9116 5176 9168 5185
rect 11048 5219 11100 5228
rect 11048 5185 11057 5219
rect 11057 5185 11091 5219
rect 11091 5185 11100 5219
rect 14176 5355 14228 5364
rect 14176 5321 14185 5355
rect 14185 5321 14219 5355
rect 14219 5321 14228 5355
rect 14176 5312 14228 5321
rect 17304 5312 17356 5364
rect 17488 5355 17540 5364
rect 17488 5321 17497 5355
rect 17497 5321 17531 5355
rect 17531 5321 17540 5355
rect 17488 5312 17540 5321
rect 18684 5312 18736 5364
rect 19052 5312 19104 5364
rect 17856 5244 17908 5296
rect 11048 5176 11100 5185
rect 11324 5108 11376 5160
rect 14176 5176 14228 5228
rect 17764 5176 17816 5228
rect 18316 5219 18368 5228
rect 18316 5185 18325 5219
rect 18325 5185 18359 5219
rect 18359 5185 18368 5219
rect 20340 5312 20392 5364
rect 22456 5312 22508 5364
rect 23560 5355 23612 5364
rect 23560 5321 23569 5355
rect 23569 5321 23603 5355
rect 23603 5321 23612 5355
rect 23560 5312 23612 5321
rect 24388 5312 24440 5364
rect 18316 5176 18368 5185
rect 20248 5176 20300 5228
rect 20616 5176 20668 5228
rect 10956 5083 11008 5092
rect 10956 5049 10965 5083
rect 10965 5049 10999 5083
rect 10999 5049 11008 5083
rect 10956 5040 11008 5049
rect 12888 5108 12940 5160
rect 14360 5108 14412 5160
rect 17672 5108 17724 5160
rect 19512 5151 19564 5160
rect 19512 5117 19521 5151
rect 19521 5117 19555 5151
rect 19555 5117 19564 5151
rect 19512 5108 19564 5117
rect 19880 5108 19932 5160
rect 21444 5108 21496 5160
rect 23468 5176 23520 5228
rect 23560 5108 23612 5160
rect 24480 5176 24532 5228
rect 12612 5040 12664 5092
rect 15280 5040 15332 5092
rect 16660 5040 16712 5092
rect 16844 5040 16896 5092
rect 19144 5040 19196 5092
rect 20064 5040 20116 5092
rect 23192 5040 23244 5092
rect 8012 5015 8064 5024
rect 8012 4981 8021 5015
rect 8021 4981 8055 5015
rect 8055 4981 8064 5015
rect 8012 4972 8064 4981
rect 8380 5015 8432 5024
rect 8380 4981 8389 5015
rect 8389 4981 8423 5015
rect 8423 4981 8432 5015
rect 8380 4972 8432 4981
rect 9300 4972 9352 5024
rect 9760 4972 9812 5024
rect 14544 4972 14596 5024
rect 16568 5015 16620 5024
rect 16568 4981 16577 5015
rect 16577 4981 16611 5015
rect 16611 4981 16620 5015
rect 16568 4972 16620 4981
rect 19236 5015 19288 5024
rect 19236 4981 19245 5015
rect 19245 4981 19279 5015
rect 19279 4981 19288 5015
rect 19236 4972 19288 4981
rect 19880 5015 19932 5024
rect 19880 4981 19889 5015
rect 19889 4981 19923 5015
rect 19923 4981 19932 5015
rect 19880 4972 19932 4981
rect 23652 4972 23704 5024
rect 25308 5015 25360 5024
rect 25308 4981 25317 5015
rect 25317 4981 25351 5015
rect 25351 4981 25360 5015
rect 25308 4972 25360 4981
rect 25952 4972 26004 5024
rect 10027 4870 10079 4922
rect 10091 4870 10143 4922
rect 10155 4870 10207 4922
rect 10219 4870 10271 4922
rect 19360 4870 19412 4922
rect 19424 4870 19476 4922
rect 19488 4870 19540 4922
rect 19552 4870 19604 4922
rect 7828 4811 7880 4820
rect 7828 4777 7837 4811
rect 7837 4777 7871 4811
rect 7871 4777 7880 4811
rect 7828 4768 7880 4777
rect 8104 4811 8156 4820
rect 8104 4777 8113 4811
rect 8113 4777 8147 4811
rect 8147 4777 8156 4811
rect 8104 4768 8156 4777
rect 9852 4811 9904 4820
rect 9852 4777 9861 4811
rect 9861 4777 9895 4811
rect 9895 4777 9904 4811
rect 9852 4768 9904 4777
rect 11508 4811 11560 4820
rect 11508 4777 11517 4811
rect 11517 4777 11551 4811
rect 11551 4777 11560 4811
rect 11508 4768 11560 4777
rect 12704 4768 12756 4820
rect 14176 4768 14228 4820
rect 15280 4811 15332 4820
rect 15280 4777 15289 4811
rect 15289 4777 15323 4811
rect 15323 4777 15332 4811
rect 15280 4768 15332 4777
rect 15648 4811 15700 4820
rect 15648 4777 15657 4811
rect 15657 4777 15691 4811
rect 15691 4777 15700 4811
rect 15648 4768 15700 4777
rect 10680 4632 10732 4684
rect 12060 4632 12112 4684
rect 14544 4700 14596 4752
rect 15004 4700 15056 4752
rect 16200 4768 16252 4820
rect 17212 4811 17264 4820
rect 17212 4777 17221 4811
rect 17221 4777 17255 4811
rect 17255 4777 17264 4811
rect 17212 4768 17264 4777
rect 18316 4811 18368 4820
rect 18316 4777 18325 4811
rect 18325 4777 18359 4811
rect 18359 4777 18368 4811
rect 18316 4768 18368 4777
rect 17488 4700 17540 4752
rect 17672 4743 17724 4752
rect 17672 4709 17681 4743
rect 17681 4709 17715 4743
rect 17715 4709 17724 4743
rect 18960 4768 19012 4820
rect 17672 4700 17724 4709
rect 18592 4700 18644 4752
rect 19236 4700 19288 4752
rect 20340 4768 20392 4820
rect 22088 4811 22140 4820
rect 22088 4777 22097 4811
rect 22097 4777 22131 4811
rect 22131 4777 22140 4811
rect 22088 4768 22140 4777
rect 23192 4811 23244 4820
rect 23192 4777 23201 4811
rect 23201 4777 23235 4811
rect 23235 4777 23244 4811
rect 23192 4768 23244 4777
rect 23376 4768 23428 4820
rect 24664 4768 24716 4820
rect 19972 4700 20024 4752
rect 22272 4700 22324 4752
rect 25032 4700 25084 4752
rect 13532 4632 13584 4684
rect 16384 4632 16436 4684
rect 17120 4632 17172 4684
rect 21996 4675 22048 4684
rect 8288 4607 8340 4616
rect 8288 4573 8297 4607
rect 8297 4573 8331 4607
rect 8331 4573 8340 4607
rect 8288 4564 8340 4573
rect 10128 4607 10180 4616
rect 10128 4573 10137 4607
rect 10137 4573 10171 4607
rect 10171 4573 10180 4607
rect 10128 4564 10180 4573
rect 13808 4607 13860 4616
rect 13808 4573 13817 4607
rect 13817 4573 13851 4607
rect 13851 4573 13860 4607
rect 13808 4564 13860 4573
rect 9300 4496 9352 4548
rect 12796 4496 12848 4548
rect 13624 4496 13676 4548
rect 14084 4564 14136 4616
rect 16568 4564 16620 4616
rect 17488 4564 17540 4616
rect 16476 4496 16528 4548
rect 19144 4564 19196 4616
rect 21996 4641 22005 4675
rect 22005 4641 22039 4675
rect 22039 4641 22048 4675
rect 21996 4632 22048 4641
rect 24756 4675 24808 4684
rect 24756 4641 24765 4675
rect 24765 4641 24799 4675
rect 24799 4641 24808 4675
rect 24756 4632 24808 4641
rect 20616 4607 20668 4616
rect 20616 4573 20625 4607
rect 20625 4573 20659 4607
rect 20659 4573 20668 4607
rect 20616 4564 20668 4573
rect 22272 4607 22324 4616
rect 22272 4573 22281 4607
rect 22281 4573 22315 4607
rect 22315 4573 22324 4607
rect 22272 4564 22324 4573
rect 19052 4496 19104 4548
rect 23744 4607 23796 4616
rect 23744 4573 23753 4607
rect 23753 4573 23787 4607
rect 23787 4573 23796 4607
rect 23744 4564 23796 4573
rect 9668 4428 9720 4480
rect 12612 4471 12664 4480
rect 12612 4437 12621 4471
rect 12621 4437 12655 4471
rect 12655 4437 12664 4471
rect 12612 4428 12664 4437
rect 12704 4471 12756 4480
rect 12704 4437 12713 4471
rect 12713 4437 12747 4471
rect 12747 4437 12756 4471
rect 18592 4471 18644 4480
rect 12704 4428 12756 4437
rect 18592 4437 18601 4471
rect 18601 4437 18635 4471
rect 18635 4437 18644 4471
rect 18592 4428 18644 4437
rect 18776 4471 18828 4480
rect 18776 4437 18785 4471
rect 18785 4437 18819 4471
rect 18819 4437 18828 4471
rect 18776 4428 18828 4437
rect 21536 4428 21588 4480
rect 22640 4471 22692 4480
rect 22640 4437 22649 4471
rect 22649 4437 22683 4471
rect 22683 4437 22692 4471
rect 22640 4428 22692 4437
rect 22916 4428 22968 4480
rect 23192 4428 23244 4480
rect 24664 4471 24716 4480
rect 24664 4437 24673 4471
rect 24673 4437 24707 4471
rect 24707 4437 24716 4471
rect 24664 4428 24716 4437
rect 5360 4326 5412 4378
rect 5424 4326 5476 4378
rect 5488 4326 5540 4378
rect 5552 4326 5604 4378
rect 14694 4326 14746 4378
rect 14758 4326 14810 4378
rect 14822 4326 14874 4378
rect 14886 4326 14938 4378
rect 24027 4326 24079 4378
rect 24091 4326 24143 4378
rect 24155 4326 24207 4378
rect 24219 4326 24271 4378
rect 14084 4224 14136 4276
rect 7644 4088 7696 4140
rect 10680 4156 10732 4208
rect 9668 4131 9720 4140
rect 9668 4097 9677 4131
rect 9677 4097 9711 4131
rect 9711 4097 9720 4131
rect 9668 4088 9720 4097
rect 11600 4131 11652 4140
rect 8932 4020 8984 4072
rect 11600 4097 11609 4131
rect 11609 4097 11643 4131
rect 11643 4097 11652 4131
rect 11600 4088 11652 4097
rect 12796 4131 12848 4140
rect 12796 4097 12805 4131
rect 12805 4097 12839 4131
rect 12839 4097 12848 4131
rect 12796 4088 12848 4097
rect 11876 4063 11928 4072
rect 11876 4029 11885 4063
rect 11885 4029 11919 4063
rect 11919 4029 11928 4063
rect 11876 4020 11928 4029
rect 12704 4020 12756 4072
rect 13900 4063 13952 4072
rect 13900 4029 13909 4063
rect 13909 4029 13943 4063
rect 13943 4029 13952 4063
rect 13900 4020 13952 4029
rect 13992 4020 14044 4072
rect 16568 4224 16620 4276
rect 21996 4224 22048 4276
rect 23376 4224 23428 4276
rect 23928 4267 23980 4276
rect 23928 4233 23937 4267
rect 23937 4233 23971 4267
rect 23971 4233 23980 4267
rect 23928 4224 23980 4233
rect 24756 4224 24808 4276
rect 16292 4131 16344 4140
rect 16292 4097 16301 4131
rect 16301 4097 16335 4131
rect 16335 4097 16344 4131
rect 16292 4088 16344 4097
rect 17304 4088 17356 4140
rect 18592 4088 18644 4140
rect 18960 4088 19012 4140
rect 20340 4156 20392 4208
rect 22272 4156 22324 4208
rect 23100 4156 23152 4208
rect 20708 4131 20760 4140
rect 20708 4097 20717 4131
rect 20717 4097 20751 4131
rect 20751 4097 20760 4131
rect 20708 4088 20760 4097
rect 23284 4088 23336 4140
rect 24664 4156 24716 4208
rect 7552 3927 7604 3936
rect 7552 3893 7561 3927
rect 7561 3893 7595 3927
rect 7595 3893 7604 3927
rect 7552 3884 7604 3893
rect 8656 3927 8708 3936
rect 8656 3893 8665 3927
rect 8665 3893 8699 3927
rect 8699 3893 8708 3927
rect 8656 3884 8708 3893
rect 8932 3927 8984 3936
rect 8932 3893 8941 3927
rect 8941 3893 8975 3927
rect 8975 3893 8984 3927
rect 8932 3884 8984 3893
rect 9392 3952 9444 4004
rect 10128 3952 10180 4004
rect 11324 3952 11376 4004
rect 20892 4020 20944 4072
rect 18132 3995 18184 4004
rect 18132 3961 18141 3995
rect 18141 3961 18175 3995
rect 18175 3961 18184 3995
rect 18132 3952 18184 3961
rect 19236 3952 19288 4004
rect 24480 4020 24532 4072
rect 21720 3952 21772 4004
rect 24572 3952 24624 4004
rect 9300 3884 9352 3936
rect 9576 3927 9628 3936
rect 9576 3893 9585 3927
rect 9585 3893 9619 3927
rect 9619 3893 9628 3927
rect 9576 3884 9628 3893
rect 11140 3927 11192 3936
rect 11140 3893 11149 3927
rect 11149 3893 11183 3927
rect 11183 3893 11192 3927
rect 11140 3884 11192 3893
rect 12152 3927 12204 3936
rect 12152 3893 12161 3927
rect 12161 3893 12195 3927
rect 12195 3893 12204 3927
rect 12612 3927 12664 3936
rect 12152 3884 12204 3893
rect 12612 3893 12621 3927
rect 12621 3893 12655 3927
rect 12655 3893 12664 3927
rect 12612 3884 12664 3893
rect 13348 3927 13400 3936
rect 13348 3893 13357 3927
rect 13357 3893 13391 3927
rect 13391 3893 13400 3927
rect 13348 3884 13400 3893
rect 13808 3927 13860 3936
rect 13808 3893 13817 3927
rect 13817 3893 13851 3927
rect 13851 3893 13860 3927
rect 13808 3884 13860 3893
rect 15464 3884 15516 3936
rect 16200 3884 16252 3936
rect 17120 3927 17172 3936
rect 17120 3893 17129 3927
rect 17129 3893 17163 3927
rect 17163 3893 17172 3927
rect 17120 3884 17172 3893
rect 17488 3927 17540 3936
rect 17488 3893 17497 3927
rect 17497 3893 17531 3927
rect 17531 3893 17540 3927
rect 17488 3884 17540 3893
rect 17764 3927 17816 3936
rect 17764 3893 17773 3927
rect 17773 3893 17807 3927
rect 17807 3893 17816 3927
rect 17764 3884 17816 3893
rect 19788 3884 19840 3936
rect 19972 3927 20024 3936
rect 19972 3893 19981 3927
rect 19981 3893 20015 3927
rect 20015 3893 20024 3927
rect 19972 3884 20024 3893
rect 20064 3927 20116 3936
rect 20064 3893 20073 3927
rect 20073 3893 20107 3927
rect 20107 3893 20116 3927
rect 21168 3927 21220 3936
rect 20064 3884 20116 3893
rect 21168 3893 21177 3927
rect 21177 3893 21211 3927
rect 21211 3893 21220 3927
rect 21168 3884 21220 3893
rect 21536 3927 21588 3936
rect 21536 3893 21545 3927
rect 21545 3893 21579 3927
rect 21579 3893 21588 3927
rect 21536 3884 21588 3893
rect 10027 3782 10079 3834
rect 10091 3782 10143 3834
rect 10155 3782 10207 3834
rect 10219 3782 10271 3834
rect 19360 3782 19412 3834
rect 19424 3782 19476 3834
rect 19488 3782 19540 3834
rect 19552 3782 19604 3834
rect 7644 3723 7696 3732
rect 7644 3689 7653 3723
rect 7653 3689 7687 3723
rect 7687 3689 7696 3723
rect 7644 3680 7696 3689
rect 10680 3680 10732 3732
rect 11324 3723 11376 3732
rect 11324 3689 11333 3723
rect 11333 3689 11367 3723
rect 11367 3689 11376 3723
rect 11324 3680 11376 3689
rect 12796 3680 12848 3732
rect 13992 3723 14044 3732
rect 13992 3689 14001 3723
rect 14001 3689 14035 3723
rect 14035 3689 14044 3723
rect 13992 3680 14044 3689
rect 14544 3680 14596 3732
rect 14820 3723 14872 3732
rect 14820 3689 14829 3723
rect 14829 3689 14863 3723
rect 14863 3689 14872 3723
rect 14820 3680 14872 3689
rect 16016 3723 16068 3732
rect 16016 3689 16025 3723
rect 16025 3689 16059 3723
rect 16059 3689 16068 3723
rect 16016 3680 16068 3689
rect 16384 3680 16436 3732
rect 17028 3723 17080 3732
rect 17028 3689 17037 3723
rect 17037 3689 17071 3723
rect 17071 3689 17080 3723
rect 17028 3680 17080 3689
rect 17672 3723 17724 3732
rect 17672 3689 17681 3723
rect 17681 3689 17715 3723
rect 17715 3689 17724 3723
rect 17672 3680 17724 3689
rect 18224 3680 18276 3732
rect 18776 3680 18828 3732
rect 21168 3723 21220 3732
rect 21168 3689 21177 3723
rect 21177 3689 21211 3723
rect 21211 3689 21220 3723
rect 21168 3680 21220 3689
rect 22088 3680 22140 3732
rect 23744 3680 23796 3732
rect 9300 3612 9352 3664
rect 9668 3655 9720 3664
rect 9668 3621 9702 3655
rect 9702 3621 9720 3655
rect 9668 3612 9720 3621
rect 8472 3544 8524 3596
rect 16844 3612 16896 3664
rect 17764 3612 17816 3664
rect 18960 3612 19012 3664
rect 19144 3655 19196 3664
rect 19144 3621 19153 3655
rect 19153 3621 19187 3655
rect 19187 3621 19196 3655
rect 19144 3612 19196 3621
rect 23560 3655 23612 3664
rect 23560 3621 23594 3655
rect 23594 3621 23612 3655
rect 23560 3612 23612 3621
rect 11968 3544 12020 3596
rect 12152 3587 12204 3596
rect 12152 3553 12186 3587
rect 12186 3553 12204 3587
rect 15372 3587 15424 3596
rect 12152 3544 12204 3553
rect 15372 3553 15381 3587
rect 15381 3553 15415 3587
rect 15415 3553 15424 3587
rect 15372 3544 15424 3553
rect 15464 3587 15516 3596
rect 15464 3553 15473 3587
rect 15473 3553 15507 3587
rect 15507 3553 15516 3587
rect 15464 3544 15516 3553
rect 16384 3544 16436 3596
rect 18132 3544 18184 3596
rect 22640 3587 22692 3596
rect 22640 3553 22649 3587
rect 22649 3553 22683 3587
rect 22683 3553 22692 3587
rect 22640 3544 22692 3553
rect 24572 3544 24624 3596
rect 9392 3519 9444 3528
rect 8564 3340 8616 3392
rect 8656 3340 8708 3392
rect 9392 3485 9401 3519
rect 9401 3485 9435 3519
rect 9435 3485 9444 3519
rect 15556 3519 15608 3528
rect 9392 3476 9444 3485
rect 15556 3485 15565 3519
rect 15565 3485 15599 3519
rect 15599 3485 15608 3519
rect 15556 3476 15608 3485
rect 17212 3519 17264 3528
rect 17212 3485 17221 3519
rect 17221 3485 17255 3519
rect 17255 3485 17264 3519
rect 17212 3476 17264 3485
rect 18684 3519 18736 3528
rect 18684 3485 18693 3519
rect 18693 3485 18727 3519
rect 18727 3485 18736 3519
rect 18684 3476 18736 3485
rect 21260 3519 21312 3528
rect 21260 3485 21269 3519
rect 21269 3485 21303 3519
rect 21303 3485 21312 3519
rect 21260 3476 21312 3485
rect 21352 3519 21404 3528
rect 21352 3485 21361 3519
rect 21361 3485 21395 3519
rect 21395 3485 21404 3519
rect 21352 3476 21404 3485
rect 9576 3340 9628 3392
rect 10496 3340 10548 3392
rect 12888 3340 12940 3392
rect 15004 3383 15056 3392
rect 15004 3349 15013 3383
rect 15013 3349 15047 3383
rect 15047 3349 15056 3383
rect 15004 3340 15056 3349
rect 17304 3340 17356 3392
rect 19144 3340 19196 3392
rect 19972 3340 20024 3392
rect 20800 3383 20852 3392
rect 20800 3349 20809 3383
rect 20809 3349 20843 3383
rect 20843 3349 20852 3383
rect 20800 3340 20852 3349
rect 24664 3383 24716 3392
rect 24664 3349 24673 3383
rect 24673 3349 24707 3383
rect 24707 3349 24716 3383
rect 24664 3340 24716 3349
rect 5360 3238 5412 3290
rect 5424 3238 5476 3290
rect 5488 3238 5540 3290
rect 5552 3238 5604 3290
rect 14694 3238 14746 3290
rect 14758 3238 14810 3290
rect 14822 3238 14874 3290
rect 14886 3238 14938 3290
rect 24027 3238 24079 3290
rect 24091 3238 24143 3290
rect 24155 3238 24207 3290
rect 24219 3238 24271 3290
rect 8656 3136 8708 3188
rect 8840 3179 8892 3188
rect 8840 3145 8849 3179
rect 8849 3145 8883 3179
rect 8883 3145 8892 3179
rect 8840 3136 8892 3145
rect 9668 3136 9720 3188
rect 12428 3179 12480 3188
rect 12428 3145 12437 3179
rect 12437 3145 12471 3179
rect 12471 3145 12480 3179
rect 12428 3136 12480 3145
rect 15556 3136 15608 3188
rect 16384 3179 16436 3188
rect 16384 3145 16393 3179
rect 16393 3145 16427 3179
rect 16427 3145 16436 3179
rect 16384 3136 16436 3145
rect 16844 3136 16896 3188
rect 18684 3136 18736 3188
rect 21260 3136 21312 3188
rect 23192 3179 23244 3188
rect 23192 3145 23201 3179
rect 23201 3145 23235 3179
rect 23235 3145 23244 3179
rect 23192 3136 23244 3145
rect 8472 3068 8524 3120
rect 8840 2932 8892 2984
rect 15096 3068 15148 3120
rect 17028 3111 17080 3120
rect 17028 3077 17037 3111
rect 17037 3077 17071 3111
rect 17071 3077 17080 3111
rect 17028 3068 17080 3077
rect 13072 3043 13124 3052
rect 13072 3009 13081 3043
rect 13081 3009 13115 3043
rect 13115 3009 13124 3043
rect 13072 3000 13124 3009
rect 13900 3000 13952 3052
rect 15372 3000 15424 3052
rect 20248 3043 20300 3052
rect 20248 3009 20257 3043
rect 20257 3009 20291 3043
rect 20291 3009 20300 3043
rect 20248 3000 20300 3009
rect 23560 3000 23612 3052
rect 23928 3043 23980 3052
rect 23928 3009 23937 3043
rect 23937 3009 23971 3043
rect 23971 3009 23980 3043
rect 23928 3000 23980 3009
rect 24664 3000 24716 3052
rect 10404 2932 10456 2984
rect 12152 2932 12204 2984
rect 13532 2932 13584 2984
rect 16016 2932 16068 2984
rect 17764 2975 17816 2984
rect 17764 2941 17773 2975
rect 17773 2941 17807 2975
rect 17807 2941 17816 2975
rect 17764 2932 17816 2941
rect 7184 2907 7236 2916
rect 7184 2873 7193 2907
rect 7193 2873 7227 2907
rect 7227 2873 7236 2907
rect 7184 2864 7236 2873
rect 11876 2907 11928 2916
rect 11876 2873 11885 2907
rect 11885 2873 11919 2907
rect 11919 2873 11928 2907
rect 11876 2864 11928 2873
rect 12888 2907 12940 2916
rect 12888 2873 12897 2907
rect 12897 2873 12931 2907
rect 12931 2873 12940 2907
rect 12888 2864 12940 2873
rect 14544 2864 14596 2916
rect 17304 2864 17356 2916
rect 19052 2864 19104 2916
rect 20248 2864 20300 2916
rect 21352 2932 21404 2984
rect 23468 2932 23520 2984
rect 23192 2864 23244 2916
rect 23836 2907 23888 2916
rect 23836 2873 23845 2907
rect 23845 2873 23879 2907
rect 23879 2873 23888 2907
rect 23836 2864 23888 2873
rect 24572 2864 24624 2916
rect 8656 2796 8708 2848
rect 10404 2796 10456 2848
rect 13716 2796 13768 2848
rect 21720 2796 21772 2848
rect 25124 2839 25176 2848
rect 25124 2805 25133 2839
rect 25133 2805 25167 2839
rect 25167 2805 25176 2839
rect 25124 2796 25176 2805
rect 25768 2796 25820 2848
rect 10027 2694 10079 2746
rect 10091 2694 10143 2746
rect 10155 2694 10207 2746
rect 10219 2694 10271 2746
rect 19360 2694 19412 2746
rect 19424 2694 19476 2746
rect 19488 2694 19540 2746
rect 19552 2694 19604 2746
rect 9300 2635 9352 2644
rect 9300 2601 9309 2635
rect 9309 2601 9343 2635
rect 9343 2601 9352 2635
rect 9300 2592 9352 2601
rect 10680 2635 10732 2644
rect 10680 2601 10689 2635
rect 10689 2601 10723 2635
rect 10723 2601 10732 2635
rect 10680 2592 10732 2601
rect 8196 2499 8248 2508
rect 8196 2465 8205 2499
rect 8205 2465 8239 2499
rect 8239 2465 8248 2499
rect 8196 2456 8248 2465
rect 10956 2524 11008 2576
rect 10404 2456 10456 2508
rect 10496 2456 10548 2508
rect 8288 2431 8340 2440
rect 8288 2397 8297 2431
rect 8297 2397 8331 2431
rect 8331 2397 8340 2431
rect 8288 2388 8340 2397
rect 8472 2431 8524 2440
rect 8472 2397 8481 2431
rect 8481 2397 8515 2431
rect 8515 2397 8524 2431
rect 8472 2388 8524 2397
rect 12060 2592 12112 2644
rect 13532 2592 13584 2644
rect 16568 2635 16620 2644
rect 16568 2601 16577 2635
rect 16577 2601 16611 2635
rect 16611 2601 16620 2635
rect 16568 2592 16620 2601
rect 17212 2635 17264 2644
rect 17212 2601 17221 2635
rect 17221 2601 17255 2635
rect 17255 2601 17264 2635
rect 17212 2592 17264 2601
rect 19052 2592 19104 2644
rect 20708 2635 20760 2644
rect 20708 2601 20717 2635
rect 20717 2601 20751 2635
rect 20751 2601 20760 2635
rect 20708 2592 20760 2601
rect 21352 2592 21404 2644
rect 23008 2592 23060 2644
rect 24204 2635 24256 2644
rect 24204 2601 24213 2635
rect 24213 2601 24247 2635
rect 24247 2601 24256 2635
rect 24204 2592 24256 2601
rect 25768 2635 25820 2644
rect 25768 2601 25777 2635
rect 25777 2601 25811 2635
rect 25811 2601 25820 2635
rect 25768 2592 25820 2601
rect 13072 2524 13124 2576
rect 15556 2524 15608 2576
rect 11968 2456 12020 2508
rect 13900 2456 13952 2508
rect 18316 2499 18368 2508
rect 18316 2465 18350 2499
rect 18350 2465 18368 2499
rect 18316 2456 18368 2465
rect 20432 2456 20484 2508
rect 21720 2456 21772 2508
rect 24112 2499 24164 2508
rect 17764 2388 17816 2440
rect 7828 2363 7880 2372
rect 7828 2329 7837 2363
rect 7837 2329 7871 2363
rect 7871 2329 7880 2363
rect 7828 2320 7880 2329
rect 24112 2465 24121 2499
rect 24121 2465 24155 2499
rect 24155 2465 24164 2499
rect 24112 2456 24164 2465
rect 24572 2388 24624 2440
rect 10404 2252 10456 2304
rect 10496 2295 10548 2304
rect 10496 2261 10505 2295
rect 10505 2261 10539 2295
rect 10539 2261 10548 2295
rect 20248 2295 20300 2304
rect 10496 2252 10548 2261
rect 20248 2261 20257 2295
rect 20257 2261 20291 2295
rect 20291 2261 20300 2295
rect 20248 2252 20300 2261
rect 23468 2295 23520 2304
rect 23468 2261 23477 2295
rect 23477 2261 23511 2295
rect 23511 2261 23520 2295
rect 23468 2252 23520 2261
rect 5360 2150 5412 2202
rect 5424 2150 5476 2202
rect 5488 2150 5540 2202
rect 5552 2150 5604 2202
rect 14694 2150 14746 2202
rect 14758 2150 14810 2202
rect 14822 2150 14874 2202
rect 14886 2150 14938 2202
rect 24027 2150 24079 2202
rect 24091 2150 24143 2202
rect 24155 2150 24207 2202
rect 24219 2150 24271 2202
rect 21628 1980 21680 2032
rect 24020 1980 24072 2032
rect 17488 552 17540 604
rect 18040 552 18092 604
rect 18132 552 18184 604
rect 18592 552 18644 604
rect 22088 552 22140 604
rect 25216 552 25268 604
rect 25952 552 26004 604
rect 26320 552 26372 604
<< metal2 >>
rect 2490 27520 2546 28000
rect 8010 27520 8066 28000
rect 13622 27520 13678 28000
rect 19234 27520 19290 28000
rect 24846 27520 24902 28000
rect 2504 23526 2532 27520
rect 5334 25052 5630 25072
rect 5390 25050 5414 25052
rect 5470 25050 5494 25052
rect 5550 25050 5574 25052
rect 5412 24998 5414 25050
rect 5476 24998 5488 25050
rect 5550 24998 5552 25050
rect 5390 24996 5414 24998
rect 5470 24996 5494 24998
rect 5550 24996 5574 24998
rect 5334 24976 5630 24996
rect 5334 23964 5630 23984
rect 5390 23962 5414 23964
rect 5470 23962 5494 23964
rect 5550 23962 5574 23964
rect 5412 23910 5414 23962
rect 5476 23910 5488 23962
rect 5550 23910 5552 23962
rect 5390 23908 5414 23910
rect 5470 23908 5494 23910
rect 5550 23908 5574 23910
rect 5334 23888 5630 23908
rect 2492 23520 2544 23526
rect 2492 23462 2544 23468
rect 3780 23520 3832 23526
rect 3780 23462 3832 23468
rect 3792 14521 3820 23462
rect 5334 22876 5630 22896
rect 5390 22874 5414 22876
rect 5470 22874 5494 22876
rect 5550 22874 5574 22876
rect 5412 22822 5414 22874
rect 5476 22822 5488 22874
rect 5550 22822 5552 22874
rect 5390 22820 5414 22822
rect 5470 22820 5494 22822
rect 5550 22820 5574 22822
rect 5334 22800 5630 22820
rect 5334 21788 5630 21808
rect 5390 21786 5414 21788
rect 5470 21786 5494 21788
rect 5550 21786 5574 21788
rect 5412 21734 5414 21786
rect 5476 21734 5488 21786
rect 5550 21734 5552 21786
rect 5390 21732 5414 21734
rect 5470 21732 5494 21734
rect 5550 21732 5574 21734
rect 5334 21712 5630 21732
rect 5334 20700 5630 20720
rect 5390 20698 5414 20700
rect 5470 20698 5494 20700
rect 5550 20698 5574 20700
rect 5412 20646 5414 20698
rect 5476 20646 5488 20698
rect 5550 20646 5552 20698
rect 5390 20644 5414 20646
rect 5470 20644 5494 20646
rect 5550 20644 5574 20646
rect 5334 20624 5630 20644
rect 5334 19612 5630 19632
rect 5390 19610 5414 19612
rect 5470 19610 5494 19612
rect 5550 19610 5574 19612
rect 5412 19558 5414 19610
rect 5476 19558 5488 19610
rect 5550 19558 5552 19610
rect 5390 19556 5414 19558
rect 5470 19556 5494 19558
rect 5550 19556 5574 19558
rect 5334 19536 5630 19556
rect 5334 18524 5630 18544
rect 5390 18522 5414 18524
rect 5470 18522 5494 18524
rect 5550 18522 5574 18524
rect 5412 18470 5414 18522
rect 5476 18470 5488 18522
rect 5550 18470 5552 18522
rect 5390 18468 5414 18470
rect 5470 18468 5494 18470
rect 5550 18468 5574 18470
rect 5334 18448 5630 18468
rect 5334 17436 5630 17456
rect 5390 17434 5414 17436
rect 5470 17434 5494 17436
rect 5550 17434 5574 17436
rect 5412 17382 5414 17434
rect 5476 17382 5488 17434
rect 5550 17382 5552 17434
rect 5390 17380 5414 17382
rect 5470 17380 5494 17382
rect 5550 17380 5574 17382
rect 5334 17360 5630 17380
rect 7550 16960 7606 16969
rect 7550 16895 7606 16904
rect 5334 16348 5630 16368
rect 5390 16346 5414 16348
rect 5470 16346 5494 16348
rect 5550 16346 5574 16348
rect 5412 16294 5414 16346
rect 5476 16294 5488 16346
rect 5550 16294 5552 16346
rect 5390 16292 5414 16294
rect 5470 16292 5494 16294
rect 5550 16292 5574 16294
rect 5334 16272 5630 16292
rect 5334 15260 5630 15280
rect 5390 15258 5414 15260
rect 5470 15258 5494 15260
rect 5550 15258 5574 15260
rect 5412 15206 5414 15258
rect 5476 15206 5488 15258
rect 5550 15206 5552 15258
rect 5390 15204 5414 15206
rect 5470 15204 5494 15206
rect 5550 15204 5574 15206
rect 5334 15184 5630 15204
rect 3778 14512 3834 14521
rect 3778 14447 3834 14456
rect 5334 14172 5630 14192
rect 5390 14170 5414 14172
rect 5470 14170 5494 14172
rect 5550 14170 5574 14172
rect 5412 14118 5414 14170
rect 5476 14118 5488 14170
rect 5550 14118 5552 14170
rect 5390 14116 5414 14118
rect 5470 14116 5494 14118
rect 5550 14116 5574 14118
rect 5334 14096 5630 14116
rect 5334 13084 5630 13104
rect 5390 13082 5414 13084
rect 5470 13082 5494 13084
rect 5550 13082 5574 13084
rect 5412 13030 5414 13082
rect 5476 13030 5488 13082
rect 5550 13030 5552 13082
rect 5390 13028 5414 13030
rect 5470 13028 5494 13030
rect 5550 13028 5574 13030
rect 5334 13008 5630 13028
rect 3870 12744 3926 12753
rect 3870 12679 3926 12688
rect 1294 8392 1350 8401
rect 1294 8327 1350 8336
rect 650 6352 706 6361
rect 650 6287 706 6296
rect 6 4176 62 4185
rect 6 4111 62 4120
rect 20 480 48 4111
rect 664 480 692 6287
rect 1308 480 1336 8327
rect 3884 7546 3912 12679
rect 5334 11996 5630 12016
rect 5390 11994 5414 11996
rect 5470 11994 5494 11996
rect 5550 11994 5574 11996
rect 5412 11942 5414 11994
rect 5476 11942 5488 11994
rect 5550 11942 5552 11994
rect 5390 11940 5414 11942
rect 5470 11940 5494 11942
rect 5550 11940 5574 11942
rect 5334 11920 5630 11940
rect 5334 10908 5630 10928
rect 5390 10906 5414 10908
rect 5470 10906 5494 10908
rect 5550 10906 5574 10908
rect 5412 10854 5414 10906
rect 5476 10854 5488 10906
rect 5550 10854 5552 10906
rect 5390 10852 5414 10854
rect 5470 10852 5494 10854
rect 5550 10852 5574 10854
rect 5334 10832 5630 10852
rect 5334 9820 5630 9840
rect 5390 9818 5414 9820
rect 5470 9818 5494 9820
rect 5550 9818 5574 9820
rect 5412 9766 5414 9818
rect 5476 9766 5488 9818
rect 5550 9766 5552 9818
rect 5390 9764 5414 9766
rect 5470 9764 5494 9766
rect 5550 9764 5574 9766
rect 5334 9744 5630 9764
rect 5802 9480 5858 9489
rect 5802 9415 5858 9424
rect 5334 8732 5630 8752
rect 5390 8730 5414 8732
rect 5470 8730 5494 8732
rect 5550 8730 5574 8732
rect 5412 8678 5414 8730
rect 5476 8678 5488 8730
rect 5550 8678 5552 8730
rect 5390 8676 5414 8678
rect 5470 8676 5494 8678
rect 5550 8676 5574 8678
rect 5334 8656 5630 8676
rect 5066 7984 5122 7993
rect 5066 7919 5122 7928
rect 3872 7540 3924 7546
rect 3872 7482 3924 7488
rect 1938 7304 1994 7313
rect 1938 7239 1994 7248
rect 1952 480 1980 7239
rect 4514 5264 4570 5273
rect 4514 5199 4570 5208
rect 3226 4176 3282 4185
rect 3226 4111 3282 4120
rect 2582 3904 2638 3913
rect 2582 3839 2638 3848
rect 2596 480 2624 3839
rect 3240 480 3268 4111
rect 3962 3496 4018 3505
rect 3962 3431 4018 3440
rect 3976 626 4004 3431
rect 3884 598 4004 626
rect 3884 480 3912 598
rect 4528 480 4556 5199
rect 5080 4457 5108 7919
rect 5334 7644 5630 7664
rect 5390 7642 5414 7644
rect 5470 7642 5494 7644
rect 5550 7642 5574 7644
rect 5412 7590 5414 7642
rect 5476 7590 5488 7642
rect 5550 7590 5552 7642
rect 5390 7588 5414 7590
rect 5470 7588 5494 7590
rect 5550 7588 5574 7590
rect 5334 7568 5630 7588
rect 5160 7540 5212 7546
rect 5160 7482 5212 7488
rect 5066 4448 5122 4457
rect 5066 4383 5122 4392
rect 5172 480 5200 7482
rect 5334 6556 5630 6576
rect 5390 6554 5414 6556
rect 5470 6554 5494 6556
rect 5550 6554 5574 6556
rect 5412 6502 5414 6554
rect 5476 6502 5488 6554
rect 5550 6502 5552 6554
rect 5390 6500 5414 6502
rect 5470 6500 5494 6502
rect 5550 6500 5574 6502
rect 5334 6480 5630 6500
rect 5334 5468 5630 5488
rect 5390 5466 5414 5468
rect 5470 5466 5494 5468
rect 5550 5466 5574 5468
rect 5412 5414 5414 5466
rect 5476 5414 5488 5466
rect 5550 5414 5552 5466
rect 5390 5412 5414 5414
rect 5470 5412 5494 5414
rect 5550 5412 5574 5414
rect 5334 5392 5630 5412
rect 5334 4380 5630 4400
rect 5390 4378 5414 4380
rect 5470 4378 5494 4380
rect 5550 4378 5574 4380
rect 5412 4326 5414 4378
rect 5476 4326 5488 4378
rect 5550 4326 5552 4378
rect 5390 4324 5414 4326
rect 5470 4324 5494 4326
rect 5550 4324 5574 4326
rect 5334 4304 5630 4324
rect 5334 3292 5630 3312
rect 5390 3290 5414 3292
rect 5470 3290 5494 3292
rect 5550 3290 5574 3292
rect 5412 3238 5414 3290
rect 5476 3238 5488 3290
rect 5550 3238 5552 3290
rect 5390 3236 5414 3238
rect 5470 3236 5494 3238
rect 5550 3236 5574 3238
rect 5334 3216 5630 3236
rect 5334 2204 5630 2224
rect 5390 2202 5414 2204
rect 5470 2202 5494 2204
rect 5550 2202 5574 2204
rect 5412 2150 5414 2202
rect 5476 2150 5488 2202
rect 5550 2150 5552 2202
rect 5390 2148 5414 2150
rect 5470 2148 5494 2150
rect 5550 2148 5574 2150
rect 5334 2128 5630 2148
rect 5816 480 5844 9415
rect 6908 6860 6960 6866
rect 6908 6802 6960 6808
rect 6920 6458 6948 6802
rect 6908 6452 6960 6458
rect 6908 6394 6960 6400
rect 6920 5914 6948 6394
rect 6908 5908 6960 5914
rect 6908 5850 6960 5856
rect 7090 4992 7146 5001
rect 7090 4927 7146 4936
rect 6446 4448 6502 4457
rect 6446 4383 6502 4392
rect 6460 480 6488 4383
rect 7104 480 7132 4927
rect 7564 3942 7592 16895
rect 7828 7744 7880 7750
rect 7828 7686 7880 7692
rect 7642 7576 7698 7585
rect 7642 7511 7698 7520
rect 7656 5234 7684 7511
rect 7840 7342 7868 7686
rect 8024 7546 8052 27520
rect 13636 27418 13664 27520
rect 13544 27390 13664 27418
rect 10001 25596 10297 25616
rect 10057 25594 10081 25596
rect 10137 25594 10161 25596
rect 10217 25594 10241 25596
rect 10079 25542 10081 25594
rect 10143 25542 10155 25594
rect 10217 25542 10219 25594
rect 10057 25540 10081 25542
rect 10137 25540 10161 25542
rect 10217 25540 10241 25542
rect 10001 25520 10297 25540
rect 10001 24508 10297 24528
rect 10057 24506 10081 24508
rect 10137 24506 10161 24508
rect 10217 24506 10241 24508
rect 10079 24454 10081 24506
rect 10143 24454 10155 24506
rect 10217 24454 10219 24506
rect 10057 24452 10081 24454
rect 10137 24452 10161 24454
rect 10217 24452 10241 24454
rect 10001 24432 10297 24452
rect 10678 23624 10734 23633
rect 10678 23559 10734 23568
rect 10001 23420 10297 23440
rect 10057 23418 10081 23420
rect 10137 23418 10161 23420
rect 10217 23418 10241 23420
rect 10079 23366 10081 23418
rect 10143 23366 10155 23418
rect 10217 23366 10219 23418
rect 10057 23364 10081 23366
rect 10137 23364 10161 23366
rect 10217 23364 10241 23366
rect 10001 23344 10297 23364
rect 10692 23322 10720 23559
rect 10680 23316 10732 23322
rect 10680 23258 10732 23264
rect 10496 23180 10548 23186
rect 10496 23122 10548 23128
rect 10508 22438 10536 23122
rect 10586 22536 10642 22545
rect 10586 22471 10642 22480
rect 9760 22432 9812 22438
rect 9760 22374 9812 22380
rect 10496 22432 10548 22438
rect 10496 22374 10548 22380
rect 9772 22166 9800 22374
rect 10001 22332 10297 22352
rect 10057 22330 10081 22332
rect 10137 22330 10161 22332
rect 10217 22330 10241 22332
rect 10079 22278 10081 22330
rect 10143 22278 10155 22330
rect 10217 22278 10219 22330
rect 10057 22276 10081 22278
rect 10137 22276 10161 22278
rect 10217 22276 10241 22278
rect 10001 22256 10297 22276
rect 9760 22160 9812 22166
rect 9760 22102 9812 22108
rect 9392 22092 9444 22098
rect 9392 22034 9444 22040
rect 9404 21350 9432 22034
rect 9392 21344 9444 21350
rect 9392 21286 9444 21292
rect 8470 7848 8526 7857
rect 8470 7783 8526 7792
rect 8012 7540 8064 7546
rect 8012 7482 8064 7488
rect 7828 7336 7880 7342
rect 7828 7278 7880 7284
rect 7840 6934 7868 7278
rect 8024 7274 8052 7482
rect 8012 7268 8064 7274
rect 8012 7210 8064 7216
rect 7828 6928 7880 6934
rect 7828 6870 7880 6876
rect 7734 6624 7790 6633
rect 7734 6559 7790 6568
rect 7748 5642 7776 6559
rect 7840 6254 7868 6870
rect 8196 6860 8248 6866
rect 8196 6802 8248 6808
rect 7828 6248 7880 6254
rect 7828 6190 7880 6196
rect 8104 6248 8156 6254
rect 8104 6190 8156 6196
rect 8012 5772 8064 5778
rect 8012 5714 8064 5720
rect 7920 5704 7972 5710
rect 7826 5672 7882 5681
rect 7736 5636 7788 5642
rect 7920 5646 7972 5652
rect 7826 5607 7828 5616
rect 7736 5578 7788 5584
rect 7880 5607 7882 5616
rect 7828 5578 7880 5584
rect 7644 5228 7696 5234
rect 7644 5170 7696 5176
rect 7840 4826 7868 5578
rect 7932 5370 7960 5646
rect 7920 5364 7972 5370
rect 7920 5306 7972 5312
rect 8024 5030 8052 5714
rect 8012 5024 8064 5030
rect 8010 4992 8012 5001
rect 8064 4992 8066 5001
rect 8010 4927 8066 4936
rect 8116 4826 8144 6190
rect 8208 5710 8236 6802
rect 8196 5704 8248 5710
rect 8196 5646 8248 5652
rect 8380 5024 8432 5030
rect 8380 4966 8432 4972
rect 7828 4820 7880 4826
rect 7828 4762 7880 4768
rect 8104 4820 8156 4826
rect 8104 4762 8156 4768
rect 8288 4616 8340 4622
rect 8288 4558 8340 4564
rect 7644 4140 7696 4146
rect 7644 4082 7696 4088
rect 7552 3936 7604 3942
rect 7552 3878 7604 3884
rect 7656 3738 7684 4082
rect 8300 4049 8328 4558
rect 8286 4040 8342 4049
rect 8286 3975 8342 3984
rect 8392 3913 8420 4966
rect 8378 3904 8434 3913
rect 8378 3839 8434 3848
rect 7734 3768 7790 3777
rect 7644 3732 7696 3738
rect 7734 3703 7790 3712
rect 7644 3674 7696 3680
rect 7182 2952 7238 2961
rect 7182 2887 7184 2896
rect 7236 2887 7238 2896
rect 7184 2858 7236 2864
rect 7748 480 7776 3703
rect 8484 3602 8512 7783
rect 9208 7472 9260 7478
rect 9206 7440 9208 7449
rect 9260 7440 9262 7449
rect 9206 7375 9262 7384
rect 9208 7200 9260 7206
rect 9208 7142 9260 7148
rect 9220 6254 9248 7142
rect 9404 6730 9432 21286
rect 10001 21244 10297 21264
rect 10057 21242 10081 21244
rect 10137 21242 10161 21244
rect 10217 21242 10241 21244
rect 10079 21190 10081 21242
rect 10143 21190 10155 21242
rect 10217 21190 10219 21242
rect 10057 21188 10081 21190
rect 10137 21188 10161 21190
rect 10217 21188 10241 21190
rect 10001 21168 10297 21188
rect 9666 21040 9722 21049
rect 9666 20975 9722 20984
rect 9680 12458 9708 20975
rect 10001 20156 10297 20176
rect 10057 20154 10081 20156
rect 10137 20154 10161 20156
rect 10217 20154 10241 20156
rect 10079 20102 10081 20154
rect 10143 20102 10155 20154
rect 10217 20102 10219 20154
rect 10057 20100 10081 20102
rect 10137 20100 10161 20102
rect 10217 20100 10241 20102
rect 10001 20080 10297 20100
rect 10001 19068 10297 19088
rect 10057 19066 10081 19068
rect 10137 19066 10161 19068
rect 10217 19066 10241 19068
rect 10079 19014 10081 19066
rect 10143 19014 10155 19066
rect 10217 19014 10219 19066
rect 10057 19012 10081 19014
rect 10137 19012 10161 19014
rect 10217 19012 10241 19014
rect 10001 18992 10297 19012
rect 10001 17980 10297 18000
rect 10057 17978 10081 17980
rect 10137 17978 10161 17980
rect 10217 17978 10241 17980
rect 10079 17926 10081 17978
rect 10143 17926 10155 17978
rect 10217 17926 10219 17978
rect 10057 17924 10081 17926
rect 10137 17924 10161 17926
rect 10217 17924 10241 17926
rect 10001 17904 10297 17924
rect 9852 17740 9904 17746
rect 9852 17682 9904 17688
rect 9864 16998 9892 17682
rect 9852 16992 9904 16998
rect 9850 16960 9852 16969
rect 9904 16960 9906 16969
rect 9850 16895 9906 16904
rect 10001 16892 10297 16912
rect 10057 16890 10081 16892
rect 10137 16890 10161 16892
rect 10217 16890 10241 16892
rect 10079 16838 10081 16890
rect 10143 16838 10155 16890
rect 10217 16838 10219 16890
rect 10057 16836 10081 16838
rect 10137 16836 10161 16838
rect 10217 16836 10241 16838
rect 10001 16816 10297 16836
rect 10001 15804 10297 15824
rect 10057 15802 10081 15804
rect 10137 15802 10161 15804
rect 10217 15802 10241 15804
rect 10079 15750 10081 15802
rect 10143 15750 10155 15802
rect 10217 15750 10219 15802
rect 10057 15748 10081 15750
rect 10137 15748 10161 15750
rect 10217 15748 10241 15750
rect 10001 15728 10297 15748
rect 10001 14716 10297 14736
rect 10057 14714 10081 14716
rect 10137 14714 10161 14716
rect 10217 14714 10241 14716
rect 10079 14662 10081 14714
rect 10143 14662 10155 14714
rect 10217 14662 10219 14714
rect 10057 14660 10081 14662
rect 10137 14660 10161 14662
rect 10217 14660 10241 14662
rect 10001 14640 10297 14660
rect 10001 13628 10297 13648
rect 10057 13626 10081 13628
rect 10137 13626 10161 13628
rect 10217 13626 10241 13628
rect 10079 13574 10081 13626
rect 10143 13574 10155 13626
rect 10217 13574 10219 13626
rect 10057 13572 10081 13574
rect 10137 13572 10161 13574
rect 10217 13572 10241 13574
rect 10001 13552 10297 13572
rect 10001 12540 10297 12560
rect 10057 12538 10081 12540
rect 10137 12538 10161 12540
rect 10217 12538 10241 12540
rect 10079 12486 10081 12538
rect 10143 12486 10155 12538
rect 10217 12486 10219 12538
rect 10057 12484 10081 12486
rect 10137 12484 10161 12486
rect 10217 12484 10241 12486
rect 10001 12464 10297 12484
rect 9680 12430 9892 12458
rect 9576 8356 9628 8362
rect 9576 8298 9628 8304
rect 9588 6730 9616 8298
rect 9760 7880 9812 7886
rect 9760 7822 9812 7828
rect 9772 7002 9800 7822
rect 9760 6996 9812 7002
rect 9760 6938 9812 6944
rect 9668 6792 9720 6798
rect 9668 6734 9720 6740
rect 9392 6724 9444 6730
rect 9392 6666 9444 6672
rect 9576 6724 9628 6730
rect 9576 6666 9628 6672
rect 9208 6248 9260 6254
rect 9208 6190 9260 6196
rect 9300 6180 9352 6186
rect 9300 6122 9352 6128
rect 9392 6180 9444 6186
rect 9392 6122 9444 6128
rect 9116 5908 9168 5914
rect 9116 5850 9168 5856
rect 9128 5234 9156 5850
rect 9312 5778 9340 6122
rect 9300 5772 9352 5778
rect 9300 5714 9352 5720
rect 9404 5370 9432 6122
rect 9484 6112 9536 6118
rect 9484 6054 9536 6060
rect 9496 5914 9524 6054
rect 9588 5914 9616 6666
rect 9680 6186 9708 6734
rect 9772 6458 9800 6938
rect 9760 6452 9812 6458
rect 9760 6394 9812 6400
rect 9668 6180 9720 6186
rect 9668 6122 9720 6128
rect 9864 5914 9892 12430
rect 10001 11452 10297 11472
rect 10057 11450 10081 11452
rect 10137 11450 10161 11452
rect 10217 11450 10241 11452
rect 10079 11398 10081 11450
rect 10143 11398 10155 11450
rect 10217 11398 10219 11450
rect 10057 11396 10081 11398
rect 10137 11396 10161 11398
rect 10217 11396 10241 11398
rect 10001 11376 10297 11396
rect 10001 10364 10297 10384
rect 10057 10362 10081 10364
rect 10137 10362 10161 10364
rect 10217 10362 10241 10364
rect 10079 10310 10081 10362
rect 10143 10310 10155 10362
rect 10217 10310 10219 10362
rect 10057 10308 10081 10310
rect 10137 10308 10161 10310
rect 10217 10308 10241 10310
rect 10001 10288 10297 10308
rect 10001 9276 10297 9296
rect 10057 9274 10081 9276
rect 10137 9274 10161 9276
rect 10217 9274 10241 9276
rect 10079 9222 10081 9274
rect 10143 9222 10155 9274
rect 10217 9222 10219 9274
rect 10057 9220 10081 9222
rect 10137 9220 10161 9222
rect 10217 9220 10241 9222
rect 10001 9200 10297 9220
rect 10600 9178 10628 22471
rect 12336 22092 12388 22098
rect 12336 22034 12388 22040
rect 12242 21448 12298 21457
rect 12242 21383 12298 21392
rect 11138 19816 11194 19825
rect 11138 19751 11194 19760
rect 11152 18970 11180 19751
rect 11140 18964 11192 18970
rect 11140 18906 11192 18912
rect 10772 18828 10824 18834
rect 10772 18770 10824 18776
rect 10784 18086 10812 18770
rect 10772 18080 10824 18086
rect 10692 18028 10772 18034
rect 10692 18022 10824 18028
rect 10692 18006 10812 18022
rect 10692 17814 10720 18006
rect 10680 17808 10732 17814
rect 10680 17750 10732 17756
rect 12152 17128 12204 17134
rect 12152 17070 12204 17076
rect 10956 9376 11008 9382
rect 10956 9318 11008 9324
rect 10588 9172 10640 9178
rect 10588 9114 10640 9120
rect 10968 9042 10996 9318
rect 10956 9036 11008 9042
rect 10956 8978 11008 8984
rect 10496 8832 10548 8838
rect 10496 8774 10548 8780
rect 10001 8188 10297 8208
rect 10057 8186 10081 8188
rect 10137 8186 10161 8188
rect 10217 8186 10241 8188
rect 10079 8134 10081 8186
rect 10143 8134 10155 8186
rect 10217 8134 10219 8186
rect 10057 8132 10081 8134
rect 10137 8132 10161 8134
rect 10217 8132 10241 8134
rect 10001 8112 10297 8132
rect 10508 7546 10536 8774
rect 10968 8634 10996 8978
rect 11784 8968 11836 8974
rect 12060 8968 12112 8974
rect 11784 8910 11836 8916
rect 11874 8936 11930 8945
rect 11796 8634 11824 8910
rect 12060 8910 12112 8916
rect 11874 8871 11930 8880
rect 10956 8628 11008 8634
rect 10956 8570 11008 8576
rect 11784 8628 11836 8634
rect 11784 8570 11836 8576
rect 10680 8424 10732 8430
rect 10680 8366 10732 8372
rect 10692 7886 10720 8366
rect 10956 8288 11008 8294
rect 10956 8230 11008 8236
rect 10968 7954 10996 8230
rect 11796 8090 11824 8570
rect 11784 8084 11836 8090
rect 11784 8026 11836 8032
rect 10956 7948 11008 7954
rect 10956 7890 11008 7896
rect 10680 7880 10732 7886
rect 10680 7822 10732 7828
rect 10496 7540 10548 7546
rect 10496 7482 10548 7488
rect 10310 7304 10366 7313
rect 10310 7239 10312 7248
rect 10364 7239 10366 7248
rect 10312 7210 10364 7216
rect 10692 7206 10720 7822
rect 10968 7410 10996 7890
rect 10956 7404 11008 7410
rect 10956 7346 11008 7352
rect 10680 7200 10732 7206
rect 10680 7142 10732 7148
rect 10772 7200 10824 7206
rect 10772 7142 10824 7148
rect 10001 7100 10297 7120
rect 10057 7098 10081 7100
rect 10137 7098 10161 7100
rect 10217 7098 10241 7100
rect 10079 7046 10081 7098
rect 10143 7046 10155 7098
rect 10217 7046 10219 7098
rect 10057 7044 10081 7046
rect 10137 7044 10161 7046
rect 10217 7044 10241 7046
rect 10001 7024 10297 7044
rect 10692 6934 10720 7142
rect 10680 6928 10732 6934
rect 10680 6870 10732 6876
rect 10784 6866 10812 7142
rect 10772 6860 10824 6866
rect 10772 6802 10824 6808
rect 11324 6860 11376 6866
rect 11324 6802 11376 6808
rect 11416 6860 11468 6866
rect 11416 6802 11468 6808
rect 11692 6860 11744 6866
rect 11692 6802 11744 6808
rect 10784 6769 10812 6802
rect 10770 6760 10826 6769
rect 10770 6695 10826 6704
rect 11048 6112 11100 6118
rect 11048 6054 11100 6060
rect 10001 6012 10297 6032
rect 10057 6010 10081 6012
rect 10137 6010 10161 6012
rect 10217 6010 10241 6012
rect 10079 5958 10081 6010
rect 10143 5958 10155 6010
rect 10217 5958 10219 6010
rect 10057 5956 10081 5958
rect 10137 5956 10161 5958
rect 10217 5956 10241 5958
rect 10001 5936 10297 5956
rect 11060 5914 11088 6054
rect 9484 5908 9536 5914
rect 9484 5850 9536 5856
rect 9576 5908 9628 5914
rect 9576 5850 9628 5856
rect 9852 5908 9904 5914
rect 9852 5850 9904 5856
rect 11048 5908 11100 5914
rect 11048 5850 11100 5856
rect 11336 5846 11364 6802
rect 9668 5840 9720 5846
rect 9668 5782 9720 5788
rect 11324 5840 11376 5846
rect 11324 5782 11376 5788
rect 9680 5370 9708 5782
rect 9852 5772 9904 5778
rect 9852 5714 9904 5720
rect 11048 5772 11100 5778
rect 11048 5714 11100 5720
rect 9392 5364 9444 5370
rect 9392 5306 9444 5312
rect 9668 5364 9720 5370
rect 9668 5306 9720 5312
rect 9116 5228 9168 5234
rect 9116 5170 9168 5176
rect 9300 5024 9352 5030
rect 9300 4966 9352 4972
rect 9760 5024 9812 5030
rect 9760 4966 9812 4972
rect 8838 4584 8894 4593
rect 9312 4554 9340 4966
rect 8838 4519 8894 4528
rect 9300 4548 9352 4554
rect 8656 3936 8708 3942
rect 8656 3878 8708 3884
rect 8472 3596 8524 3602
rect 8472 3538 8524 3544
rect 8484 3126 8512 3538
rect 8668 3398 8696 3878
rect 8564 3392 8616 3398
rect 8564 3334 8616 3340
rect 8656 3392 8708 3398
rect 8656 3334 8708 3340
rect 8472 3120 8524 3126
rect 8472 3062 8524 3068
rect 8196 2508 8248 2514
rect 8196 2450 8248 2456
rect 7826 2408 7882 2417
rect 7826 2343 7828 2352
rect 7880 2343 7882 2352
rect 7828 2314 7880 2320
rect 8208 1737 8236 2450
rect 8288 2440 8340 2446
rect 8288 2382 8340 2388
rect 8472 2440 8524 2446
rect 8472 2382 8524 2388
rect 8300 2281 8328 2382
rect 8286 2272 8342 2281
rect 8286 2207 8342 2216
rect 8378 2136 8434 2145
rect 8378 2071 8434 2080
rect 8194 1728 8250 1737
rect 8194 1663 8250 1672
rect 8392 480 8420 2071
rect 8484 1601 8512 2382
rect 8576 1873 8604 3334
rect 8668 3194 8696 3334
rect 8852 3194 8880 4519
rect 9300 4490 9352 4496
rect 8932 4072 8984 4078
rect 8932 4014 8984 4020
rect 8944 3942 8972 4014
rect 9312 3942 9340 4490
rect 9668 4480 9720 4486
rect 9668 4422 9720 4428
rect 9680 4146 9708 4422
rect 9772 4185 9800 4966
rect 9864 4826 9892 5714
rect 10312 5704 10364 5710
rect 10312 5646 10364 5652
rect 10324 5370 10352 5646
rect 11060 5574 11088 5714
rect 11428 5710 11456 6802
rect 11704 6746 11732 6802
rect 11520 6718 11732 6746
rect 11520 6118 11548 6718
rect 11508 6112 11560 6118
rect 11508 6054 11560 6060
rect 11416 5704 11468 5710
rect 11520 5681 11548 6054
rect 11888 5794 11916 8871
rect 12072 7410 12100 8910
rect 12060 7404 12112 7410
rect 12060 7346 12112 7352
rect 12072 6934 12100 7346
rect 12060 6928 12112 6934
rect 12060 6870 12112 6876
rect 11796 5766 11916 5794
rect 12060 5840 12112 5846
rect 12060 5782 12112 5788
rect 11416 5646 11468 5652
rect 11506 5672 11562 5681
rect 11506 5607 11562 5616
rect 11048 5568 11100 5574
rect 11048 5510 11100 5516
rect 10312 5364 10364 5370
rect 10312 5306 10364 5312
rect 11060 5234 11088 5510
rect 11048 5228 11100 5234
rect 11048 5170 11100 5176
rect 11324 5160 11376 5166
rect 10954 5128 11010 5137
rect 11324 5102 11376 5108
rect 10954 5063 10956 5072
rect 11008 5063 11010 5072
rect 10956 5034 11008 5040
rect 10001 4924 10297 4944
rect 10057 4922 10081 4924
rect 10137 4922 10161 4924
rect 10217 4922 10241 4924
rect 10079 4870 10081 4922
rect 10143 4870 10155 4922
rect 10217 4870 10219 4922
rect 10057 4868 10081 4870
rect 10137 4868 10161 4870
rect 10217 4868 10241 4870
rect 10001 4848 10297 4868
rect 9852 4820 9904 4826
rect 9852 4762 9904 4768
rect 10680 4684 10732 4690
rect 10680 4626 10732 4632
rect 10128 4616 10180 4622
rect 10128 4558 10180 4564
rect 9758 4176 9814 4185
rect 9668 4140 9720 4146
rect 9758 4111 9814 4120
rect 9668 4082 9720 4088
rect 9392 4004 9444 4010
rect 9392 3946 9444 3952
rect 8932 3936 8984 3942
rect 8932 3878 8984 3884
rect 9300 3936 9352 3942
rect 9300 3878 9352 3884
rect 8944 3777 8972 3878
rect 8930 3768 8986 3777
rect 8930 3703 8986 3712
rect 9300 3664 9352 3670
rect 9022 3632 9078 3641
rect 9300 3606 9352 3612
rect 9022 3567 9078 3576
rect 8656 3188 8708 3194
rect 8656 3130 8708 3136
rect 8840 3188 8892 3194
rect 8840 3130 8892 3136
rect 8852 2990 8880 3130
rect 8840 2984 8892 2990
rect 8840 2926 8892 2932
rect 8656 2848 8708 2854
rect 8656 2790 8708 2796
rect 8668 2009 8696 2790
rect 8654 2000 8710 2009
rect 8654 1935 8710 1944
rect 8562 1864 8618 1873
rect 8562 1799 8618 1808
rect 8470 1592 8526 1601
rect 8470 1527 8526 1536
rect 9036 480 9064 3567
rect 9312 2650 9340 3606
rect 9404 3534 9432 3946
rect 9576 3936 9628 3942
rect 9576 3878 9628 3884
rect 9392 3528 9444 3534
rect 9392 3470 9444 3476
rect 9588 3398 9616 3878
rect 9680 3670 9708 4082
rect 10140 4010 10168 4558
rect 10692 4214 10720 4626
rect 10680 4208 10732 4214
rect 10680 4150 10732 4156
rect 10128 4004 10180 4010
rect 10128 3946 10180 3952
rect 10402 3904 10458 3913
rect 10001 3836 10297 3856
rect 10402 3839 10458 3848
rect 10057 3834 10081 3836
rect 10137 3834 10161 3836
rect 10217 3834 10241 3836
rect 10079 3782 10081 3834
rect 10143 3782 10155 3834
rect 10217 3782 10219 3834
rect 10057 3780 10081 3782
rect 10137 3780 10161 3782
rect 10217 3780 10241 3782
rect 10001 3760 10297 3780
rect 9668 3664 9720 3670
rect 9668 3606 9720 3612
rect 9576 3392 9628 3398
rect 9576 3334 9628 3340
rect 9680 3194 9708 3606
rect 9850 3360 9906 3369
rect 9850 3295 9906 3304
rect 9668 3188 9720 3194
rect 9668 3130 9720 3136
rect 9300 2644 9352 2650
rect 9300 2586 9352 2592
rect 9864 626 9892 3295
rect 10416 2990 10444 3839
rect 10692 3738 10720 4150
rect 10680 3732 10732 3738
rect 10680 3674 10732 3680
rect 10496 3392 10548 3398
rect 10496 3334 10548 3340
rect 10404 2984 10456 2990
rect 10404 2926 10456 2932
rect 10404 2848 10456 2854
rect 10508 2825 10536 3334
rect 10404 2790 10456 2796
rect 10494 2816 10550 2825
rect 10001 2748 10297 2768
rect 10057 2746 10081 2748
rect 10137 2746 10161 2748
rect 10217 2746 10241 2748
rect 10079 2694 10081 2746
rect 10143 2694 10155 2746
rect 10217 2694 10219 2746
rect 10057 2692 10081 2694
rect 10137 2692 10161 2694
rect 10217 2692 10241 2694
rect 10001 2672 10297 2692
rect 10416 2514 10444 2790
rect 10494 2751 10550 2760
rect 10678 2680 10734 2689
rect 10678 2615 10680 2624
rect 10732 2615 10734 2624
rect 10680 2586 10732 2592
rect 10968 2582 10996 5034
rect 11046 4720 11102 4729
rect 11046 4655 11102 4664
rect 10956 2576 11008 2582
rect 10956 2518 11008 2524
rect 10404 2508 10456 2514
rect 10404 2450 10456 2456
rect 10496 2508 10548 2514
rect 10496 2450 10548 2456
rect 10508 2310 10536 2450
rect 10404 2304 10456 2310
rect 10310 2272 10366 2281
rect 10404 2246 10456 2252
rect 10496 2304 10548 2310
rect 10496 2246 10548 2252
rect 10310 2207 10366 2216
rect 10324 1306 10352 2207
rect 10416 1465 10444 2246
rect 10508 2145 10536 2246
rect 10494 2136 10550 2145
rect 10494 2071 10550 2080
rect 10402 1456 10458 1465
rect 10402 1391 10458 1400
rect 10324 1278 10444 1306
rect 9772 598 9892 626
rect 9772 480 9800 598
rect 10416 480 10444 1278
rect 11060 480 11088 4655
rect 11336 4010 11364 5102
rect 11520 4826 11548 5607
rect 11508 4820 11560 4826
rect 11508 4762 11560 4768
rect 11598 4176 11654 4185
rect 11598 4111 11600 4120
rect 11652 4111 11654 4120
rect 11600 4082 11652 4088
rect 11324 4004 11376 4010
rect 11324 3946 11376 3952
rect 11140 3936 11192 3942
rect 11140 3878 11192 3884
rect 11152 3777 11180 3878
rect 11138 3768 11194 3777
rect 11336 3738 11364 3946
rect 11138 3703 11194 3712
rect 11324 3732 11376 3738
rect 11324 3674 11376 3680
rect 11796 626 11824 5766
rect 12072 4690 12100 5782
rect 12060 4684 12112 4690
rect 12060 4626 12112 4632
rect 11876 4072 11928 4078
rect 11874 4040 11876 4049
rect 11928 4040 11930 4049
rect 11874 3975 11930 3984
rect 12164 3942 12192 17070
rect 12256 6458 12284 21383
rect 12348 21350 12376 22034
rect 12428 22024 12480 22030
rect 12426 21992 12428 22001
rect 12480 21992 12482 22001
rect 12426 21927 12482 21936
rect 12336 21344 12388 21350
rect 12336 21286 12388 21292
rect 12348 21049 12376 21286
rect 12334 21040 12390 21049
rect 12334 20975 12390 20984
rect 12886 17096 12942 17105
rect 12886 17031 12888 17040
rect 12940 17031 12942 17040
rect 12888 17002 12940 17008
rect 13544 16561 13572 27390
rect 14668 25052 14964 25072
rect 14724 25050 14748 25052
rect 14804 25050 14828 25052
rect 14884 25050 14908 25052
rect 14746 24998 14748 25050
rect 14810 24998 14822 25050
rect 14884 24998 14886 25050
rect 14724 24996 14748 24998
rect 14804 24996 14828 24998
rect 14884 24996 14908 24998
rect 14668 24976 14964 24996
rect 14668 23964 14964 23984
rect 14724 23962 14748 23964
rect 14804 23962 14828 23964
rect 14884 23962 14908 23964
rect 14746 23910 14748 23962
rect 14810 23910 14822 23962
rect 14884 23910 14886 23962
rect 14724 23908 14748 23910
rect 14804 23908 14828 23910
rect 14884 23908 14908 23910
rect 14668 23888 14964 23908
rect 19248 23225 19276 27520
rect 23558 27160 23614 27169
rect 23558 27095 23614 27104
rect 23466 26616 23522 26625
rect 23466 26551 23522 26560
rect 19334 25596 19630 25616
rect 19390 25594 19414 25596
rect 19470 25594 19494 25596
rect 19550 25594 19574 25596
rect 19412 25542 19414 25594
rect 19476 25542 19488 25594
rect 19550 25542 19552 25594
rect 19390 25540 19414 25542
rect 19470 25540 19494 25542
rect 19550 25540 19574 25542
rect 19334 25520 19630 25540
rect 19334 24508 19630 24528
rect 19390 24506 19414 24508
rect 19470 24506 19494 24508
rect 19550 24506 19574 24508
rect 19412 24454 19414 24506
rect 19476 24454 19488 24506
rect 19550 24454 19552 24506
rect 19390 24452 19414 24454
rect 19470 24452 19494 24454
rect 19550 24452 19574 24454
rect 19334 24432 19630 24452
rect 19334 23420 19630 23440
rect 19390 23418 19414 23420
rect 19470 23418 19494 23420
rect 19550 23418 19574 23420
rect 19412 23366 19414 23418
rect 19476 23366 19488 23418
rect 19550 23366 19552 23418
rect 19390 23364 19414 23366
rect 19470 23364 19494 23366
rect 19550 23364 19574 23366
rect 19334 23344 19630 23364
rect 19234 23216 19290 23225
rect 19234 23151 19290 23160
rect 14668 22876 14964 22896
rect 14724 22874 14748 22876
rect 14804 22874 14828 22876
rect 14884 22874 14908 22876
rect 14746 22822 14748 22874
rect 14810 22822 14822 22874
rect 14884 22822 14886 22874
rect 14724 22820 14748 22822
rect 14804 22820 14828 22822
rect 14884 22820 14908 22822
rect 14668 22800 14964 22820
rect 23190 22536 23246 22545
rect 23190 22471 23192 22480
rect 23244 22471 23246 22480
rect 23192 22442 23244 22448
rect 19334 22332 19630 22352
rect 19390 22330 19414 22332
rect 19470 22330 19494 22332
rect 19550 22330 19574 22332
rect 19412 22278 19414 22330
rect 19476 22278 19488 22330
rect 19550 22278 19552 22330
rect 19390 22276 19414 22278
rect 19470 22276 19494 22278
rect 19550 22276 19574 22278
rect 19334 22256 19630 22276
rect 23480 21842 23508 26551
rect 23296 21814 23508 21842
rect 14668 21788 14964 21808
rect 14724 21786 14748 21788
rect 14804 21786 14828 21788
rect 14884 21786 14908 21788
rect 14746 21734 14748 21786
rect 14810 21734 14822 21786
rect 14884 21734 14886 21786
rect 14724 21732 14748 21734
rect 14804 21732 14828 21734
rect 14884 21732 14908 21734
rect 14668 21712 14964 21732
rect 14728 21480 14780 21486
rect 14726 21448 14728 21457
rect 14780 21448 14782 21457
rect 14726 21383 14782 21392
rect 15002 21448 15058 21457
rect 15002 21383 15004 21392
rect 15056 21383 15058 21392
rect 15004 21354 15056 21360
rect 19334 21244 19630 21264
rect 19390 21242 19414 21244
rect 19470 21242 19494 21244
rect 19550 21242 19574 21244
rect 19412 21190 19414 21242
rect 19476 21190 19488 21242
rect 19550 21190 19552 21242
rect 19390 21188 19414 21190
rect 19470 21188 19494 21190
rect 19550 21188 19574 21190
rect 19334 21168 19630 21188
rect 23192 21004 23244 21010
rect 23192 20946 23244 20952
rect 14668 20700 14964 20720
rect 14724 20698 14748 20700
rect 14804 20698 14828 20700
rect 14884 20698 14908 20700
rect 14746 20646 14748 20698
rect 14810 20646 14822 20698
rect 14884 20646 14886 20698
rect 14724 20644 14748 20646
rect 14804 20644 14828 20646
rect 14884 20644 14908 20646
rect 14668 20624 14964 20644
rect 23204 20398 23232 20946
rect 23192 20392 23244 20398
rect 15646 20360 15702 20369
rect 15646 20295 15702 20304
rect 23190 20360 23192 20369
rect 23244 20360 23246 20369
rect 23190 20295 23246 20304
rect 14668 19612 14964 19632
rect 14724 19610 14748 19612
rect 14804 19610 14828 19612
rect 14884 19610 14908 19612
rect 14746 19558 14748 19610
rect 14810 19558 14822 19610
rect 14884 19558 14886 19610
rect 14724 19556 14748 19558
rect 14804 19556 14828 19558
rect 14884 19556 14908 19558
rect 14668 19536 14964 19556
rect 15372 18828 15424 18834
rect 15372 18770 15424 18776
rect 14668 18524 14964 18544
rect 14724 18522 14748 18524
rect 14804 18522 14828 18524
rect 14884 18522 14908 18524
rect 14746 18470 14748 18522
rect 14810 18470 14822 18522
rect 14884 18470 14886 18522
rect 14724 18468 14748 18470
rect 14804 18468 14828 18470
rect 14884 18468 14908 18470
rect 14668 18448 14964 18468
rect 15384 18086 15412 18770
rect 15372 18080 15424 18086
rect 15372 18022 15424 18028
rect 14668 17436 14964 17456
rect 14724 17434 14748 17436
rect 14804 17434 14828 17436
rect 14884 17434 14908 17436
rect 14746 17382 14748 17434
rect 14810 17382 14822 17434
rect 14884 17382 14886 17434
rect 14724 17380 14748 17382
rect 14804 17380 14828 17382
rect 14884 17380 14908 17382
rect 14668 17360 14964 17380
rect 15004 16652 15056 16658
rect 15004 16594 15056 16600
rect 13530 16552 13586 16561
rect 13530 16487 13586 16496
rect 14668 16348 14964 16368
rect 14724 16346 14748 16348
rect 14804 16346 14828 16348
rect 14884 16346 14908 16348
rect 14746 16294 14748 16346
rect 14810 16294 14822 16346
rect 14884 16294 14886 16346
rect 14724 16292 14748 16294
rect 14804 16292 14828 16294
rect 14884 16292 14908 16294
rect 14668 16272 14964 16292
rect 15016 15910 15044 16594
rect 15004 15904 15056 15910
rect 12426 15872 12482 15881
rect 12426 15807 12482 15816
rect 15002 15872 15004 15881
rect 15056 15872 15058 15881
rect 15002 15807 15058 15816
rect 12336 9104 12388 9110
rect 12336 9046 12388 9052
rect 12348 8634 12376 9046
rect 12336 8628 12388 8634
rect 12336 8570 12388 8576
rect 12244 6452 12296 6458
rect 12244 6394 12296 6400
rect 12152 3936 12204 3942
rect 12152 3878 12204 3884
rect 12334 3768 12390 3777
rect 12334 3703 12390 3712
rect 11968 3596 12020 3602
rect 11968 3538 12020 3544
rect 12152 3596 12204 3602
rect 12152 3538 12204 3544
rect 11874 2952 11930 2961
rect 11874 2887 11876 2896
rect 11928 2887 11930 2896
rect 11876 2858 11928 2864
rect 11980 2514 12008 3538
rect 12164 2990 12192 3538
rect 12152 2984 12204 2990
rect 12152 2926 12204 2932
rect 12060 2644 12112 2650
rect 12164 2632 12192 2926
rect 12112 2604 12192 2632
rect 12060 2586 12112 2592
rect 11968 2508 12020 2514
rect 11968 2450 12020 2456
rect 11704 598 11824 626
rect 11704 480 11732 598
rect 12348 480 12376 3703
rect 12440 3194 12468 15807
rect 14668 15260 14964 15280
rect 14724 15258 14748 15260
rect 14804 15258 14828 15260
rect 14884 15258 14908 15260
rect 14746 15206 14748 15258
rect 14810 15206 14822 15258
rect 14884 15206 14886 15258
rect 14724 15204 14748 15206
rect 14804 15204 14828 15206
rect 14884 15204 14908 15206
rect 14668 15184 14964 15204
rect 13162 14920 13218 14929
rect 13162 14855 13218 14864
rect 12612 9376 12664 9382
rect 12612 9318 12664 9324
rect 13070 9344 13126 9353
rect 12624 9081 12652 9318
rect 13070 9279 13126 9288
rect 12610 9072 12666 9081
rect 12610 9007 12666 9016
rect 12520 8288 12572 8294
rect 12520 8230 12572 8236
rect 12532 7954 12560 8230
rect 12520 7948 12572 7954
rect 12520 7890 12572 7896
rect 12532 7546 12560 7890
rect 12980 7812 13032 7818
rect 12980 7754 13032 7760
rect 12520 7540 12572 7546
rect 12520 7482 12572 7488
rect 12992 7342 13020 7754
rect 12980 7336 13032 7342
rect 12980 7278 13032 7284
rect 12992 7002 13020 7278
rect 12980 6996 13032 7002
rect 12980 6938 13032 6944
rect 13084 6882 13112 9279
rect 13176 8090 13204 14855
rect 15186 14512 15242 14521
rect 15186 14447 15242 14456
rect 14668 14172 14964 14192
rect 14724 14170 14748 14172
rect 14804 14170 14828 14172
rect 14884 14170 14908 14172
rect 14746 14118 14748 14170
rect 14810 14118 14822 14170
rect 14884 14118 14886 14170
rect 14724 14116 14748 14118
rect 14804 14116 14828 14118
rect 14884 14116 14908 14118
rect 14668 14096 14964 14116
rect 15002 13288 15058 13297
rect 15002 13223 15058 13232
rect 14668 13084 14964 13104
rect 14724 13082 14748 13084
rect 14804 13082 14828 13084
rect 14884 13082 14908 13084
rect 14746 13030 14748 13082
rect 14810 13030 14822 13082
rect 14884 13030 14886 13082
rect 14724 13028 14748 13030
rect 14804 13028 14828 13030
rect 14884 13028 14908 13030
rect 14668 13008 14964 13028
rect 14668 11996 14964 12016
rect 14724 11994 14748 11996
rect 14804 11994 14828 11996
rect 14884 11994 14908 11996
rect 14746 11942 14748 11994
rect 14810 11942 14822 11994
rect 14884 11942 14886 11994
rect 14724 11940 14748 11942
rect 14804 11940 14828 11942
rect 14884 11940 14908 11942
rect 14668 11920 14964 11940
rect 13622 11656 13678 11665
rect 13622 11591 13678 11600
rect 13636 11218 13664 11591
rect 15016 11393 15044 13223
rect 14450 11384 14506 11393
rect 14450 11319 14506 11328
rect 15002 11384 15058 11393
rect 15002 11319 15058 11328
rect 13624 11212 13676 11218
rect 13624 11154 13676 11160
rect 13636 11098 13664 11154
rect 13452 11070 13664 11098
rect 13716 11144 13768 11150
rect 13716 11086 13768 11092
rect 13452 10810 13480 11070
rect 13440 10804 13492 10810
rect 13440 10746 13492 10752
rect 13624 9920 13676 9926
rect 13624 9862 13676 9868
rect 13636 9586 13664 9862
rect 13624 9580 13676 9586
rect 13624 9522 13676 9528
rect 13532 9444 13584 9450
rect 13532 9386 13584 9392
rect 13544 9178 13572 9386
rect 13532 9172 13584 9178
rect 13532 9114 13584 9120
rect 13636 9110 13664 9522
rect 13624 9104 13676 9110
rect 13624 9046 13676 9052
rect 13346 8392 13402 8401
rect 13346 8327 13348 8336
rect 13400 8327 13402 8336
rect 13348 8298 13400 8304
rect 13164 8084 13216 8090
rect 13164 8026 13216 8032
rect 13624 7880 13676 7886
rect 13624 7822 13676 7828
rect 12992 6854 13112 6882
rect 12888 6316 12940 6322
rect 12888 6258 12940 6264
rect 12612 6112 12664 6118
rect 12612 6054 12664 6060
rect 12704 6112 12756 6118
rect 12704 6054 12756 6060
rect 12624 5914 12652 6054
rect 12612 5908 12664 5914
rect 12612 5850 12664 5856
rect 12612 5636 12664 5642
rect 12612 5578 12664 5584
rect 12624 5098 12652 5578
rect 12612 5092 12664 5098
rect 12612 5034 12664 5040
rect 12624 4570 12652 5034
rect 12716 4826 12744 6054
rect 12900 5166 12928 6258
rect 12888 5160 12940 5166
rect 12888 5102 12940 5108
rect 12704 4820 12756 4826
rect 12704 4762 12756 4768
rect 12624 4542 12744 4570
rect 12716 4486 12744 4542
rect 12796 4548 12848 4554
rect 12796 4490 12848 4496
rect 12612 4480 12664 4486
rect 12612 4422 12664 4428
rect 12704 4480 12756 4486
rect 12704 4422 12756 4428
rect 12624 3942 12652 4422
rect 12716 4078 12744 4422
rect 12808 4146 12836 4490
rect 12796 4140 12848 4146
rect 12796 4082 12848 4088
rect 12704 4072 12756 4078
rect 12704 4014 12756 4020
rect 12612 3936 12664 3942
rect 12808 3913 12836 4082
rect 12612 3878 12664 3884
rect 12794 3904 12850 3913
rect 12428 3188 12480 3194
rect 12428 3130 12480 3136
rect 12624 2689 12652 3878
rect 12794 3839 12850 3848
rect 12808 3738 12836 3839
rect 12796 3732 12848 3738
rect 12796 3674 12848 3680
rect 12888 3392 12940 3398
rect 12888 3334 12940 3340
rect 12900 2961 12928 3334
rect 12886 2952 12942 2961
rect 12886 2887 12888 2896
rect 12940 2887 12942 2896
rect 12888 2858 12940 2864
rect 12610 2680 12666 2689
rect 12610 2615 12666 2624
rect 12992 480 13020 6854
rect 13636 6662 13664 7822
rect 13624 6656 13676 6662
rect 13622 6624 13624 6633
rect 13676 6624 13678 6633
rect 13622 6559 13678 6568
rect 13624 6112 13676 6118
rect 13624 6054 13676 6060
rect 13532 4684 13584 4690
rect 13532 4626 13584 4632
rect 13544 4060 13572 4626
rect 13636 4554 13664 6054
rect 13624 4548 13676 4554
rect 13624 4490 13676 4496
rect 13360 4032 13572 4060
rect 13360 3942 13388 4032
rect 13348 3936 13400 3942
rect 13348 3878 13400 3884
rect 13360 3505 13388 3878
rect 13346 3496 13402 3505
rect 13346 3431 13402 3440
rect 13072 3052 13124 3058
rect 13072 2994 13124 3000
rect 13084 2689 13112 2994
rect 13532 2984 13584 2990
rect 13532 2926 13584 2932
rect 13070 2680 13126 2689
rect 13544 2650 13572 2926
rect 13728 2854 13756 11086
rect 13900 10532 13952 10538
rect 13900 10474 13952 10480
rect 13912 10266 13940 10474
rect 14360 10464 14412 10470
rect 14360 10406 14412 10412
rect 13900 10260 13952 10266
rect 13900 10202 13952 10208
rect 14372 9926 14400 10406
rect 14360 9920 14412 9926
rect 14360 9862 14412 9868
rect 14084 9172 14136 9178
rect 14084 9114 14136 9120
rect 14096 8498 14124 9114
rect 14372 8634 14400 9862
rect 14360 8628 14412 8634
rect 14360 8570 14412 8576
rect 14084 8492 14136 8498
rect 14084 8434 14136 8440
rect 14268 8424 14320 8430
rect 14268 8366 14320 8372
rect 14280 7002 14308 8366
rect 14358 8120 14414 8129
rect 14358 8055 14414 8064
rect 14372 7857 14400 8055
rect 14358 7848 14414 7857
rect 14358 7783 14414 7792
rect 14360 7472 14412 7478
rect 14360 7414 14412 7420
rect 14268 6996 14320 7002
rect 14268 6938 14320 6944
rect 13900 6792 13952 6798
rect 13900 6734 13952 6740
rect 13808 6656 13860 6662
rect 13808 6598 13860 6604
rect 13820 6254 13848 6598
rect 13808 6248 13860 6254
rect 13808 6190 13860 6196
rect 13820 5642 13848 6190
rect 13808 5636 13860 5642
rect 13808 5578 13860 5584
rect 13912 5001 13940 6734
rect 14176 5636 14228 5642
rect 14176 5578 14228 5584
rect 14188 5370 14216 5578
rect 14176 5364 14228 5370
rect 14176 5306 14228 5312
rect 14188 5234 14216 5306
rect 14176 5228 14228 5234
rect 14176 5170 14228 5176
rect 13898 4992 13954 5001
rect 13898 4927 13954 4936
rect 14188 4826 14216 5170
rect 14372 5166 14400 7414
rect 14360 5160 14412 5166
rect 14360 5102 14412 5108
rect 14464 4978 14492 11319
rect 15004 11212 15056 11218
rect 15004 11154 15056 11160
rect 14668 10908 14964 10928
rect 14724 10906 14748 10908
rect 14804 10906 14828 10908
rect 14884 10906 14908 10908
rect 14746 10854 14748 10906
rect 14810 10854 14822 10906
rect 14884 10854 14886 10906
rect 14724 10852 14748 10854
rect 14804 10852 14828 10854
rect 14884 10852 14908 10854
rect 14668 10832 14964 10852
rect 15016 10742 15044 11154
rect 15004 10736 15056 10742
rect 15004 10678 15056 10684
rect 14728 10668 14780 10674
rect 14728 10610 14780 10616
rect 14740 10198 14768 10610
rect 14728 10192 14780 10198
rect 14728 10134 14780 10140
rect 15004 10192 15056 10198
rect 15004 10134 15056 10140
rect 14668 9820 14964 9840
rect 14724 9818 14748 9820
rect 14804 9818 14828 9820
rect 14884 9818 14908 9820
rect 14746 9766 14748 9818
rect 14810 9766 14822 9818
rect 14884 9766 14886 9818
rect 14724 9764 14748 9766
rect 14804 9764 14828 9766
rect 14884 9764 14908 9766
rect 14668 9744 14964 9764
rect 15016 9722 15044 10134
rect 15096 10124 15148 10130
rect 15096 10066 15148 10072
rect 15004 9716 15056 9722
rect 15004 9658 15056 9664
rect 14668 8732 14964 8752
rect 14724 8730 14748 8732
rect 14804 8730 14828 8732
rect 14884 8730 14908 8732
rect 14746 8678 14748 8730
rect 14810 8678 14822 8730
rect 14884 8678 14886 8730
rect 14724 8676 14748 8678
rect 14804 8676 14828 8678
rect 14884 8676 14908 8678
rect 14668 8656 14964 8676
rect 15108 8498 15136 10066
rect 15096 8492 15148 8498
rect 15016 8452 15096 8480
rect 14820 8356 14872 8362
rect 14820 8298 14872 8304
rect 14832 8090 14860 8298
rect 14820 8084 14872 8090
rect 14820 8026 14872 8032
rect 14544 7948 14596 7954
rect 14544 7890 14596 7896
rect 14556 7206 14584 7890
rect 15016 7886 15044 8452
rect 15096 8434 15148 8440
rect 15004 7880 15056 7886
rect 15004 7822 15056 7828
rect 14668 7644 14964 7664
rect 14724 7642 14748 7644
rect 14804 7642 14828 7644
rect 14884 7642 14908 7644
rect 14746 7590 14748 7642
rect 14810 7590 14822 7642
rect 14884 7590 14886 7642
rect 14724 7588 14748 7590
rect 14804 7588 14828 7590
rect 14884 7588 14908 7590
rect 14668 7568 14964 7588
rect 15200 7546 15228 14447
rect 15278 11248 15334 11257
rect 15278 11183 15280 11192
rect 15332 11183 15334 11192
rect 15280 11154 15332 11160
rect 15384 9178 15412 18022
rect 15372 9172 15424 9178
rect 15372 9114 15424 9120
rect 15370 9072 15426 9081
rect 15370 9007 15372 9016
rect 15424 9007 15426 9016
rect 15464 9036 15516 9042
rect 15372 8978 15424 8984
rect 15464 8978 15516 8984
rect 15384 8634 15412 8978
rect 15372 8628 15424 8634
rect 15372 8570 15424 8576
rect 15188 7540 15240 7546
rect 15188 7482 15240 7488
rect 15200 7342 15228 7482
rect 15188 7336 15240 7342
rect 15188 7278 15240 7284
rect 14544 7200 14596 7206
rect 14544 7142 14596 7148
rect 14556 6798 14584 7142
rect 15370 6896 15426 6905
rect 15370 6831 15426 6840
rect 14544 6792 14596 6798
rect 14544 6734 14596 6740
rect 14556 5914 14584 6734
rect 15384 6730 15412 6831
rect 15476 6730 15504 8978
rect 15556 8968 15608 8974
rect 15556 8910 15608 8916
rect 15568 8362 15596 8910
rect 15556 8356 15608 8362
rect 15556 8298 15608 8304
rect 15556 6996 15608 7002
rect 15556 6938 15608 6944
rect 15372 6724 15424 6730
rect 15372 6666 15424 6672
rect 15464 6724 15516 6730
rect 15464 6666 15516 6672
rect 14668 6556 14964 6576
rect 14724 6554 14748 6556
rect 14804 6554 14828 6556
rect 14884 6554 14908 6556
rect 14746 6502 14748 6554
rect 14810 6502 14822 6554
rect 14884 6502 14886 6554
rect 14724 6500 14748 6502
rect 14804 6500 14828 6502
rect 14884 6500 14908 6502
rect 14668 6480 14964 6500
rect 15568 6497 15596 6938
rect 15554 6488 15610 6497
rect 15554 6423 15610 6432
rect 15568 5914 15596 6423
rect 14544 5908 14596 5914
rect 14544 5850 14596 5856
rect 15556 5908 15608 5914
rect 15556 5850 15608 5856
rect 15002 5808 15058 5817
rect 15002 5743 15004 5752
rect 15056 5743 15058 5752
rect 15004 5714 15056 5720
rect 14668 5468 14964 5488
rect 14724 5466 14748 5468
rect 14804 5466 14828 5468
rect 14884 5466 14908 5468
rect 14746 5414 14748 5466
rect 14810 5414 14822 5466
rect 14884 5414 14886 5466
rect 14724 5412 14748 5414
rect 14804 5412 14828 5414
rect 14884 5412 14908 5414
rect 14668 5392 14964 5412
rect 15280 5092 15332 5098
rect 15280 5034 15332 5040
rect 14280 4950 14492 4978
rect 14544 5024 14596 5030
rect 14544 4966 14596 4972
rect 14176 4820 14228 4826
rect 14176 4762 14228 4768
rect 13808 4616 13860 4622
rect 13808 4558 13860 4564
rect 14084 4616 14136 4622
rect 14084 4558 14136 4564
rect 13820 3942 13848 4558
rect 14096 4282 14124 4558
rect 14084 4276 14136 4282
rect 14084 4218 14136 4224
rect 13900 4072 13952 4078
rect 13900 4014 13952 4020
rect 13992 4072 14044 4078
rect 13992 4014 14044 4020
rect 13808 3936 13860 3942
rect 13808 3878 13860 3884
rect 13912 3058 13940 4014
rect 14004 3738 14032 4014
rect 13992 3732 14044 3738
rect 13992 3674 14044 3680
rect 13900 3052 13952 3058
rect 13900 2994 13952 3000
rect 13716 2848 13768 2854
rect 13716 2790 13768 2796
rect 13070 2615 13126 2624
rect 13532 2644 13584 2650
rect 13084 2582 13112 2615
rect 13532 2586 13584 2592
rect 13072 2576 13124 2582
rect 13072 2518 13124 2524
rect 13912 2514 13940 2994
rect 13900 2508 13952 2514
rect 13900 2450 13952 2456
rect 13622 1456 13678 1465
rect 13622 1391 13678 1400
rect 13636 480 13664 1391
rect 14280 480 14308 4950
rect 14358 4856 14414 4865
rect 14358 4791 14414 4800
rect 14372 4457 14400 4791
rect 14556 4758 14584 4966
rect 15292 4826 15320 5034
rect 15660 4826 15688 20295
rect 21442 20224 21498 20233
rect 19334 20156 19630 20176
rect 21442 20159 21498 20168
rect 19390 20154 19414 20156
rect 19470 20154 19494 20156
rect 19550 20154 19574 20156
rect 19412 20102 19414 20154
rect 19476 20102 19488 20154
rect 19550 20102 19552 20154
rect 19390 20100 19414 20102
rect 19470 20100 19494 20102
rect 19550 20100 19574 20102
rect 19334 20080 19630 20100
rect 21456 19990 21484 20159
rect 21444 19984 21496 19990
rect 21444 19926 21496 19932
rect 21168 19916 21220 19922
rect 21168 19858 21220 19864
rect 22456 19916 22508 19922
rect 22456 19858 22508 19864
rect 21180 19174 21208 19858
rect 22468 19174 22496 19858
rect 20616 19168 20668 19174
rect 20616 19110 20668 19116
rect 21168 19168 21220 19174
rect 21168 19110 21220 19116
rect 22456 19168 22508 19174
rect 22456 19110 22508 19116
rect 19334 19068 19630 19088
rect 19390 19066 19414 19068
rect 19470 19066 19494 19068
rect 19550 19066 19574 19068
rect 19412 19014 19414 19066
rect 19476 19014 19488 19066
rect 19550 19014 19552 19066
rect 19390 19012 19414 19014
rect 19470 19012 19494 19014
rect 19550 19012 19574 19014
rect 19334 18992 19630 19012
rect 15738 18864 15794 18873
rect 15738 18799 15740 18808
rect 15792 18799 15794 18808
rect 15740 18770 15792 18776
rect 19334 17980 19630 18000
rect 19390 17978 19414 17980
rect 19470 17978 19494 17980
rect 19550 17978 19574 17980
rect 19412 17926 19414 17978
rect 19476 17926 19488 17978
rect 19550 17926 19552 17978
rect 19390 17924 19414 17926
rect 19470 17924 19494 17926
rect 19550 17924 19574 17926
rect 19334 17904 19630 17924
rect 15832 17740 15884 17746
rect 15832 17682 15884 17688
rect 15844 16998 15872 17682
rect 16014 17640 16070 17649
rect 16014 17575 16016 17584
rect 16068 17575 16070 17584
rect 16016 17546 16068 17552
rect 16106 17368 16162 17377
rect 16106 17303 16162 17312
rect 15832 16992 15884 16998
rect 15832 16934 15884 16940
rect 15844 16726 15872 16934
rect 15832 16720 15884 16726
rect 15832 16662 15884 16668
rect 15922 11792 15978 11801
rect 15922 11727 15924 11736
rect 15976 11727 15978 11736
rect 15924 11698 15976 11704
rect 16016 11620 16068 11626
rect 16016 11562 16068 11568
rect 15832 11212 15884 11218
rect 15832 11154 15884 11160
rect 15738 10160 15794 10169
rect 15844 10130 15872 11154
rect 15738 10095 15794 10104
rect 15832 10124 15884 10130
rect 15280 4820 15332 4826
rect 15280 4762 15332 4768
rect 15648 4820 15700 4826
rect 15648 4762 15700 4768
rect 14544 4752 14596 4758
rect 14544 4694 14596 4700
rect 15004 4752 15056 4758
rect 15004 4694 15056 4700
rect 14358 4448 14414 4457
rect 14358 4383 14414 4392
rect 14556 3738 14584 4694
rect 14668 4380 14964 4400
rect 14724 4378 14748 4380
rect 14804 4378 14828 4380
rect 14884 4378 14908 4380
rect 14746 4326 14748 4378
rect 14810 4326 14822 4378
rect 14884 4326 14886 4378
rect 14724 4324 14748 4326
rect 14804 4324 14828 4326
rect 14884 4324 14908 4326
rect 14668 4304 14964 4324
rect 15016 4264 15044 4694
rect 15292 4457 15320 4762
rect 15278 4448 15334 4457
rect 15278 4383 15334 4392
rect 14832 4236 15044 4264
rect 14832 3738 14860 4236
rect 15464 3936 15516 3942
rect 15464 3878 15516 3884
rect 14544 3732 14596 3738
rect 14544 3674 14596 3680
rect 14820 3732 14872 3738
rect 14820 3674 14872 3680
rect 15370 3632 15426 3641
rect 15476 3602 15504 3878
rect 15370 3567 15372 3576
rect 15424 3567 15426 3576
rect 15464 3596 15516 3602
rect 15372 3538 15424 3544
rect 15464 3538 15516 3544
rect 14542 3496 14598 3505
rect 14542 3431 14598 3440
rect 14556 2922 14584 3431
rect 15004 3392 15056 3398
rect 15004 3334 15056 3340
rect 14668 3292 14964 3312
rect 14724 3290 14748 3292
rect 14804 3290 14828 3292
rect 14884 3290 14908 3292
rect 14746 3238 14748 3290
rect 14810 3238 14822 3290
rect 14884 3238 14886 3290
rect 14724 3236 14748 3238
rect 14804 3236 14828 3238
rect 14884 3236 14908 3238
rect 14668 3216 14964 3236
rect 15016 2961 15044 3334
rect 15096 3120 15148 3126
rect 15096 3062 15148 3068
rect 15002 2952 15058 2961
rect 14544 2916 14596 2922
rect 15002 2887 15058 2896
rect 14544 2858 14596 2864
rect 14668 2204 14964 2224
rect 14724 2202 14748 2204
rect 14804 2202 14828 2204
rect 14884 2202 14908 2204
rect 14746 2150 14748 2202
rect 14810 2150 14822 2202
rect 14884 2150 14886 2202
rect 14724 2148 14748 2150
rect 14804 2148 14828 2150
rect 14884 2148 14908 2150
rect 14668 2128 14964 2148
rect 15108 1578 15136 3062
rect 15384 3058 15412 3538
rect 15556 3528 15608 3534
rect 15556 3470 15608 3476
rect 15568 3194 15596 3470
rect 15556 3188 15608 3194
rect 15556 3130 15608 3136
rect 15372 3052 15424 3058
rect 15372 2994 15424 3000
rect 15568 2582 15596 3130
rect 15752 2802 15780 10095
rect 15832 10066 15884 10072
rect 15924 9376 15976 9382
rect 15924 9318 15976 9324
rect 15832 6860 15884 6866
rect 15832 6802 15884 6808
rect 15844 6254 15872 6802
rect 15936 6361 15964 9318
rect 15922 6352 15978 6361
rect 15922 6287 15978 6296
rect 15832 6248 15884 6254
rect 15830 6216 15832 6225
rect 15884 6216 15886 6225
rect 15830 6151 15886 6160
rect 16028 3738 16056 11562
rect 16120 10810 16148 17303
rect 19334 16892 19630 16912
rect 19390 16890 19414 16892
rect 19470 16890 19494 16892
rect 19550 16890 19574 16892
rect 19412 16838 19414 16890
rect 19476 16838 19488 16890
rect 19550 16838 19552 16890
rect 19390 16836 19414 16838
rect 19470 16836 19494 16838
rect 19550 16836 19574 16838
rect 19334 16816 19630 16836
rect 18222 16688 18278 16697
rect 18222 16623 18278 16632
rect 18236 16114 18264 16623
rect 18224 16108 18276 16114
rect 18224 16050 18276 16056
rect 18868 15904 18920 15910
rect 18868 15846 18920 15852
rect 18590 13968 18646 13977
rect 18590 13903 18592 13912
rect 18644 13903 18646 13912
rect 18592 13874 18644 13880
rect 18776 13864 18828 13870
rect 18776 13806 18828 13812
rect 16658 12880 16714 12889
rect 16658 12815 16714 12824
rect 16476 12640 16528 12646
rect 16476 12582 16528 12588
rect 16384 12300 16436 12306
rect 16384 12242 16436 12248
rect 16396 11830 16424 12242
rect 16384 11824 16436 11830
rect 16384 11766 16436 11772
rect 16198 11112 16254 11121
rect 16198 11047 16254 11056
rect 16108 10804 16160 10810
rect 16108 10746 16160 10752
rect 16212 9654 16240 11047
rect 16488 10606 16516 12582
rect 16672 12374 16700 12815
rect 18590 12744 18646 12753
rect 18590 12679 18592 12688
rect 18644 12679 18646 12688
rect 18592 12650 18644 12656
rect 18500 12436 18552 12442
rect 18500 12378 18552 12384
rect 16660 12368 16712 12374
rect 16660 12310 16712 12316
rect 17856 12368 17908 12374
rect 17856 12310 17908 12316
rect 17868 11762 17896 12310
rect 17856 11756 17908 11762
rect 17856 11698 17908 11704
rect 17868 11558 17896 11698
rect 17856 11552 17908 11558
rect 17856 11494 17908 11500
rect 18316 11552 18368 11558
rect 18316 11494 18368 11500
rect 17868 11354 17896 11494
rect 17856 11348 17908 11354
rect 17856 11290 17908 11296
rect 17396 11280 17448 11286
rect 17396 11222 17448 11228
rect 16568 11212 16620 11218
rect 16568 11154 16620 11160
rect 16580 10606 16608 11154
rect 16660 11008 16712 11014
rect 16660 10950 16712 10956
rect 16842 10976 16898 10985
rect 16672 10674 16700 10950
rect 16842 10911 16898 10920
rect 16660 10668 16712 10674
rect 16660 10610 16712 10616
rect 16476 10600 16528 10606
rect 16476 10542 16528 10548
rect 16568 10600 16620 10606
rect 16568 10542 16620 10548
rect 16580 9926 16608 10542
rect 16660 10464 16712 10470
rect 16660 10406 16712 10412
rect 16568 9920 16620 9926
rect 16568 9862 16620 9868
rect 16200 9648 16252 9654
rect 16200 9590 16252 9596
rect 16580 9586 16608 9862
rect 16672 9722 16700 10406
rect 16660 9716 16712 9722
rect 16660 9658 16712 9664
rect 16568 9580 16620 9586
rect 16568 9522 16620 9528
rect 16580 9178 16608 9522
rect 16660 9376 16712 9382
rect 16660 9318 16712 9324
rect 16568 9172 16620 9178
rect 16568 9114 16620 9120
rect 16672 9110 16700 9318
rect 16660 9104 16712 9110
rect 16660 9046 16712 9052
rect 16752 9036 16804 9042
rect 16752 8978 16804 8984
rect 16764 8362 16792 8978
rect 16752 8356 16804 8362
rect 16752 8298 16804 8304
rect 16384 8288 16436 8294
rect 16384 8230 16436 8236
rect 16396 8090 16424 8230
rect 16384 8084 16436 8090
rect 16384 8026 16436 8032
rect 16764 7478 16792 8298
rect 16752 7472 16804 7478
rect 16474 7440 16530 7449
rect 16752 7414 16804 7420
rect 16474 7375 16530 7384
rect 16108 6928 16160 6934
rect 16108 6870 16160 6876
rect 16120 6118 16148 6870
rect 16488 6866 16516 7375
rect 16476 6860 16528 6866
rect 16528 6820 16608 6848
rect 16476 6802 16528 6808
rect 16580 6168 16608 6820
rect 16660 6180 16712 6186
rect 16580 6140 16660 6168
rect 16108 6112 16160 6118
rect 16108 6054 16160 6060
rect 16120 4865 16148 6054
rect 16384 5772 16436 5778
rect 16384 5714 16436 5720
rect 16198 5536 16254 5545
rect 16198 5471 16254 5480
rect 16106 4856 16162 4865
rect 16212 4826 16240 5471
rect 16396 5137 16424 5714
rect 16580 5710 16608 6140
rect 16660 6122 16712 6128
rect 16752 6112 16804 6118
rect 16752 6054 16804 6060
rect 16476 5704 16528 5710
rect 16476 5646 16528 5652
rect 16568 5704 16620 5710
rect 16568 5646 16620 5652
rect 16382 5128 16438 5137
rect 16382 5063 16438 5072
rect 16106 4791 16162 4800
rect 16200 4820 16252 4826
rect 16200 4762 16252 4768
rect 16384 4684 16436 4690
rect 16384 4626 16436 4632
rect 16290 4312 16346 4321
rect 16290 4247 16346 4256
rect 16304 4146 16332 4247
rect 16292 4140 16344 4146
rect 16292 4082 16344 4088
rect 16200 3936 16252 3942
rect 16200 3878 16252 3884
rect 16016 3732 16068 3738
rect 16016 3674 16068 3680
rect 16028 2990 16056 3674
rect 16016 2984 16068 2990
rect 16016 2926 16068 2932
rect 15752 2774 15872 2802
rect 15556 2576 15608 2582
rect 15556 2518 15608 2524
rect 15844 2428 15872 2774
rect 14924 1550 15136 1578
rect 15568 2400 15872 2428
rect 14924 480 14952 1550
rect 15568 480 15596 2400
rect 16212 480 16240 3878
rect 16396 3738 16424 4626
rect 16488 4554 16516 5646
rect 16660 5092 16712 5098
rect 16660 5034 16712 5040
rect 16568 5024 16620 5030
rect 16568 4966 16620 4972
rect 16580 4622 16608 4966
rect 16568 4616 16620 4622
rect 16568 4558 16620 4564
rect 16476 4548 16528 4554
rect 16476 4490 16528 4496
rect 16580 4282 16608 4558
rect 16568 4276 16620 4282
rect 16568 4218 16620 4224
rect 16384 3732 16436 3738
rect 16384 3674 16436 3680
rect 16384 3596 16436 3602
rect 16384 3538 16436 3544
rect 16396 3233 16424 3538
rect 16382 3224 16438 3233
rect 16382 3159 16384 3168
rect 16436 3159 16438 3168
rect 16384 3130 16436 3136
rect 16672 2802 16700 5034
rect 16764 2961 16792 6054
rect 16856 5098 16884 10911
rect 17408 10606 17436 11222
rect 18328 11121 18356 11494
rect 18314 11112 18370 11121
rect 18314 11047 18316 11056
rect 18368 11047 18370 11056
rect 18316 11018 18368 11024
rect 17672 10668 17724 10674
rect 17672 10610 17724 10616
rect 17396 10600 17448 10606
rect 17396 10542 17448 10548
rect 17408 10266 17436 10542
rect 17396 10260 17448 10266
rect 17396 10202 17448 10208
rect 17408 9194 17436 10202
rect 17580 9988 17632 9994
rect 17580 9930 17632 9936
rect 17486 9480 17542 9489
rect 17486 9415 17488 9424
rect 17540 9415 17542 9424
rect 17488 9386 17540 9392
rect 17224 9166 17436 9194
rect 17488 9172 17540 9178
rect 17224 8906 17252 9166
rect 17592 9160 17620 9930
rect 17684 9178 17712 10610
rect 17764 10464 17816 10470
rect 17764 10406 17816 10412
rect 17540 9132 17620 9160
rect 17672 9172 17724 9178
rect 17488 9114 17540 9120
rect 17672 9114 17724 9120
rect 17396 9104 17448 9110
rect 17396 9046 17448 9052
rect 17212 8900 17264 8906
rect 17212 8842 17264 8848
rect 17408 8634 17436 9046
rect 17396 8628 17448 8634
rect 17396 8570 17448 8576
rect 17776 8090 17804 10406
rect 17856 10056 17908 10062
rect 17856 9998 17908 10004
rect 17868 9625 17896 9998
rect 18316 9920 18368 9926
rect 18316 9862 18368 9868
rect 18328 9654 18356 9862
rect 18512 9704 18540 12378
rect 18684 12300 18736 12306
rect 18684 12242 18736 12248
rect 18696 11694 18724 12242
rect 18684 11688 18736 11694
rect 18684 11630 18736 11636
rect 18696 10674 18724 11630
rect 18684 10668 18736 10674
rect 18684 10610 18736 10616
rect 18420 9676 18540 9704
rect 18316 9648 18368 9654
rect 17854 9616 17910 9625
rect 18420 9636 18448 9676
rect 18420 9608 18540 9636
rect 18316 9590 18368 9596
rect 17854 9551 17910 9560
rect 17948 9580 18000 9586
rect 17948 9522 18000 9528
rect 17854 9480 17910 9489
rect 17854 9415 17910 9424
rect 17868 8129 17896 9415
rect 17960 9110 17988 9522
rect 18512 9382 18540 9608
rect 18592 9444 18644 9450
rect 18592 9386 18644 9392
rect 18224 9376 18276 9382
rect 18224 9318 18276 9324
rect 18316 9376 18368 9382
rect 18316 9318 18368 9324
rect 18500 9376 18552 9382
rect 18500 9318 18552 9324
rect 17948 9104 18000 9110
rect 17948 9046 18000 9052
rect 17946 8800 18002 8809
rect 17946 8735 18002 8744
rect 17854 8120 17910 8129
rect 17764 8084 17816 8090
rect 17854 8055 17910 8064
rect 17764 8026 17816 8032
rect 17212 7744 17264 7750
rect 17212 7686 17264 7692
rect 17120 7200 17172 7206
rect 17120 7142 17172 7148
rect 17132 6769 17160 7142
rect 17118 6760 17174 6769
rect 17118 6695 17174 6704
rect 17120 6656 17172 6662
rect 17120 6598 17172 6604
rect 17132 6118 17160 6598
rect 17120 6112 17172 6118
rect 17120 6054 17172 6060
rect 17132 5710 17160 6054
rect 17120 5704 17172 5710
rect 17120 5646 17172 5652
rect 17026 5264 17082 5273
rect 17026 5199 17082 5208
rect 16934 5128 16990 5137
rect 16844 5092 16896 5098
rect 16934 5063 16990 5072
rect 16844 5034 16896 5040
rect 16842 4992 16898 5001
rect 16842 4927 16898 4936
rect 16856 3670 16884 4927
rect 16948 4185 16976 5063
rect 16934 4176 16990 4185
rect 16934 4111 16990 4120
rect 17040 3738 17068 5199
rect 17224 4826 17252 7686
rect 17672 7200 17724 7206
rect 17672 7142 17724 7148
rect 17302 6760 17358 6769
rect 17302 6695 17358 6704
rect 17316 6458 17344 6695
rect 17304 6452 17356 6458
rect 17304 6394 17356 6400
rect 17488 6180 17540 6186
rect 17488 6122 17540 6128
rect 17304 5772 17356 5778
rect 17304 5714 17356 5720
rect 17316 5409 17344 5714
rect 17302 5400 17358 5409
rect 17500 5370 17528 6122
rect 17580 5908 17632 5914
rect 17684 5896 17712 7142
rect 17776 7002 17804 8026
rect 17856 7948 17908 7954
rect 17856 7890 17908 7896
rect 17764 6996 17816 7002
rect 17764 6938 17816 6944
rect 17868 6730 17896 7890
rect 17856 6724 17908 6730
rect 17856 6666 17908 6672
rect 17632 5868 17712 5896
rect 17580 5850 17632 5856
rect 17302 5335 17304 5344
rect 17356 5335 17358 5344
rect 17488 5364 17540 5370
rect 17304 5306 17356 5312
rect 17488 5306 17540 5312
rect 17212 4820 17264 4826
rect 17212 4762 17264 4768
rect 17500 4758 17528 5306
rect 17684 5166 17712 5868
rect 17868 5846 17896 6666
rect 17856 5840 17908 5846
rect 17856 5782 17908 5788
rect 17764 5568 17816 5574
rect 17764 5510 17816 5516
rect 17776 5234 17804 5510
rect 17868 5302 17896 5782
rect 17856 5296 17908 5302
rect 17856 5238 17908 5244
rect 17764 5228 17816 5234
rect 17764 5170 17816 5176
rect 17672 5160 17724 5166
rect 17672 5102 17724 5108
rect 17488 4752 17540 4758
rect 17488 4694 17540 4700
rect 17672 4752 17724 4758
rect 17672 4694 17724 4700
rect 17120 4684 17172 4690
rect 17120 4626 17172 4632
rect 17132 3942 17160 4626
rect 17500 4622 17528 4694
rect 17488 4616 17540 4622
rect 17488 4558 17540 4564
rect 17210 4448 17266 4457
rect 17210 4383 17266 4392
rect 17120 3936 17172 3942
rect 17120 3878 17172 3884
rect 17132 3777 17160 3878
rect 17118 3768 17174 3777
rect 17028 3732 17080 3738
rect 17118 3703 17174 3712
rect 17028 3674 17080 3680
rect 16844 3664 16896 3670
rect 16844 3606 16896 3612
rect 16856 3194 16884 3606
rect 16844 3188 16896 3194
rect 16844 3130 16896 3136
rect 17040 3126 17068 3674
rect 17224 3534 17252 4383
rect 17304 4140 17356 4146
rect 17304 4082 17356 4088
rect 17212 3528 17264 3534
rect 17212 3470 17264 3476
rect 17028 3120 17080 3126
rect 17028 3062 17080 3068
rect 16750 2952 16806 2961
rect 16750 2887 16806 2896
rect 16672 2774 16792 2802
rect 16566 2680 16622 2689
rect 16764 2666 16792 2774
rect 16764 2638 16884 2666
rect 17224 2650 17252 3470
rect 17316 3398 17344 4082
rect 17488 3936 17540 3942
rect 17488 3878 17540 3884
rect 17304 3392 17356 3398
rect 17304 3334 17356 3340
rect 17316 2922 17344 3334
rect 17500 3097 17528 3878
rect 17684 3738 17712 4694
rect 17960 4321 17988 8735
rect 18236 8242 18264 9318
rect 18144 8214 18264 8242
rect 18144 7206 18172 8214
rect 18328 7886 18356 9318
rect 18500 9172 18552 9178
rect 18500 9114 18552 9120
rect 18512 8634 18540 9114
rect 18500 8628 18552 8634
rect 18500 8570 18552 8576
rect 18512 8430 18540 8570
rect 18604 8498 18632 9386
rect 18592 8492 18644 8498
rect 18592 8434 18644 8440
rect 18500 8424 18552 8430
rect 18500 8366 18552 8372
rect 18316 7880 18368 7886
rect 18316 7822 18368 7828
rect 18592 7880 18644 7886
rect 18592 7822 18644 7828
rect 18316 7744 18368 7750
rect 18222 7712 18278 7721
rect 18316 7686 18368 7692
rect 18222 7647 18278 7656
rect 18132 7200 18184 7206
rect 18132 7142 18184 7148
rect 18236 6440 18264 7647
rect 18328 7449 18356 7686
rect 18314 7440 18370 7449
rect 18314 7375 18316 7384
rect 18368 7375 18370 7384
rect 18316 7346 18368 7352
rect 18498 7304 18554 7313
rect 18498 7239 18554 7248
rect 18316 6792 18368 6798
rect 18316 6734 18368 6740
rect 18144 6412 18264 6440
rect 18040 6112 18092 6118
rect 18040 6054 18092 6060
rect 18052 5273 18080 6054
rect 18038 5264 18094 5273
rect 18038 5199 18094 5208
rect 17946 4312 18002 4321
rect 17946 4247 18002 4256
rect 18144 4128 18172 6412
rect 18328 5352 18356 6734
rect 18512 6458 18540 7239
rect 18604 6798 18632 7822
rect 18592 6792 18644 6798
rect 18592 6734 18644 6740
rect 18788 6730 18816 13806
rect 18880 12442 18908 15846
rect 19334 15804 19630 15824
rect 19390 15802 19414 15804
rect 19470 15802 19494 15804
rect 19550 15802 19574 15804
rect 19412 15750 19414 15802
rect 19476 15750 19488 15802
rect 19550 15750 19552 15802
rect 19390 15748 19414 15750
rect 19470 15748 19494 15750
rect 19550 15748 19574 15750
rect 19334 15728 19630 15748
rect 19334 14716 19630 14736
rect 19390 14714 19414 14716
rect 19470 14714 19494 14716
rect 19550 14714 19574 14716
rect 19412 14662 19414 14714
rect 19476 14662 19488 14714
rect 19550 14662 19552 14714
rect 19390 14660 19414 14662
rect 19470 14660 19494 14662
rect 19550 14660 19574 14662
rect 19334 14640 19630 14660
rect 20432 13728 20484 13734
rect 20432 13670 20484 13676
rect 19334 13628 19630 13648
rect 19390 13626 19414 13628
rect 19470 13626 19494 13628
rect 19550 13626 19574 13628
rect 19412 13574 19414 13626
rect 19476 13574 19488 13626
rect 19550 13574 19552 13626
rect 19390 13572 19414 13574
rect 19470 13572 19494 13574
rect 19550 13572 19574 13574
rect 19334 13552 19630 13572
rect 19236 13320 19288 13326
rect 19236 13262 19288 13268
rect 18958 13152 19014 13161
rect 18958 13087 19014 13096
rect 18972 12986 19000 13087
rect 18960 12980 19012 12986
rect 18960 12922 19012 12928
rect 19144 12844 19196 12850
rect 19144 12786 19196 12792
rect 18958 12744 19014 12753
rect 18958 12679 19014 12688
rect 18868 12436 18920 12442
rect 18868 12378 18920 12384
rect 18868 12096 18920 12102
rect 18868 12038 18920 12044
rect 18880 11286 18908 12038
rect 18972 11354 19000 12679
rect 18960 11348 19012 11354
rect 18960 11290 19012 11296
rect 19052 11348 19104 11354
rect 19052 11290 19104 11296
rect 18868 11280 18920 11286
rect 18868 11222 18920 11228
rect 18880 10606 18908 11222
rect 18960 10804 19012 10810
rect 19064 10792 19092 11290
rect 19012 10764 19092 10792
rect 18960 10746 19012 10752
rect 18868 10600 18920 10606
rect 18868 10542 18920 10548
rect 18880 10130 18908 10542
rect 19156 10198 19184 12786
rect 19248 11354 19276 13262
rect 19420 13184 19472 13190
rect 19420 13126 19472 13132
rect 19432 12850 19460 13126
rect 19420 12844 19472 12850
rect 19420 12786 19472 12792
rect 19788 12776 19840 12782
rect 19788 12718 19840 12724
rect 19334 12540 19630 12560
rect 19390 12538 19414 12540
rect 19470 12538 19494 12540
rect 19550 12538 19574 12540
rect 19412 12486 19414 12538
rect 19476 12486 19488 12538
rect 19550 12486 19552 12538
rect 19390 12484 19414 12486
rect 19470 12484 19494 12486
rect 19550 12484 19574 12486
rect 19334 12464 19630 12484
rect 19604 12096 19656 12102
rect 19604 12038 19656 12044
rect 19616 11762 19644 12038
rect 19604 11756 19656 11762
rect 19604 11698 19656 11704
rect 19696 11552 19748 11558
rect 19696 11494 19748 11500
rect 19334 11452 19630 11472
rect 19390 11450 19414 11452
rect 19470 11450 19494 11452
rect 19550 11450 19574 11452
rect 19412 11398 19414 11450
rect 19476 11398 19488 11450
rect 19550 11398 19552 11450
rect 19390 11396 19414 11398
rect 19470 11396 19494 11398
rect 19550 11396 19574 11398
rect 19334 11376 19630 11396
rect 19236 11348 19288 11354
rect 19236 11290 19288 11296
rect 19512 11144 19564 11150
rect 19708 11132 19736 11494
rect 19564 11104 19736 11132
rect 19512 11086 19564 11092
rect 19524 10538 19552 11086
rect 19512 10532 19564 10538
rect 19512 10474 19564 10480
rect 19334 10364 19630 10384
rect 19390 10362 19414 10364
rect 19470 10362 19494 10364
rect 19550 10362 19574 10364
rect 19412 10310 19414 10362
rect 19476 10310 19488 10362
rect 19550 10310 19552 10362
rect 19390 10308 19414 10310
rect 19470 10308 19494 10310
rect 19550 10308 19574 10310
rect 19334 10288 19630 10308
rect 19144 10192 19196 10198
rect 19144 10134 19196 10140
rect 18868 10124 18920 10130
rect 18868 10066 18920 10072
rect 19052 10124 19104 10130
rect 19052 10066 19104 10072
rect 18960 9920 19012 9926
rect 18960 9862 19012 9868
rect 18972 9518 19000 9862
rect 18960 9512 19012 9518
rect 18960 9454 19012 9460
rect 18868 9376 18920 9382
rect 18866 9344 18868 9353
rect 18920 9344 18922 9353
rect 19064 9330 19092 10066
rect 18922 9302 19092 9330
rect 18866 9279 18922 9288
rect 19156 8838 19184 10134
rect 19800 9518 19828 12718
rect 20444 11354 20472 13670
rect 20628 13530 20656 19110
rect 22468 17377 22496 19110
rect 23192 18216 23244 18222
rect 23112 18164 23192 18170
rect 23112 18158 23244 18164
rect 23112 18142 23232 18158
rect 22454 17368 22510 17377
rect 22454 17303 22510 17312
rect 21534 16552 21590 16561
rect 21534 16487 21590 16496
rect 20984 14408 21036 14414
rect 20984 14350 21036 14356
rect 20996 13530 21024 14350
rect 20616 13524 20668 13530
rect 20616 13466 20668 13472
rect 20984 13524 21036 13530
rect 20984 13466 21036 13472
rect 20524 13184 20576 13190
rect 20522 13152 20524 13161
rect 20576 13152 20578 13161
rect 20522 13087 20578 13096
rect 20996 12986 21024 13466
rect 21352 13320 21404 13326
rect 21352 13262 21404 13268
rect 21074 13016 21130 13025
rect 20984 12980 21036 12986
rect 21074 12951 21130 12960
rect 20984 12922 21036 12928
rect 21088 12782 21116 12951
rect 21168 12844 21220 12850
rect 21168 12786 21220 12792
rect 21076 12776 21128 12782
rect 21076 12718 21128 12724
rect 20524 12640 20576 12646
rect 20524 12582 20576 12588
rect 20432 11348 20484 11354
rect 20432 11290 20484 11296
rect 19880 11212 19932 11218
rect 19880 11154 19932 11160
rect 19892 10266 19920 11154
rect 20444 10810 20472 11290
rect 20536 11286 20564 12582
rect 21180 12306 21208 12786
rect 21364 12442 21392 13262
rect 21352 12436 21404 12442
rect 21352 12378 21404 12384
rect 21168 12300 21220 12306
rect 21168 12242 21220 12248
rect 21180 11898 21208 12242
rect 21168 11892 21220 11898
rect 21168 11834 21220 11840
rect 20614 11656 20670 11665
rect 20614 11591 20670 11600
rect 20524 11280 20576 11286
rect 20524 11222 20576 11228
rect 20432 10804 20484 10810
rect 20432 10746 20484 10752
rect 20536 10266 20564 11222
rect 20628 11082 20656 11591
rect 21168 11144 21220 11150
rect 21168 11086 21220 11092
rect 20616 11076 20668 11082
rect 20616 11018 20668 11024
rect 21180 10810 21208 11086
rect 21168 10804 21220 10810
rect 21168 10746 21220 10752
rect 19880 10260 19932 10266
rect 19880 10202 19932 10208
rect 20524 10260 20576 10266
rect 20524 10202 20576 10208
rect 21168 10124 21220 10130
rect 21168 10066 21220 10072
rect 19604 9512 19656 9518
rect 19788 9512 19840 9518
rect 19656 9460 19736 9466
rect 19604 9454 19736 9460
rect 19788 9454 19840 9460
rect 19616 9438 19736 9454
rect 19334 9276 19630 9296
rect 19390 9274 19414 9276
rect 19470 9274 19494 9276
rect 19550 9274 19574 9276
rect 19412 9222 19414 9274
rect 19476 9222 19488 9274
rect 19550 9222 19552 9274
rect 19390 9220 19414 9222
rect 19470 9220 19494 9222
rect 19550 9220 19574 9222
rect 19334 9200 19630 9220
rect 19144 8832 19196 8838
rect 19144 8774 19196 8780
rect 18958 8392 19014 8401
rect 18958 8327 19014 8336
rect 18972 7857 19000 8327
rect 19334 8188 19630 8208
rect 19390 8186 19414 8188
rect 19470 8186 19494 8188
rect 19550 8186 19574 8188
rect 19412 8134 19414 8186
rect 19476 8134 19488 8186
rect 19550 8134 19552 8186
rect 19390 8132 19414 8134
rect 19470 8132 19494 8134
rect 19550 8132 19574 8134
rect 19334 8112 19630 8132
rect 18958 7848 19014 7857
rect 18958 7783 19014 7792
rect 19236 7812 19288 7818
rect 19236 7754 19288 7760
rect 19144 7472 19196 7478
rect 19144 7414 19196 7420
rect 18868 7200 18920 7206
rect 18868 7142 18920 7148
rect 18880 6934 18908 7142
rect 18868 6928 18920 6934
rect 18868 6870 18920 6876
rect 18776 6724 18828 6730
rect 18776 6666 18828 6672
rect 18684 6656 18736 6662
rect 18684 6598 18736 6604
rect 18500 6452 18552 6458
rect 18500 6394 18552 6400
rect 18512 6254 18540 6394
rect 18500 6248 18552 6254
rect 18500 6190 18552 6196
rect 18696 5370 18724 6598
rect 18774 6352 18830 6361
rect 18774 6287 18830 6296
rect 18052 4100 18172 4128
rect 18236 5324 18356 5352
rect 18684 5364 18736 5370
rect 17764 3936 17816 3942
rect 17764 3878 17816 3884
rect 17672 3732 17724 3738
rect 17672 3674 17724 3680
rect 17776 3670 17804 3878
rect 17764 3664 17816 3670
rect 17764 3606 17816 3612
rect 17486 3088 17542 3097
rect 17486 3023 17542 3032
rect 17764 2984 17816 2990
rect 17764 2926 17816 2932
rect 17304 2916 17356 2922
rect 17304 2858 17356 2864
rect 16566 2615 16568 2624
rect 16620 2615 16622 2624
rect 16568 2586 16620 2592
rect 16856 480 16884 2638
rect 17212 2644 17264 2650
rect 17212 2586 17264 2592
rect 17776 2446 17804 2926
rect 17764 2440 17816 2446
rect 17764 2382 17816 2388
rect 18052 610 18080 4100
rect 18130 4040 18186 4049
rect 18130 3975 18132 3984
rect 18184 3975 18186 3984
rect 18132 3946 18184 3952
rect 18144 3602 18172 3946
rect 18236 3738 18264 5324
rect 18684 5306 18736 5312
rect 18316 5228 18368 5234
rect 18316 5170 18368 5176
rect 18328 4826 18356 5170
rect 18316 4820 18368 4826
rect 18316 4762 18368 4768
rect 18592 4752 18644 4758
rect 18592 4694 18644 4700
rect 18604 4486 18632 4694
rect 18788 4570 18816 6287
rect 18960 6248 19012 6254
rect 18960 6190 19012 6196
rect 18972 5658 19000 6190
rect 19052 6180 19104 6186
rect 19052 6122 19104 6128
rect 19064 5914 19092 6122
rect 19052 5908 19104 5914
rect 19052 5850 19104 5856
rect 18972 5630 19092 5658
rect 19064 5370 19092 5630
rect 19156 5545 19184 7414
rect 19248 7002 19276 7754
rect 19334 7100 19630 7120
rect 19390 7098 19414 7100
rect 19470 7098 19494 7100
rect 19550 7098 19574 7100
rect 19412 7046 19414 7098
rect 19476 7046 19488 7098
rect 19550 7046 19552 7098
rect 19390 7044 19414 7046
rect 19470 7044 19494 7046
rect 19550 7044 19574 7046
rect 19334 7024 19630 7044
rect 19236 6996 19288 7002
rect 19236 6938 19288 6944
rect 19420 6792 19472 6798
rect 19420 6734 19472 6740
rect 19432 6186 19460 6734
rect 19420 6180 19472 6186
rect 19420 6122 19472 6128
rect 19334 6012 19630 6032
rect 19390 6010 19414 6012
rect 19470 6010 19494 6012
rect 19550 6010 19574 6012
rect 19412 5958 19414 6010
rect 19476 5958 19488 6010
rect 19550 5958 19552 6010
rect 19390 5956 19414 5958
rect 19470 5956 19494 5958
rect 19550 5956 19574 5958
rect 19334 5936 19630 5956
rect 19708 5681 19736 9438
rect 19800 9178 19828 9454
rect 20340 9444 20392 9450
rect 20340 9386 20392 9392
rect 20352 9330 20380 9386
rect 20352 9302 20472 9330
rect 19788 9172 19840 9178
rect 19788 9114 19840 9120
rect 19800 8634 19828 9114
rect 19788 8628 19840 8634
rect 19788 8570 19840 8576
rect 20340 8560 20392 8566
rect 20340 8502 20392 8508
rect 20352 8090 20380 8502
rect 20340 8084 20392 8090
rect 20340 8026 20392 8032
rect 20444 8022 20472 9302
rect 21180 9178 21208 10066
rect 21260 10056 21312 10062
rect 21260 9998 21312 10004
rect 21272 9450 21300 9998
rect 21364 9654 21392 12378
rect 21352 9648 21404 9654
rect 21352 9590 21404 9596
rect 21260 9444 21312 9450
rect 21260 9386 21312 9392
rect 21168 9172 21220 9178
rect 21168 9114 21220 9120
rect 20984 9036 21036 9042
rect 20628 8974 20656 9005
rect 20984 8978 21036 8984
rect 20616 8968 20668 8974
rect 20614 8936 20616 8945
rect 20668 8936 20670 8945
rect 20614 8871 20670 8880
rect 20800 8900 20852 8906
rect 20628 8634 20656 8871
rect 20800 8842 20852 8848
rect 20616 8628 20668 8634
rect 20616 8570 20668 8576
rect 20432 8016 20484 8022
rect 20432 7958 20484 7964
rect 19880 7880 19932 7886
rect 19880 7822 19932 7828
rect 19786 7168 19842 7177
rect 19786 7103 19842 7112
rect 19510 5672 19566 5681
rect 19510 5607 19566 5616
rect 19694 5672 19750 5681
rect 19694 5607 19750 5616
rect 19142 5536 19198 5545
rect 19142 5471 19198 5480
rect 19052 5364 19104 5370
rect 19052 5306 19104 5312
rect 19524 5166 19552 5607
rect 19512 5160 19564 5166
rect 19512 5102 19564 5108
rect 19144 5092 19196 5098
rect 19144 5034 19196 5040
rect 18960 4820 19012 4826
rect 18960 4762 19012 4768
rect 18696 4542 18816 4570
rect 18592 4480 18644 4486
rect 18592 4422 18644 4428
rect 18604 4146 18632 4422
rect 18592 4140 18644 4146
rect 18592 4082 18644 4088
rect 18224 3732 18276 3738
rect 18224 3674 18276 3680
rect 18696 3618 18724 4542
rect 18776 4480 18828 4486
rect 18776 4422 18828 4428
rect 18788 3738 18816 4422
rect 18866 4312 18922 4321
rect 18866 4247 18922 4256
rect 18776 3732 18828 3738
rect 18776 3674 18828 3680
rect 18132 3596 18184 3602
rect 18132 3538 18184 3544
rect 18604 3590 18724 3618
rect 18314 2544 18370 2553
rect 18314 2479 18316 2488
rect 18368 2479 18370 2488
rect 18316 2450 18368 2456
rect 18604 610 18632 3590
rect 18684 3528 18736 3534
rect 18682 3496 18684 3505
rect 18736 3496 18738 3505
rect 18682 3431 18738 3440
rect 18696 3194 18724 3431
rect 18684 3188 18736 3194
rect 18684 3130 18736 3136
rect 17488 604 17540 610
rect 17488 546 17540 552
rect 18040 604 18092 610
rect 18040 546 18092 552
rect 18132 604 18184 610
rect 18132 546 18184 552
rect 18592 604 18644 610
rect 18592 546 18644 552
rect 17500 480 17528 546
rect 18144 480 18172 546
rect 18880 480 18908 4247
rect 18972 4146 19000 4762
rect 19156 4622 19184 5034
rect 19236 5024 19288 5030
rect 19236 4966 19288 4972
rect 19248 4758 19276 4966
rect 19334 4924 19630 4944
rect 19390 4922 19414 4924
rect 19470 4922 19494 4924
rect 19550 4922 19574 4924
rect 19412 4870 19414 4922
rect 19476 4870 19488 4922
rect 19550 4870 19552 4922
rect 19390 4868 19414 4870
rect 19470 4868 19494 4870
rect 19550 4868 19574 4870
rect 19334 4848 19630 4868
rect 19236 4752 19288 4758
rect 19236 4694 19288 4700
rect 19144 4616 19196 4622
rect 19144 4558 19196 4564
rect 19052 4548 19104 4554
rect 19052 4490 19104 4496
rect 18960 4140 19012 4146
rect 18960 4082 19012 4088
rect 19064 3754 19092 4490
rect 18972 3726 19092 3754
rect 18972 3670 19000 3726
rect 19156 3670 19184 4558
rect 19236 4004 19288 4010
rect 19236 3946 19288 3952
rect 18960 3664 19012 3670
rect 18960 3606 19012 3612
rect 19144 3664 19196 3670
rect 19144 3606 19196 3612
rect 19144 3392 19196 3398
rect 19144 3334 19196 3340
rect 19052 2916 19104 2922
rect 19052 2858 19104 2864
rect 19064 2650 19092 2858
rect 19156 2825 19184 3334
rect 19248 3233 19276 3946
rect 19800 3942 19828 7103
rect 19892 5914 19920 7822
rect 20812 7750 20840 8842
rect 20892 8832 20944 8838
rect 20892 8774 20944 8780
rect 20904 8242 20932 8774
rect 20996 8401 21024 8978
rect 20982 8392 21038 8401
rect 20982 8327 20984 8336
rect 21036 8327 21038 8336
rect 20984 8298 21036 8304
rect 20904 8214 21024 8242
rect 20800 7744 20852 7750
rect 20800 7686 20852 7692
rect 20892 7744 20944 7750
rect 20892 7686 20944 7692
rect 20812 7546 20840 7686
rect 20800 7540 20852 7546
rect 20800 7482 20852 7488
rect 19970 7440 20026 7449
rect 19970 7375 19972 7384
rect 20024 7375 20026 7384
rect 20156 7404 20208 7410
rect 19972 7346 20024 7352
rect 20156 7346 20208 7352
rect 20064 7336 20116 7342
rect 20064 7278 20116 7284
rect 19972 7268 20024 7274
rect 19972 7210 20024 7216
rect 19880 5908 19932 5914
rect 19880 5850 19932 5856
rect 19892 5166 19920 5850
rect 19880 5160 19932 5166
rect 19880 5102 19932 5108
rect 19880 5024 19932 5030
rect 19880 4966 19932 4972
rect 19892 4185 19920 4966
rect 19984 4865 20012 7210
rect 20076 5098 20104 7278
rect 20168 7002 20196 7346
rect 20904 7342 20932 7686
rect 20892 7336 20944 7342
rect 20892 7278 20944 7284
rect 20156 6996 20208 7002
rect 20156 6938 20208 6944
rect 20064 5092 20116 5098
rect 20064 5034 20116 5040
rect 19970 4856 20026 4865
rect 19970 4791 20026 4800
rect 19984 4758 20012 4791
rect 19972 4752 20024 4758
rect 19972 4694 20024 4700
rect 20168 4457 20196 6938
rect 20996 6866 21024 8214
rect 21272 7546 21300 9386
rect 21364 7954 21392 9590
rect 21548 8634 21576 16487
rect 22732 15564 22784 15570
rect 22732 15506 22784 15512
rect 22744 14822 22772 15506
rect 23112 14929 23140 18142
rect 23098 14920 23154 14929
rect 23098 14855 23154 14864
rect 22732 14816 22784 14822
rect 22732 14758 22784 14764
rect 21812 13864 21864 13870
rect 21640 13812 21812 13818
rect 21640 13806 21864 13812
rect 21640 13790 21852 13806
rect 21640 10266 21668 13790
rect 21904 13728 21956 13734
rect 21904 13670 21956 13676
rect 21812 12640 21864 12646
rect 21812 12582 21864 12588
rect 21718 11792 21774 11801
rect 21718 11727 21774 11736
rect 21732 10742 21760 11727
rect 21720 10736 21772 10742
rect 21720 10678 21772 10684
rect 21628 10260 21680 10266
rect 21628 10202 21680 10208
rect 21720 10056 21772 10062
rect 21720 9998 21772 10004
rect 21732 9382 21760 9998
rect 21720 9376 21772 9382
rect 21720 9318 21772 9324
rect 21628 8900 21680 8906
rect 21628 8842 21680 8848
rect 21536 8628 21588 8634
rect 21536 8570 21588 8576
rect 21640 8022 21668 8842
rect 21732 8786 21760 9318
rect 21824 9178 21852 12582
rect 21916 10810 21944 13670
rect 22180 13184 22232 13190
rect 22180 13126 22232 13132
rect 21996 12164 22048 12170
rect 21996 12106 22048 12112
rect 22008 11150 22036 12106
rect 22088 12096 22140 12102
rect 22088 12038 22140 12044
rect 22100 11558 22128 12038
rect 22088 11552 22140 11558
rect 22088 11494 22140 11500
rect 22100 11150 22128 11494
rect 21996 11144 22048 11150
rect 21996 11086 22048 11092
rect 22088 11144 22140 11150
rect 22088 11086 22140 11092
rect 21904 10804 21956 10810
rect 21904 10746 21956 10752
rect 21916 10538 21944 10746
rect 21904 10532 21956 10538
rect 21904 10474 21956 10480
rect 22100 10146 22128 11086
rect 22192 10606 22220 13126
rect 22744 12481 22772 14758
rect 23100 14476 23152 14482
rect 23100 14418 23152 14424
rect 23112 13870 23140 14418
rect 23100 13864 23152 13870
rect 23100 13806 23152 13812
rect 23190 13832 23246 13841
rect 23190 13767 23246 13776
rect 23204 13530 23232 13767
rect 23296 13530 23324 21814
rect 23572 21706 23600 27095
rect 24478 25392 24534 25401
rect 24478 25327 24534 25336
rect 24001 25052 24297 25072
rect 24057 25050 24081 25052
rect 24137 25050 24161 25052
rect 24217 25050 24241 25052
rect 24079 24998 24081 25050
rect 24143 24998 24155 25050
rect 24217 24998 24219 25050
rect 24057 24996 24081 24998
rect 24137 24996 24161 24998
rect 24217 24996 24241 24998
rect 24001 24976 24297 24996
rect 24386 24304 24442 24313
rect 24386 24239 24442 24248
rect 24001 23964 24297 23984
rect 24057 23962 24081 23964
rect 24137 23962 24161 23964
rect 24217 23962 24241 23964
rect 24079 23910 24081 23962
rect 24143 23910 24155 23962
rect 24217 23910 24219 23962
rect 24057 23908 24081 23910
rect 24137 23908 24161 23910
rect 24217 23908 24241 23910
rect 24001 23888 24297 23908
rect 23742 23760 23798 23769
rect 23742 23695 23798 23704
rect 23652 23656 23704 23662
rect 23652 23598 23704 23604
rect 23664 22642 23692 23598
rect 23652 22636 23704 22642
rect 23652 22578 23704 22584
rect 23756 21962 23784 23695
rect 23836 23180 23888 23186
rect 23836 23122 23888 23128
rect 23848 22438 23876 23122
rect 24001 22876 24297 22896
rect 24057 22874 24081 22876
rect 24137 22874 24161 22876
rect 24217 22874 24241 22876
rect 24079 22822 24081 22874
rect 24143 22822 24155 22874
rect 24217 22822 24219 22874
rect 24057 22820 24081 22822
rect 24137 22820 24161 22822
rect 24217 22820 24241 22822
rect 24001 22800 24297 22820
rect 24400 22794 24428 24239
rect 24492 23866 24520 25327
rect 24860 24410 24888 27520
rect 25122 26072 25178 26081
rect 25122 26007 25178 26016
rect 24848 24404 24900 24410
rect 24848 24346 24900 24352
rect 24480 23860 24532 23866
rect 24480 23802 24532 23808
rect 24480 23316 24532 23322
rect 24480 23258 24532 23264
rect 24492 23225 24520 23258
rect 24478 23216 24534 23225
rect 24478 23151 24534 23160
rect 24400 22778 24612 22794
rect 24400 22772 24624 22778
rect 24400 22766 24572 22772
rect 24572 22714 24624 22720
rect 24478 22672 24534 22681
rect 24478 22607 24534 22616
rect 23836 22432 23888 22438
rect 24388 22432 24440 22438
rect 23836 22374 23888 22380
rect 24386 22400 24388 22409
rect 24440 22400 24442 22409
rect 24386 22335 24442 22344
rect 24388 22092 24440 22098
rect 24388 22034 24440 22040
rect 23744 21956 23796 21962
rect 23744 21898 23796 21904
rect 24001 21788 24297 21808
rect 24057 21786 24081 21788
rect 24137 21786 24161 21788
rect 24217 21786 24241 21788
rect 24079 21734 24081 21786
rect 24143 21734 24155 21786
rect 24217 21734 24219 21786
rect 24057 21732 24081 21734
rect 24137 21732 24161 21734
rect 24217 21732 24241 21734
rect 24001 21712 24297 21732
rect 23480 21678 23600 21706
rect 23376 20392 23428 20398
rect 23376 20334 23428 20340
rect 23388 19990 23416 20334
rect 23376 19984 23428 19990
rect 23376 19926 23428 19932
rect 23480 14074 23508 21678
rect 23558 21584 23614 21593
rect 24400 21554 24428 22034
rect 24492 21690 24520 22607
rect 24664 22568 24716 22574
rect 24664 22510 24716 22516
rect 24754 22536 24810 22545
rect 24676 22001 24704 22510
rect 24754 22471 24810 22480
rect 24662 21992 24718 22001
rect 24662 21927 24718 21936
rect 24480 21684 24532 21690
rect 24480 21626 24532 21632
rect 23558 21519 23614 21528
rect 24388 21548 24440 21554
rect 23572 20602 23600 21519
rect 24388 21490 24440 21496
rect 24112 21480 24164 21486
rect 24110 21448 24112 21457
rect 24296 21480 24348 21486
rect 24164 21448 24166 21457
rect 24296 21422 24348 21428
rect 24386 21448 24442 21457
rect 24110 21383 24166 21392
rect 24308 21078 24336 21422
rect 24386 21383 24442 21392
rect 24296 21072 24348 21078
rect 24296 21014 24348 21020
rect 24001 20700 24297 20720
rect 24057 20698 24081 20700
rect 24137 20698 24161 20700
rect 24217 20698 24241 20700
rect 24079 20646 24081 20698
rect 24143 20646 24155 20698
rect 24217 20646 24219 20698
rect 24057 20644 24081 20646
rect 24137 20644 24161 20646
rect 24217 20644 24241 20646
rect 24001 20624 24297 20644
rect 23560 20596 23612 20602
rect 23560 20538 23612 20544
rect 24400 20058 24428 21383
rect 24768 21146 24796 22471
rect 24756 21140 24808 21146
rect 24756 21082 24808 21088
rect 24572 21004 24624 21010
rect 24572 20946 24624 20952
rect 24478 20904 24534 20913
rect 24478 20839 24534 20848
rect 24388 20052 24440 20058
rect 24388 19994 24440 20000
rect 24388 19916 24440 19922
rect 24388 19858 24440 19864
rect 24001 19612 24297 19632
rect 24057 19610 24081 19612
rect 24137 19610 24161 19612
rect 24217 19610 24241 19612
rect 24079 19558 24081 19610
rect 24143 19558 24155 19610
rect 24217 19558 24219 19610
rect 24057 19556 24081 19558
rect 24137 19556 24161 19558
rect 24217 19556 24241 19558
rect 24001 19536 24297 19556
rect 23834 19408 23890 19417
rect 23890 19366 23968 19394
rect 23834 19343 23890 19352
rect 23652 19304 23704 19310
rect 23652 19246 23704 19252
rect 23664 18290 23692 19246
rect 23834 19136 23890 19145
rect 23834 19071 23890 19080
rect 23652 18284 23704 18290
rect 23652 18226 23704 18232
rect 23848 17649 23876 19071
rect 23834 17640 23890 17649
rect 23834 17575 23890 17584
rect 23834 17232 23890 17241
rect 23834 17167 23890 17176
rect 23848 16250 23876 17167
rect 23836 16244 23888 16250
rect 23836 16186 23888 16192
rect 23836 16040 23888 16046
rect 23836 15982 23888 15988
rect 23742 15056 23798 15065
rect 23848 15026 23876 15982
rect 23742 14991 23798 15000
rect 23836 15020 23888 15026
rect 23560 14952 23612 14958
rect 23560 14894 23612 14900
rect 23468 14068 23520 14074
rect 23468 14010 23520 14016
rect 23192 13524 23244 13530
rect 23192 13466 23244 13472
rect 23284 13524 23336 13530
rect 23284 13466 23336 13472
rect 22916 13388 22968 13394
rect 22916 13330 22968 13336
rect 22928 12986 22956 13330
rect 23100 13320 23152 13326
rect 23100 13262 23152 13268
rect 22916 12980 22968 12986
rect 22916 12922 22968 12928
rect 22730 12472 22786 12481
rect 22640 12436 22692 12442
rect 22730 12407 22786 12416
rect 22640 12378 22692 12384
rect 22364 11552 22416 11558
rect 22364 11494 22416 11500
rect 22376 11121 22404 11494
rect 22652 11286 22680 12378
rect 22822 12336 22878 12345
rect 22822 12271 22878 12280
rect 22836 11898 22864 12271
rect 22824 11892 22876 11898
rect 22824 11834 22876 11840
rect 22836 11694 22864 11834
rect 22824 11688 22876 11694
rect 22824 11630 22876 11636
rect 22928 11626 22956 12922
rect 23006 12472 23062 12481
rect 23112 12442 23140 13262
rect 23204 12986 23232 13466
rect 23376 13184 23428 13190
rect 23376 13126 23428 13132
rect 23192 12980 23244 12986
rect 23192 12922 23244 12928
rect 23388 12782 23416 13126
rect 23376 12776 23428 12782
rect 23374 12744 23376 12753
rect 23428 12744 23430 12753
rect 23374 12679 23430 12688
rect 23006 12407 23062 12416
rect 23100 12436 23152 12442
rect 22916 11620 22968 11626
rect 22916 11562 22968 11568
rect 22640 11280 22692 11286
rect 22640 11222 22692 11228
rect 22362 11112 22418 11121
rect 22362 11047 22418 11056
rect 22272 11008 22324 11014
rect 22272 10950 22324 10956
rect 22284 10674 22312 10950
rect 22652 10810 22680 11222
rect 22822 11112 22878 11121
rect 22822 11047 22878 11056
rect 22640 10804 22692 10810
rect 22640 10746 22692 10752
rect 22272 10668 22324 10674
rect 22272 10610 22324 10616
rect 22180 10600 22232 10606
rect 22180 10542 22232 10548
rect 22192 10266 22220 10542
rect 22180 10260 22232 10266
rect 22180 10202 22232 10208
rect 22100 10118 22312 10146
rect 22284 9926 22312 10118
rect 22272 9920 22324 9926
rect 22272 9862 22324 9868
rect 21812 9172 21864 9178
rect 21812 9114 21864 9120
rect 21824 8888 21852 9114
rect 22284 8906 22312 9862
rect 22836 9654 22864 11047
rect 22824 9648 22876 9654
rect 22824 9590 22876 9596
rect 22364 9376 22416 9382
rect 22364 9318 22416 9324
rect 22272 8900 22324 8906
rect 21824 8860 21944 8888
rect 21732 8758 21852 8786
rect 21628 8016 21680 8022
rect 21628 7958 21680 7964
rect 21352 7948 21404 7954
rect 21352 7890 21404 7896
rect 21364 7546 21392 7890
rect 21260 7540 21312 7546
rect 21260 7482 21312 7488
rect 21352 7540 21404 7546
rect 21352 7482 21404 7488
rect 21444 7404 21496 7410
rect 21444 7346 21496 7352
rect 21260 7200 21312 7206
rect 21260 7142 21312 7148
rect 21272 7002 21300 7142
rect 21260 6996 21312 7002
rect 21260 6938 21312 6944
rect 20984 6860 21036 6866
rect 20984 6802 21036 6808
rect 20892 6792 20944 6798
rect 20892 6734 20944 6740
rect 20340 6724 20392 6730
rect 20340 6666 20392 6672
rect 20352 6458 20380 6666
rect 20904 6497 20932 6734
rect 20890 6488 20946 6497
rect 20340 6452 20392 6458
rect 20890 6423 20892 6432
rect 20340 6394 20392 6400
rect 20944 6423 20946 6432
rect 20892 6394 20944 6400
rect 20352 5846 20380 6394
rect 20340 5840 20392 5846
rect 20340 5782 20392 5788
rect 20352 5370 20380 5782
rect 20616 5704 20668 5710
rect 20616 5646 20668 5652
rect 20340 5364 20392 5370
rect 20340 5306 20392 5312
rect 20248 5228 20300 5234
rect 20248 5170 20300 5176
rect 20154 4448 20210 4457
rect 20154 4383 20210 4392
rect 19878 4176 19934 4185
rect 19878 4111 19934 4120
rect 19788 3936 19840 3942
rect 19788 3878 19840 3884
rect 19972 3936 20024 3942
rect 20064 3936 20116 3942
rect 19972 3878 20024 3884
rect 20062 3904 20064 3913
rect 20116 3904 20118 3913
rect 19334 3836 19630 3856
rect 19390 3834 19414 3836
rect 19470 3834 19494 3836
rect 19550 3834 19574 3836
rect 19412 3782 19414 3834
rect 19476 3782 19488 3834
rect 19550 3782 19552 3834
rect 19390 3780 19414 3782
rect 19470 3780 19494 3782
rect 19550 3780 19574 3782
rect 19334 3760 19630 3780
rect 19694 3632 19750 3641
rect 19694 3567 19750 3576
rect 19234 3224 19290 3233
rect 19234 3159 19290 3168
rect 19142 2816 19198 2825
rect 19142 2751 19198 2760
rect 19334 2748 19630 2768
rect 19390 2746 19414 2748
rect 19470 2746 19494 2748
rect 19550 2746 19574 2748
rect 19412 2694 19414 2746
rect 19476 2694 19488 2746
rect 19550 2694 19552 2746
rect 19390 2692 19414 2694
rect 19470 2692 19494 2694
rect 19550 2692 19574 2694
rect 19334 2672 19630 2692
rect 19052 2644 19104 2650
rect 19052 2586 19104 2592
rect 19708 2530 19736 3567
rect 19984 3398 20012 3878
rect 20062 3839 20118 3848
rect 19972 3392 20024 3398
rect 19970 3360 19972 3369
rect 20024 3360 20026 3369
rect 19970 3295 20026 3304
rect 20260 3074 20288 5170
rect 20352 4826 20380 5306
rect 20628 5234 20656 5646
rect 20616 5228 20668 5234
rect 20616 5170 20668 5176
rect 20340 4820 20392 4826
rect 20340 4762 20392 4768
rect 20352 4214 20380 4762
rect 20616 4616 20668 4622
rect 20616 4558 20668 4564
rect 20340 4208 20392 4214
rect 20340 4150 20392 4156
rect 20628 4049 20656 4558
rect 20708 4140 20760 4146
rect 20708 4082 20760 4088
rect 20614 4040 20670 4049
rect 20614 3975 20670 3984
rect 20720 3097 20748 4082
rect 20904 4078 20932 6394
rect 20996 5574 21024 6802
rect 21456 5914 21484 7346
rect 21536 7200 21588 7206
rect 21534 7168 21536 7177
rect 21588 7168 21590 7177
rect 21534 7103 21590 7112
rect 21824 7018 21852 8758
rect 21916 8430 21944 8860
rect 22272 8842 22324 8848
rect 22180 8832 22232 8838
rect 22180 8774 22232 8780
rect 22192 8498 22220 8774
rect 22180 8492 22232 8498
rect 22180 8434 22232 8440
rect 21904 8424 21956 8430
rect 21904 8366 21956 8372
rect 21996 7744 22048 7750
rect 21996 7686 22048 7692
rect 22180 7744 22232 7750
rect 22180 7686 22232 7692
rect 22008 7449 22036 7686
rect 21994 7440 22050 7449
rect 21994 7375 22050 7384
rect 22192 7206 22220 7686
rect 22180 7200 22232 7206
rect 22180 7142 22232 7148
rect 21824 6990 21944 7018
rect 21812 6928 21864 6934
rect 21626 6896 21682 6905
rect 21812 6870 21864 6876
rect 21626 6831 21682 6840
rect 21534 6624 21590 6633
rect 21534 6559 21590 6568
rect 21548 6458 21576 6559
rect 21536 6452 21588 6458
rect 21536 6394 21588 6400
rect 21548 6118 21576 6394
rect 21536 6112 21588 6118
rect 21536 6054 21588 6060
rect 21444 5908 21496 5914
rect 21444 5850 21496 5856
rect 20984 5568 21036 5574
rect 20984 5510 21036 5516
rect 21456 5166 21484 5850
rect 21536 5568 21588 5574
rect 21536 5510 21588 5516
rect 21444 5160 21496 5166
rect 21444 5102 21496 5108
rect 21548 4486 21576 5510
rect 21536 4480 21588 4486
rect 21536 4422 21588 4428
rect 21442 4176 21498 4185
rect 21442 4111 21498 4120
rect 20892 4072 20944 4078
rect 20892 4014 20944 4020
rect 21168 3936 21220 3942
rect 21168 3878 21220 3884
rect 21180 3738 21208 3878
rect 21168 3732 21220 3738
rect 21168 3674 21220 3680
rect 21260 3528 21312 3534
rect 20890 3496 20946 3505
rect 21260 3470 21312 3476
rect 21352 3528 21404 3534
rect 21352 3470 21404 3476
rect 20890 3431 20946 3440
rect 20800 3392 20852 3398
rect 20800 3334 20852 3340
rect 20706 3088 20762 3097
rect 20260 3058 20472 3074
rect 20248 3052 20472 3058
rect 20300 3046 20472 3052
rect 20248 2994 20300 3000
rect 20248 2916 20300 2922
rect 20248 2858 20300 2864
rect 19524 2502 19736 2530
rect 19524 480 19552 2502
rect 20260 2310 20288 2858
rect 20444 2514 20472 3046
rect 20706 3023 20762 3032
rect 20720 2650 20748 3023
rect 20812 2689 20840 3334
rect 20798 2680 20854 2689
rect 20708 2644 20760 2650
rect 20798 2615 20854 2624
rect 20708 2586 20760 2592
rect 20904 2530 20932 3431
rect 21272 3194 21300 3470
rect 21260 3188 21312 3194
rect 21260 3130 21312 3136
rect 21364 2990 21392 3470
rect 21352 2984 21404 2990
rect 21352 2926 21404 2932
rect 21364 2650 21392 2926
rect 21352 2644 21404 2650
rect 21352 2586 21404 2592
rect 20432 2508 20484 2514
rect 20432 2450 20484 2456
rect 20812 2502 20932 2530
rect 20248 2304 20300 2310
rect 20248 2246 20300 2252
rect 20154 1864 20210 1873
rect 20154 1799 20210 1808
rect 20168 480 20196 1799
rect 20260 1601 20288 2246
rect 20246 1592 20302 1601
rect 20246 1527 20302 1536
rect 20812 480 20840 2502
rect 21456 480 21484 4111
rect 21548 3942 21576 4422
rect 21536 3936 21588 3942
rect 21536 3878 21588 3884
rect 21548 3777 21576 3878
rect 21534 3768 21590 3777
rect 21534 3703 21590 3712
rect 21640 2038 21668 6831
rect 21824 6662 21852 6870
rect 21916 6866 21944 6990
rect 21904 6860 21956 6866
rect 21904 6802 21956 6808
rect 22088 6792 22140 6798
rect 22088 6734 22140 6740
rect 21812 6656 21864 6662
rect 21812 6598 21864 6604
rect 21718 6488 21774 6497
rect 21718 6423 21720 6432
rect 21772 6423 21774 6432
rect 21720 6394 21772 6400
rect 21824 6186 21852 6598
rect 21812 6180 21864 6186
rect 21812 6122 21864 6128
rect 22100 5778 22128 6734
rect 22180 6656 22232 6662
rect 22180 6598 22232 6604
rect 22192 6322 22220 6598
rect 22376 6361 22404 9318
rect 22456 8356 22508 8362
rect 22456 8298 22508 8304
rect 22468 7546 22496 8298
rect 22916 7744 22968 7750
rect 22916 7686 22968 7692
rect 22456 7540 22508 7546
rect 22456 7482 22508 7488
rect 22928 7342 22956 7686
rect 22916 7336 22968 7342
rect 22916 7278 22968 7284
rect 22548 6860 22600 6866
rect 22548 6802 22600 6808
rect 22560 6458 22588 6802
rect 22548 6452 22600 6458
rect 22468 6412 22548 6440
rect 22362 6352 22418 6361
rect 22180 6316 22232 6322
rect 22362 6287 22418 6296
rect 22180 6258 22232 6264
rect 22272 6180 22324 6186
rect 22272 6122 22324 6128
rect 22180 6112 22232 6118
rect 22180 6054 22232 6060
rect 22192 5953 22220 6054
rect 22178 5944 22234 5953
rect 22178 5879 22234 5888
rect 22088 5772 22140 5778
rect 22088 5714 22140 5720
rect 22086 4856 22142 4865
rect 22086 4791 22088 4800
rect 22140 4791 22142 4800
rect 22088 4762 22140 4768
rect 21994 4720 22050 4729
rect 21994 4655 21996 4664
rect 22048 4655 22050 4664
rect 21996 4626 22048 4632
rect 22008 4282 22036 4626
rect 21996 4276 22048 4282
rect 21996 4218 22048 4224
rect 21720 4004 21772 4010
rect 21720 3946 21772 3952
rect 21732 2938 21760 3946
rect 22100 3738 22128 4762
rect 22284 4758 22312 6122
rect 22468 5370 22496 6412
rect 22548 6394 22600 6400
rect 22548 5704 22600 5710
rect 22546 5672 22548 5681
rect 22600 5672 22602 5681
rect 22546 5607 22602 5616
rect 22916 5568 22968 5574
rect 22916 5510 22968 5516
rect 22456 5364 22508 5370
rect 22456 5306 22508 5312
rect 22730 5264 22786 5273
rect 22730 5199 22786 5208
rect 22272 4752 22324 4758
rect 22272 4694 22324 4700
rect 22272 4616 22324 4622
rect 22272 4558 22324 4564
rect 22284 4214 22312 4558
rect 22640 4480 22692 4486
rect 22640 4422 22692 4428
rect 22272 4208 22324 4214
rect 22272 4150 22324 4156
rect 22088 3732 22140 3738
rect 22088 3674 22140 3680
rect 22652 3602 22680 4422
rect 22640 3596 22692 3602
rect 22640 3538 22692 3544
rect 21732 2910 21852 2938
rect 21720 2848 21772 2854
rect 21720 2790 21772 2796
rect 21732 2553 21760 2790
rect 21718 2544 21774 2553
rect 21824 2530 21852 2910
rect 21902 2544 21958 2553
rect 21824 2502 21902 2530
rect 21718 2479 21720 2488
rect 21772 2479 21774 2488
rect 21902 2479 21958 2488
rect 21720 2450 21772 2456
rect 21732 2419 21760 2450
rect 21628 2032 21680 2038
rect 21628 1974 21680 1980
rect 22088 604 22140 610
rect 22088 546 22140 552
rect 22100 480 22128 546
rect 22744 480 22772 5199
rect 22928 4486 22956 5510
rect 22916 4480 22968 4486
rect 22916 4422 22968 4428
rect 23020 2650 23048 12407
rect 23100 12378 23152 12384
rect 23192 11552 23244 11558
rect 23192 11494 23244 11500
rect 23376 11552 23428 11558
rect 23376 11494 23428 11500
rect 23204 11098 23232 11494
rect 23112 11070 23232 11098
rect 23112 7993 23140 11070
rect 23284 10600 23336 10606
rect 23284 10542 23336 10548
rect 23296 10062 23324 10542
rect 23388 10266 23416 11494
rect 23376 10260 23428 10266
rect 23376 10202 23428 10208
rect 23284 10056 23336 10062
rect 23284 9998 23336 10004
rect 23388 9654 23416 10202
rect 23376 9648 23428 9654
rect 23190 9616 23246 9625
rect 23376 9590 23428 9596
rect 23190 9551 23192 9560
rect 23244 9551 23246 9560
rect 23192 9522 23244 9528
rect 23468 9376 23520 9382
rect 23468 9318 23520 9324
rect 23192 9104 23244 9110
rect 23192 9046 23244 9052
rect 23204 8566 23232 9046
rect 23376 8832 23428 8838
rect 23480 8809 23508 9318
rect 23376 8774 23428 8780
rect 23466 8800 23522 8809
rect 23192 8560 23244 8566
rect 23192 8502 23244 8508
rect 23388 8430 23416 8774
rect 23466 8735 23522 8744
rect 23192 8424 23244 8430
rect 23192 8366 23244 8372
rect 23376 8424 23428 8430
rect 23376 8366 23428 8372
rect 23204 8090 23232 8366
rect 23192 8084 23244 8090
rect 23192 8026 23244 8032
rect 23098 7984 23154 7993
rect 23098 7919 23100 7928
rect 23152 7919 23154 7928
rect 23100 7890 23152 7896
rect 23112 7478 23140 7890
rect 23100 7472 23152 7478
rect 23100 7414 23152 7420
rect 23468 7200 23520 7206
rect 23468 7142 23520 7148
rect 23376 6724 23428 6730
rect 23376 6666 23428 6672
rect 23284 6248 23336 6254
rect 23284 6190 23336 6196
rect 23100 6112 23152 6118
rect 23100 6054 23152 6060
rect 23112 4214 23140 6054
rect 23296 5710 23324 6190
rect 23388 5914 23416 6666
rect 23376 5908 23428 5914
rect 23376 5850 23428 5856
rect 23374 5808 23430 5817
rect 23374 5743 23430 5752
rect 23284 5704 23336 5710
rect 23284 5646 23336 5652
rect 23282 5400 23338 5409
rect 23282 5335 23338 5344
rect 23192 5092 23244 5098
rect 23192 5034 23244 5040
rect 23204 4826 23232 5034
rect 23192 4820 23244 4826
rect 23192 4762 23244 4768
rect 23192 4480 23244 4486
rect 23192 4422 23244 4428
rect 23204 4321 23232 4422
rect 23190 4312 23246 4321
rect 23190 4247 23246 4256
rect 23100 4208 23152 4214
rect 23100 4150 23152 4156
rect 23296 4146 23324 5335
rect 23388 4826 23416 5743
rect 23480 5234 23508 7142
rect 23572 5370 23600 14894
rect 23652 13728 23704 13734
rect 23652 13670 23704 13676
rect 23664 12850 23692 13670
rect 23756 13025 23784 14991
rect 23836 14962 23888 14968
rect 23742 13016 23798 13025
rect 23940 13002 23968 19366
rect 24400 19174 24428 19858
rect 24492 19174 24520 20839
rect 24584 20262 24612 20946
rect 24572 20256 24624 20262
rect 24570 20224 24572 20233
rect 24624 20224 24626 20233
rect 24570 20159 24626 20168
rect 24846 19680 24902 19689
rect 24846 19615 24902 19624
rect 24112 19168 24164 19174
rect 24112 19110 24164 19116
rect 24388 19168 24440 19174
rect 24388 19110 24440 19116
rect 24480 19168 24532 19174
rect 24480 19110 24532 19116
rect 24124 18873 24152 19110
rect 24110 18864 24166 18873
rect 24110 18799 24166 18808
rect 24386 18592 24442 18601
rect 24001 18524 24297 18544
rect 24386 18527 24442 18536
rect 24057 18522 24081 18524
rect 24137 18522 24161 18524
rect 24217 18522 24241 18524
rect 24079 18470 24081 18522
rect 24143 18470 24155 18522
rect 24217 18470 24219 18522
rect 24057 18468 24081 18470
rect 24137 18468 24161 18470
rect 24217 18468 24241 18470
rect 24001 18448 24297 18468
rect 24001 17436 24297 17456
rect 24057 17434 24081 17436
rect 24137 17434 24161 17436
rect 24217 17434 24241 17436
rect 24079 17382 24081 17434
rect 24143 17382 24155 17434
rect 24217 17382 24219 17434
rect 24057 17380 24081 17382
rect 24137 17380 24161 17382
rect 24217 17380 24241 17382
rect 24001 17360 24297 17380
rect 24400 17338 24428 18527
rect 24860 18426 24888 19615
rect 24848 18420 24900 18426
rect 24848 18362 24900 18368
rect 24664 18216 24716 18222
rect 24664 18158 24716 18164
rect 24478 18048 24534 18057
rect 24478 17983 24534 17992
rect 24388 17332 24440 17338
rect 24388 17274 24440 17280
rect 24296 17128 24348 17134
rect 24296 17070 24348 17076
rect 24308 16697 24336 17070
rect 24492 16794 24520 17983
rect 24676 17105 24704 18158
rect 24662 17096 24718 17105
rect 24662 17031 24718 17040
rect 24480 16788 24532 16794
rect 24480 16730 24532 16736
rect 24294 16688 24350 16697
rect 24478 16688 24534 16697
rect 24294 16623 24350 16632
rect 24388 16652 24440 16658
rect 24478 16623 24534 16632
rect 24388 16594 24440 16600
rect 24001 16348 24297 16368
rect 24057 16346 24081 16348
rect 24137 16346 24161 16348
rect 24217 16346 24241 16348
rect 24079 16294 24081 16346
rect 24143 16294 24155 16346
rect 24217 16294 24219 16346
rect 24057 16292 24081 16294
rect 24137 16292 24161 16294
rect 24217 16292 24241 16294
rect 24001 16272 24297 16292
rect 24400 15910 24428 16594
rect 24112 15904 24164 15910
rect 24112 15846 24164 15852
rect 24388 15904 24440 15910
rect 24388 15846 24440 15852
rect 24124 15638 24152 15846
rect 24386 15736 24442 15745
rect 24386 15671 24442 15680
rect 24112 15632 24164 15638
rect 24112 15574 24164 15580
rect 24400 15570 24428 15671
rect 24388 15564 24440 15570
rect 24388 15506 24440 15512
rect 24001 15260 24297 15280
rect 24057 15258 24081 15260
rect 24137 15258 24161 15260
rect 24217 15258 24241 15260
rect 24079 15206 24081 15258
rect 24143 15206 24155 15258
rect 24217 15206 24219 15258
rect 24057 15204 24081 15206
rect 24137 15204 24161 15206
rect 24217 15204 24241 15206
rect 24001 15184 24297 15204
rect 24400 15162 24428 15506
rect 24492 15178 24520 16623
rect 24662 16280 24718 16289
rect 24662 16215 24718 16224
rect 24492 15162 24612 15178
rect 24388 15156 24440 15162
rect 24492 15156 24624 15162
rect 24492 15150 24572 15156
rect 24388 15098 24440 15104
rect 24572 15098 24624 15104
rect 24676 14618 24704 16215
rect 24848 14952 24900 14958
rect 24848 14894 24900 14900
rect 24664 14612 24716 14618
rect 24664 14554 24716 14560
rect 24860 14550 24888 14894
rect 24848 14544 24900 14550
rect 24848 14486 24900 14492
rect 24388 14476 24440 14482
rect 24388 14418 24440 14424
rect 24001 14172 24297 14192
rect 24057 14170 24081 14172
rect 24137 14170 24161 14172
rect 24217 14170 24241 14172
rect 24079 14118 24081 14170
rect 24143 14118 24155 14170
rect 24217 14118 24219 14170
rect 24057 14116 24081 14118
rect 24137 14116 24161 14118
rect 24217 14116 24241 14118
rect 24001 14096 24297 14116
rect 24400 13977 24428 14418
rect 24848 14000 24900 14006
rect 24386 13968 24442 13977
rect 24386 13903 24442 13912
rect 24846 13968 24848 13977
rect 24900 13968 24902 13977
rect 24846 13903 24902 13912
rect 24388 13388 24440 13394
rect 24388 13330 24440 13336
rect 24001 13084 24297 13104
rect 24057 13082 24081 13084
rect 24137 13082 24161 13084
rect 24217 13082 24241 13084
rect 24079 13030 24081 13082
rect 24143 13030 24155 13082
rect 24217 13030 24219 13082
rect 24057 13028 24081 13030
rect 24137 13028 24161 13030
rect 24217 13028 24241 13030
rect 24001 13008 24297 13028
rect 23742 12951 23798 12960
rect 23848 12974 23968 13002
rect 23652 12844 23704 12850
rect 23652 12786 23704 12792
rect 23848 12458 23876 12974
rect 24296 12912 24348 12918
rect 24294 12880 24296 12889
rect 24348 12880 24350 12889
rect 24400 12866 24428 13330
rect 24846 13288 24902 13297
rect 24846 13223 24902 13232
rect 24860 12986 24888 13223
rect 24848 12980 24900 12986
rect 24848 12922 24900 12928
rect 24350 12838 24428 12866
rect 24478 12880 24534 12889
rect 24294 12815 24350 12824
rect 24478 12815 24534 12824
rect 23756 12430 23876 12458
rect 23756 10826 23784 12430
rect 24001 11996 24297 12016
rect 24057 11994 24081 11996
rect 24137 11994 24161 11996
rect 24217 11994 24241 11996
rect 24079 11942 24081 11994
rect 24143 11942 24155 11994
rect 24217 11942 24219 11994
rect 24057 11940 24081 11942
rect 24137 11940 24161 11942
rect 24217 11940 24241 11942
rect 24001 11920 24297 11940
rect 24492 11898 24520 12815
rect 24756 12300 24808 12306
rect 24756 12242 24808 12248
rect 24768 11898 24796 12242
rect 25136 11898 25164 26007
rect 25950 22400 26006 22409
rect 25950 22335 26006 22344
rect 25306 14648 25362 14657
rect 25306 14583 25362 14592
rect 25320 12986 25348 14583
rect 25398 13424 25454 13433
rect 25398 13359 25454 13368
rect 25308 12980 25360 12986
rect 25308 12922 25360 12928
rect 25320 12782 25348 12922
rect 25308 12776 25360 12782
rect 25308 12718 25360 12724
rect 24480 11892 24532 11898
rect 24480 11834 24532 11840
rect 24756 11892 24808 11898
rect 24756 11834 24808 11840
rect 25124 11892 25176 11898
rect 25124 11834 25176 11840
rect 24478 11792 24534 11801
rect 23928 11756 23980 11762
rect 24478 11727 24534 11736
rect 23928 11698 23980 11704
rect 23940 11014 23968 11698
rect 23928 11008 23980 11014
rect 23928 10950 23980 10956
rect 24001 10908 24297 10928
rect 24057 10906 24081 10908
rect 24137 10906 24161 10908
rect 24217 10906 24241 10908
rect 24079 10854 24081 10906
rect 24143 10854 24155 10906
rect 24217 10854 24219 10906
rect 24057 10852 24081 10854
rect 24137 10852 24161 10854
rect 24217 10852 24241 10854
rect 24001 10832 24297 10852
rect 23756 10798 23968 10826
rect 23834 10568 23890 10577
rect 23834 10503 23890 10512
rect 23744 9580 23796 9586
rect 23744 9522 23796 9528
rect 23756 9450 23784 9522
rect 23744 9444 23796 9450
rect 23744 9386 23796 9392
rect 23744 8832 23796 8838
rect 23744 8774 23796 8780
rect 23756 8362 23784 8774
rect 23744 8356 23796 8362
rect 23744 8298 23796 8304
rect 23650 8256 23706 8265
rect 23650 8191 23706 8200
rect 23664 8090 23692 8191
rect 23652 8084 23704 8090
rect 23652 8026 23704 8032
rect 23664 7546 23692 8026
rect 23756 7886 23784 8298
rect 23744 7880 23796 7886
rect 23744 7822 23796 7828
rect 23652 7540 23704 7546
rect 23652 7482 23704 7488
rect 23848 7290 23876 10503
rect 23940 7886 23968 10798
rect 24386 10024 24442 10033
rect 24492 10010 24520 11727
rect 24940 11688 24992 11694
rect 24940 11630 24992 11636
rect 24952 11257 24980 11630
rect 24938 11248 24994 11257
rect 25412 11218 25440 13359
rect 24938 11183 24994 11192
rect 25400 11212 25452 11218
rect 25400 11154 25452 11160
rect 24940 11076 24992 11082
rect 24940 11018 24992 11024
rect 24756 11008 24808 11014
rect 24756 10950 24808 10956
rect 24768 10470 24796 10950
rect 24756 10464 24808 10470
rect 24756 10406 24808 10412
rect 24768 10198 24796 10406
rect 24756 10192 24808 10198
rect 24952 10169 24980 11018
rect 25412 10810 25440 11154
rect 25400 10804 25452 10810
rect 25400 10746 25452 10752
rect 24756 10134 24808 10140
rect 24938 10160 24994 10169
rect 24492 9982 24612 10010
rect 24386 9959 24442 9968
rect 24001 9820 24297 9840
rect 24057 9818 24081 9820
rect 24137 9818 24161 9820
rect 24217 9818 24241 9820
rect 24079 9766 24081 9818
rect 24143 9766 24155 9818
rect 24217 9766 24219 9818
rect 24057 9764 24081 9766
rect 24137 9764 24161 9766
rect 24217 9764 24241 9766
rect 24001 9744 24297 9764
rect 24020 9580 24072 9586
rect 24020 9522 24072 9528
rect 24032 9110 24060 9522
rect 24020 9104 24072 9110
rect 24020 9046 24072 9052
rect 24001 8732 24297 8752
rect 24057 8730 24081 8732
rect 24137 8730 24161 8732
rect 24217 8730 24241 8732
rect 24079 8678 24081 8730
rect 24143 8678 24155 8730
rect 24217 8678 24219 8730
rect 24057 8676 24081 8678
rect 24137 8676 24161 8678
rect 24217 8676 24241 8678
rect 24001 8656 24297 8676
rect 23928 7880 23980 7886
rect 23928 7822 23980 7828
rect 23928 7744 23980 7750
rect 23928 7686 23980 7692
rect 23756 7262 23876 7290
rect 23652 6656 23704 6662
rect 23652 6598 23704 6604
rect 23664 6186 23692 6598
rect 23652 6180 23704 6186
rect 23652 6122 23704 6128
rect 23652 5840 23704 5846
rect 23652 5782 23704 5788
rect 23560 5364 23612 5370
rect 23560 5306 23612 5312
rect 23468 5228 23520 5234
rect 23468 5170 23520 5176
rect 23560 5160 23612 5166
rect 23560 5102 23612 5108
rect 23376 4820 23428 4826
rect 23376 4762 23428 4768
rect 23388 4282 23416 4762
rect 23376 4276 23428 4282
rect 23376 4218 23428 4224
rect 23284 4140 23336 4146
rect 23284 4082 23336 4088
rect 23190 3904 23246 3913
rect 23190 3839 23246 3848
rect 23204 3194 23232 3839
rect 23572 3670 23600 5102
rect 23664 5030 23692 5782
rect 23652 5024 23704 5030
rect 23756 5001 23784 7262
rect 23940 7206 23968 7686
rect 24001 7644 24297 7664
rect 24057 7642 24081 7644
rect 24137 7642 24161 7644
rect 24217 7642 24241 7644
rect 24079 7590 24081 7642
rect 24143 7590 24155 7642
rect 24217 7590 24219 7642
rect 24057 7588 24081 7590
rect 24137 7588 24161 7590
rect 24217 7588 24241 7590
rect 24001 7568 24297 7588
rect 24020 7404 24072 7410
rect 24020 7346 24072 7352
rect 23836 7200 23888 7206
rect 23836 7142 23888 7148
rect 23928 7200 23980 7206
rect 23928 7142 23980 7148
rect 23848 7002 23876 7142
rect 23836 6996 23888 7002
rect 23836 6938 23888 6944
rect 23848 6497 23876 6938
rect 23834 6488 23890 6497
rect 23834 6423 23890 6432
rect 23834 5944 23890 5953
rect 23834 5879 23890 5888
rect 23652 4966 23704 4972
rect 23742 4992 23798 5001
rect 23664 4842 23692 4966
rect 23742 4927 23798 4936
rect 23664 4814 23784 4842
rect 23756 4622 23784 4814
rect 23744 4616 23796 4622
rect 23744 4558 23796 4564
rect 23756 3738 23784 4558
rect 23744 3732 23796 3738
rect 23744 3674 23796 3680
rect 23560 3664 23612 3670
rect 23848 3618 23876 5879
rect 23940 4282 23968 7142
rect 24032 6730 24060 7346
rect 24020 6724 24072 6730
rect 24020 6666 24072 6672
rect 24001 6556 24297 6576
rect 24057 6554 24081 6556
rect 24137 6554 24161 6556
rect 24217 6554 24241 6556
rect 24079 6502 24081 6554
rect 24143 6502 24155 6554
rect 24217 6502 24219 6554
rect 24057 6500 24081 6502
rect 24137 6500 24161 6502
rect 24217 6500 24241 6502
rect 24001 6480 24297 6500
rect 24001 5468 24297 5488
rect 24057 5466 24081 5468
rect 24137 5466 24161 5468
rect 24217 5466 24241 5468
rect 24079 5414 24081 5466
rect 24143 5414 24155 5466
rect 24217 5414 24219 5466
rect 24057 5412 24081 5414
rect 24137 5412 24161 5414
rect 24217 5412 24241 5414
rect 24001 5392 24297 5412
rect 24400 5370 24428 9959
rect 24480 9920 24532 9926
rect 24480 9862 24532 9868
rect 24492 9654 24520 9862
rect 24480 9648 24532 9654
rect 24480 9590 24532 9596
rect 24478 8936 24534 8945
rect 24478 8871 24534 8880
rect 24492 6882 24520 8871
rect 24584 7954 24612 9982
rect 24768 9722 24796 10134
rect 24938 10095 24994 10104
rect 24756 9716 24808 9722
rect 24756 9658 24808 9664
rect 24664 8832 24716 8838
rect 24664 8774 24716 8780
rect 24676 8430 24704 8774
rect 24664 8424 24716 8430
rect 24664 8366 24716 8372
rect 24676 8090 24704 8366
rect 24664 8084 24716 8090
rect 24664 8026 24716 8032
rect 24572 7948 24624 7954
rect 24572 7890 24624 7896
rect 24584 7546 24612 7890
rect 24664 7880 24716 7886
rect 24664 7822 24716 7828
rect 24938 7848 24994 7857
rect 24572 7540 24624 7546
rect 24572 7482 24624 7488
rect 24492 6866 24612 6882
rect 24492 6860 24624 6866
rect 24492 6854 24572 6860
rect 24492 6440 24520 6854
rect 24572 6802 24624 6808
rect 24572 6452 24624 6458
rect 24492 6412 24572 6440
rect 24572 6394 24624 6400
rect 24480 5568 24532 5574
rect 24480 5510 24532 5516
rect 24388 5364 24440 5370
rect 24388 5306 24440 5312
rect 24492 5234 24520 5510
rect 24480 5228 24532 5234
rect 24480 5170 24532 5176
rect 24386 4856 24442 4865
rect 24676 4826 24704 7822
rect 24938 7783 24940 7792
rect 24992 7783 24994 7792
rect 24940 7754 24992 7760
rect 25674 7712 25730 7721
rect 25674 7647 25730 7656
rect 25688 7546 25716 7647
rect 25964 7546 25992 22335
rect 26320 15360 26372 15366
rect 26320 15302 26372 15308
rect 25676 7540 25728 7546
rect 25676 7482 25728 7488
rect 25952 7540 26004 7546
rect 25952 7482 26004 7488
rect 25688 7342 25716 7482
rect 25676 7336 25728 7342
rect 25676 7278 25728 7284
rect 25216 7200 25268 7206
rect 25216 7142 25268 7148
rect 24848 6724 24900 6730
rect 24848 6666 24900 6672
rect 24860 6390 24888 6666
rect 24940 6656 24992 6662
rect 24940 6598 24992 6604
rect 24848 6384 24900 6390
rect 24848 6326 24900 6332
rect 24754 4992 24810 5001
rect 24754 4927 24810 4936
rect 24664 4820 24716 4826
rect 24386 4791 24442 4800
rect 24001 4380 24297 4400
rect 24057 4378 24081 4380
rect 24137 4378 24161 4380
rect 24217 4378 24241 4380
rect 24079 4326 24081 4378
rect 24143 4326 24155 4378
rect 24217 4326 24219 4378
rect 24057 4324 24081 4326
rect 24137 4324 24161 4326
rect 24217 4324 24241 4326
rect 24001 4304 24297 4324
rect 24400 4321 24428 4791
rect 24584 4780 24664 4808
rect 24386 4312 24442 4321
rect 23928 4276 23980 4282
rect 24386 4247 24442 4256
rect 23928 4218 23980 4224
rect 24480 4072 24532 4078
rect 24480 4014 24532 4020
rect 23560 3606 23612 3612
rect 23466 3360 23522 3369
rect 23466 3295 23522 3304
rect 23192 3188 23244 3194
rect 23192 3130 23244 3136
rect 23204 2922 23232 3130
rect 23480 2990 23508 3295
rect 23572 3058 23600 3606
rect 23664 3590 23876 3618
rect 23560 3052 23612 3058
rect 23560 2994 23612 3000
rect 23468 2984 23520 2990
rect 23374 2952 23430 2961
rect 23192 2916 23244 2922
rect 23468 2926 23520 2932
rect 23374 2887 23430 2896
rect 23192 2858 23244 2864
rect 23008 2644 23060 2650
rect 23008 2586 23060 2592
rect 23388 480 23416 2887
rect 23480 2310 23508 2926
rect 23468 2304 23520 2310
rect 23468 2246 23520 2252
rect 23480 1465 23508 2246
rect 23664 1873 23692 3590
rect 24001 3292 24297 3312
rect 24057 3290 24081 3292
rect 24137 3290 24161 3292
rect 24217 3290 24241 3292
rect 24079 3238 24081 3290
rect 24143 3238 24155 3290
rect 24217 3238 24219 3290
rect 24057 3236 24081 3238
rect 24137 3236 24161 3238
rect 24217 3236 24241 3238
rect 24001 3216 24297 3236
rect 23926 3088 23982 3097
rect 23926 3023 23928 3032
rect 23980 3023 23982 3032
rect 23928 2994 23980 3000
rect 23836 2916 23888 2922
rect 23836 2858 23888 2864
rect 23650 1864 23706 1873
rect 23650 1799 23706 1808
rect 23466 1456 23522 1465
rect 23466 1391 23522 1400
rect 6 0 62 480
rect 650 0 706 480
rect 1294 0 1350 480
rect 1938 0 1994 480
rect 2582 0 2638 480
rect 3226 0 3282 480
rect 3870 0 3926 480
rect 4514 0 4570 480
rect 5158 0 5214 480
rect 5802 0 5858 480
rect 6446 0 6502 480
rect 7090 0 7146 480
rect 7734 0 7790 480
rect 8378 0 8434 480
rect 9022 0 9078 480
rect 9758 0 9814 480
rect 10402 0 10458 480
rect 11046 0 11102 480
rect 11690 0 11746 480
rect 12334 0 12390 480
rect 12978 0 13034 480
rect 13622 0 13678 480
rect 14266 0 14322 480
rect 14910 0 14966 480
rect 15554 0 15610 480
rect 16198 0 16254 480
rect 16842 0 16898 480
rect 17486 0 17542 480
rect 18130 0 18186 480
rect 18866 0 18922 480
rect 19510 0 19566 480
rect 20154 0 20210 480
rect 20798 0 20854 480
rect 21442 0 21498 480
rect 22086 0 22142 480
rect 22730 0 22786 480
rect 23374 0 23430 480
rect 23848 377 23876 2858
rect 24202 2680 24258 2689
rect 24202 2615 24204 2624
rect 24256 2615 24258 2624
rect 24204 2586 24256 2592
rect 24112 2508 24164 2514
rect 24112 2450 24164 2456
rect 24124 2417 24152 2450
rect 24110 2408 24166 2417
rect 24110 2343 24166 2352
rect 24001 2204 24297 2224
rect 24057 2202 24081 2204
rect 24137 2202 24161 2204
rect 24217 2202 24241 2204
rect 24079 2150 24081 2202
rect 24143 2150 24155 2202
rect 24217 2150 24219 2202
rect 24057 2148 24081 2150
rect 24137 2148 24161 2150
rect 24217 2148 24241 2150
rect 24001 2128 24297 2148
rect 24020 2032 24072 2038
rect 24020 1974 24072 1980
rect 24032 480 24060 1974
rect 24492 921 24520 4014
rect 24584 4010 24612 4780
rect 24664 4762 24716 4768
rect 24768 4690 24796 4927
rect 24756 4684 24808 4690
rect 24756 4626 24808 4632
rect 24664 4480 24716 4486
rect 24664 4422 24716 4428
rect 24676 4214 24704 4422
rect 24768 4282 24796 4626
rect 24952 4570 24980 6598
rect 25032 4752 25084 4758
rect 25032 4694 25084 4700
rect 24860 4542 24980 4570
rect 24756 4276 24808 4282
rect 24756 4218 24808 4224
rect 24664 4208 24716 4214
rect 24664 4150 24716 4156
rect 24572 4004 24624 4010
rect 24572 3946 24624 3952
rect 24572 3596 24624 3602
rect 24572 3538 24624 3544
rect 24584 2922 24612 3538
rect 24860 3505 24888 4542
rect 24846 3496 24902 3505
rect 24846 3431 24902 3440
rect 24664 3392 24716 3398
rect 24664 3334 24716 3340
rect 24676 3058 24704 3334
rect 25044 3233 25072 4694
rect 25030 3224 25086 3233
rect 25030 3159 25086 3168
rect 24664 3052 24716 3058
rect 24664 2994 24716 3000
rect 24662 2952 24718 2961
rect 24572 2916 24624 2922
rect 24662 2887 24718 2896
rect 24572 2858 24624 2864
rect 24572 2440 24624 2446
rect 24572 2382 24624 2388
rect 24584 1737 24612 2382
rect 24570 1728 24626 1737
rect 24570 1663 24626 1672
rect 24478 912 24534 921
rect 24478 847 24534 856
rect 24676 480 24704 2887
rect 25124 2848 25176 2854
rect 25122 2816 25124 2825
rect 25176 2816 25178 2825
rect 25122 2751 25178 2760
rect 25228 610 25256 7142
rect 25952 6112 26004 6118
rect 25952 6054 26004 6060
rect 25964 5030 25992 6054
rect 25308 5024 25360 5030
rect 25308 4966 25360 4972
rect 25952 5024 26004 5030
rect 25952 4966 26004 4972
rect 25320 3641 25348 4966
rect 25306 3632 25362 3641
rect 25306 3567 25362 3576
rect 25768 2848 25820 2854
rect 25964 2836 25992 4966
rect 25820 2808 25992 2836
rect 25768 2790 25820 2796
rect 25780 2650 25808 2790
rect 25768 2644 25820 2650
rect 25768 2586 25820 2592
rect 25306 2000 25362 2009
rect 25306 1935 25362 1944
rect 25216 604 25268 610
rect 25216 546 25268 552
rect 25320 480 25348 1935
rect 26332 610 26360 15302
rect 26596 7540 26648 7546
rect 26596 7482 26648 7488
rect 25952 604 26004 610
rect 25952 546 26004 552
rect 26320 604 26372 610
rect 26320 546 26372 552
rect 25964 480 25992 546
rect 26608 480 26636 7482
rect 27238 2816 27294 2825
rect 27238 2751 27294 2760
rect 27252 480 27280 2751
rect 23834 368 23890 377
rect 23834 303 23890 312
rect 24018 0 24074 480
rect 24662 0 24718 480
rect 25306 0 25362 480
rect 25950 0 26006 480
rect 26594 0 26650 480
rect 27238 0 27294 480
<< via2 >>
rect 5334 25050 5390 25052
rect 5414 25050 5470 25052
rect 5494 25050 5550 25052
rect 5574 25050 5630 25052
rect 5334 24998 5360 25050
rect 5360 24998 5390 25050
rect 5414 24998 5424 25050
rect 5424 24998 5470 25050
rect 5494 24998 5540 25050
rect 5540 24998 5550 25050
rect 5574 24998 5604 25050
rect 5604 24998 5630 25050
rect 5334 24996 5390 24998
rect 5414 24996 5470 24998
rect 5494 24996 5550 24998
rect 5574 24996 5630 24998
rect 5334 23962 5390 23964
rect 5414 23962 5470 23964
rect 5494 23962 5550 23964
rect 5574 23962 5630 23964
rect 5334 23910 5360 23962
rect 5360 23910 5390 23962
rect 5414 23910 5424 23962
rect 5424 23910 5470 23962
rect 5494 23910 5540 23962
rect 5540 23910 5550 23962
rect 5574 23910 5604 23962
rect 5604 23910 5630 23962
rect 5334 23908 5390 23910
rect 5414 23908 5470 23910
rect 5494 23908 5550 23910
rect 5574 23908 5630 23910
rect 5334 22874 5390 22876
rect 5414 22874 5470 22876
rect 5494 22874 5550 22876
rect 5574 22874 5630 22876
rect 5334 22822 5360 22874
rect 5360 22822 5390 22874
rect 5414 22822 5424 22874
rect 5424 22822 5470 22874
rect 5494 22822 5540 22874
rect 5540 22822 5550 22874
rect 5574 22822 5604 22874
rect 5604 22822 5630 22874
rect 5334 22820 5390 22822
rect 5414 22820 5470 22822
rect 5494 22820 5550 22822
rect 5574 22820 5630 22822
rect 5334 21786 5390 21788
rect 5414 21786 5470 21788
rect 5494 21786 5550 21788
rect 5574 21786 5630 21788
rect 5334 21734 5360 21786
rect 5360 21734 5390 21786
rect 5414 21734 5424 21786
rect 5424 21734 5470 21786
rect 5494 21734 5540 21786
rect 5540 21734 5550 21786
rect 5574 21734 5604 21786
rect 5604 21734 5630 21786
rect 5334 21732 5390 21734
rect 5414 21732 5470 21734
rect 5494 21732 5550 21734
rect 5574 21732 5630 21734
rect 5334 20698 5390 20700
rect 5414 20698 5470 20700
rect 5494 20698 5550 20700
rect 5574 20698 5630 20700
rect 5334 20646 5360 20698
rect 5360 20646 5390 20698
rect 5414 20646 5424 20698
rect 5424 20646 5470 20698
rect 5494 20646 5540 20698
rect 5540 20646 5550 20698
rect 5574 20646 5604 20698
rect 5604 20646 5630 20698
rect 5334 20644 5390 20646
rect 5414 20644 5470 20646
rect 5494 20644 5550 20646
rect 5574 20644 5630 20646
rect 5334 19610 5390 19612
rect 5414 19610 5470 19612
rect 5494 19610 5550 19612
rect 5574 19610 5630 19612
rect 5334 19558 5360 19610
rect 5360 19558 5390 19610
rect 5414 19558 5424 19610
rect 5424 19558 5470 19610
rect 5494 19558 5540 19610
rect 5540 19558 5550 19610
rect 5574 19558 5604 19610
rect 5604 19558 5630 19610
rect 5334 19556 5390 19558
rect 5414 19556 5470 19558
rect 5494 19556 5550 19558
rect 5574 19556 5630 19558
rect 5334 18522 5390 18524
rect 5414 18522 5470 18524
rect 5494 18522 5550 18524
rect 5574 18522 5630 18524
rect 5334 18470 5360 18522
rect 5360 18470 5390 18522
rect 5414 18470 5424 18522
rect 5424 18470 5470 18522
rect 5494 18470 5540 18522
rect 5540 18470 5550 18522
rect 5574 18470 5604 18522
rect 5604 18470 5630 18522
rect 5334 18468 5390 18470
rect 5414 18468 5470 18470
rect 5494 18468 5550 18470
rect 5574 18468 5630 18470
rect 5334 17434 5390 17436
rect 5414 17434 5470 17436
rect 5494 17434 5550 17436
rect 5574 17434 5630 17436
rect 5334 17382 5360 17434
rect 5360 17382 5390 17434
rect 5414 17382 5424 17434
rect 5424 17382 5470 17434
rect 5494 17382 5540 17434
rect 5540 17382 5550 17434
rect 5574 17382 5604 17434
rect 5604 17382 5630 17434
rect 5334 17380 5390 17382
rect 5414 17380 5470 17382
rect 5494 17380 5550 17382
rect 5574 17380 5630 17382
rect 7550 16904 7606 16960
rect 5334 16346 5390 16348
rect 5414 16346 5470 16348
rect 5494 16346 5550 16348
rect 5574 16346 5630 16348
rect 5334 16294 5360 16346
rect 5360 16294 5390 16346
rect 5414 16294 5424 16346
rect 5424 16294 5470 16346
rect 5494 16294 5540 16346
rect 5540 16294 5550 16346
rect 5574 16294 5604 16346
rect 5604 16294 5630 16346
rect 5334 16292 5390 16294
rect 5414 16292 5470 16294
rect 5494 16292 5550 16294
rect 5574 16292 5630 16294
rect 5334 15258 5390 15260
rect 5414 15258 5470 15260
rect 5494 15258 5550 15260
rect 5574 15258 5630 15260
rect 5334 15206 5360 15258
rect 5360 15206 5390 15258
rect 5414 15206 5424 15258
rect 5424 15206 5470 15258
rect 5494 15206 5540 15258
rect 5540 15206 5550 15258
rect 5574 15206 5604 15258
rect 5604 15206 5630 15258
rect 5334 15204 5390 15206
rect 5414 15204 5470 15206
rect 5494 15204 5550 15206
rect 5574 15204 5630 15206
rect 3778 14456 3834 14512
rect 5334 14170 5390 14172
rect 5414 14170 5470 14172
rect 5494 14170 5550 14172
rect 5574 14170 5630 14172
rect 5334 14118 5360 14170
rect 5360 14118 5390 14170
rect 5414 14118 5424 14170
rect 5424 14118 5470 14170
rect 5494 14118 5540 14170
rect 5540 14118 5550 14170
rect 5574 14118 5604 14170
rect 5604 14118 5630 14170
rect 5334 14116 5390 14118
rect 5414 14116 5470 14118
rect 5494 14116 5550 14118
rect 5574 14116 5630 14118
rect 5334 13082 5390 13084
rect 5414 13082 5470 13084
rect 5494 13082 5550 13084
rect 5574 13082 5630 13084
rect 5334 13030 5360 13082
rect 5360 13030 5390 13082
rect 5414 13030 5424 13082
rect 5424 13030 5470 13082
rect 5494 13030 5540 13082
rect 5540 13030 5550 13082
rect 5574 13030 5604 13082
rect 5604 13030 5630 13082
rect 5334 13028 5390 13030
rect 5414 13028 5470 13030
rect 5494 13028 5550 13030
rect 5574 13028 5630 13030
rect 3870 12688 3926 12744
rect 1294 8336 1350 8392
rect 650 6296 706 6352
rect 6 4120 62 4176
rect 5334 11994 5390 11996
rect 5414 11994 5470 11996
rect 5494 11994 5550 11996
rect 5574 11994 5630 11996
rect 5334 11942 5360 11994
rect 5360 11942 5390 11994
rect 5414 11942 5424 11994
rect 5424 11942 5470 11994
rect 5494 11942 5540 11994
rect 5540 11942 5550 11994
rect 5574 11942 5604 11994
rect 5604 11942 5630 11994
rect 5334 11940 5390 11942
rect 5414 11940 5470 11942
rect 5494 11940 5550 11942
rect 5574 11940 5630 11942
rect 5334 10906 5390 10908
rect 5414 10906 5470 10908
rect 5494 10906 5550 10908
rect 5574 10906 5630 10908
rect 5334 10854 5360 10906
rect 5360 10854 5390 10906
rect 5414 10854 5424 10906
rect 5424 10854 5470 10906
rect 5494 10854 5540 10906
rect 5540 10854 5550 10906
rect 5574 10854 5604 10906
rect 5604 10854 5630 10906
rect 5334 10852 5390 10854
rect 5414 10852 5470 10854
rect 5494 10852 5550 10854
rect 5574 10852 5630 10854
rect 5334 9818 5390 9820
rect 5414 9818 5470 9820
rect 5494 9818 5550 9820
rect 5574 9818 5630 9820
rect 5334 9766 5360 9818
rect 5360 9766 5390 9818
rect 5414 9766 5424 9818
rect 5424 9766 5470 9818
rect 5494 9766 5540 9818
rect 5540 9766 5550 9818
rect 5574 9766 5604 9818
rect 5604 9766 5630 9818
rect 5334 9764 5390 9766
rect 5414 9764 5470 9766
rect 5494 9764 5550 9766
rect 5574 9764 5630 9766
rect 5802 9424 5858 9480
rect 5334 8730 5390 8732
rect 5414 8730 5470 8732
rect 5494 8730 5550 8732
rect 5574 8730 5630 8732
rect 5334 8678 5360 8730
rect 5360 8678 5390 8730
rect 5414 8678 5424 8730
rect 5424 8678 5470 8730
rect 5494 8678 5540 8730
rect 5540 8678 5550 8730
rect 5574 8678 5604 8730
rect 5604 8678 5630 8730
rect 5334 8676 5390 8678
rect 5414 8676 5470 8678
rect 5494 8676 5550 8678
rect 5574 8676 5630 8678
rect 5066 7928 5122 7984
rect 1938 7248 1994 7304
rect 4514 5208 4570 5264
rect 3226 4120 3282 4176
rect 2582 3848 2638 3904
rect 3962 3440 4018 3496
rect 5334 7642 5390 7644
rect 5414 7642 5470 7644
rect 5494 7642 5550 7644
rect 5574 7642 5630 7644
rect 5334 7590 5360 7642
rect 5360 7590 5390 7642
rect 5414 7590 5424 7642
rect 5424 7590 5470 7642
rect 5494 7590 5540 7642
rect 5540 7590 5550 7642
rect 5574 7590 5604 7642
rect 5604 7590 5630 7642
rect 5334 7588 5390 7590
rect 5414 7588 5470 7590
rect 5494 7588 5550 7590
rect 5574 7588 5630 7590
rect 5066 4392 5122 4448
rect 5334 6554 5390 6556
rect 5414 6554 5470 6556
rect 5494 6554 5550 6556
rect 5574 6554 5630 6556
rect 5334 6502 5360 6554
rect 5360 6502 5390 6554
rect 5414 6502 5424 6554
rect 5424 6502 5470 6554
rect 5494 6502 5540 6554
rect 5540 6502 5550 6554
rect 5574 6502 5604 6554
rect 5604 6502 5630 6554
rect 5334 6500 5390 6502
rect 5414 6500 5470 6502
rect 5494 6500 5550 6502
rect 5574 6500 5630 6502
rect 5334 5466 5390 5468
rect 5414 5466 5470 5468
rect 5494 5466 5550 5468
rect 5574 5466 5630 5468
rect 5334 5414 5360 5466
rect 5360 5414 5390 5466
rect 5414 5414 5424 5466
rect 5424 5414 5470 5466
rect 5494 5414 5540 5466
rect 5540 5414 5550 5466
rect 5574 5414 5604 5466
rect 5604 5414 5630 5466
rect 5334 5412 5390 5414
rect 5414 5412 5470 5414
rect 5494 5412 5550 5414
rect 5574 5412 5630 5414
rect 5334 4378 5390 4380
rect 5414 4378 5470 4380
rect 5494 4378 5550 4380
rect 5574 4378 5630 4380
rect 5334 4326 5360 4378
rect 5360 4326 5390 4378
rect 5414 4326 5424 4378
rect 5424 4326 5470 4378
rect 5494 4326 5540 4378
rect 5540 4326 5550 4378
rect 5574 4326 5604 4378
rect 5604 4326 5630 4378
rect 5334 4324 5390 4326
rect 5414 4324 5470 4326
rect 5494 4324 5550 4326
rect 5574 4324 5630 4326
rect 5334 3290 5390 3292
rect 5414 3290 5470 3292
rect 5494 3290 5550 3292
rect 5574 3290 5630 3292
rect 5334 3238 5360 3290
rect 5360 3238 5390 3290
rect 5414 3238 5424 3290
rect 5424 3238 5470 3290
rect 5494 3238 5540 3290
rect 5540 3238 5550 3290
rect 5574 3238 5604 3290
rect 5604 3238 5630 3290
rect 5334 3236 5390 3238
rect 5414 3236 5470 3238
rect 5494 3236 5550 3238
rect 5574 3236 5630 3238
rect 5334 2202 5390 2204
rect 5414 2202 5470 2204
rect 5494 2202 5550 2204
rect 5574 2202 5630 2204
rect 5334 2150 5360 2202
rect 5360 2150 5390 2202
rect 5414 2150 5424 2202
rect 5424 2150 5470 2202
rect 5494 2150 5540 2202
rect 5540 2150 5550 2202
rect 5574 2150 5604 2202
rect 5604 2150 5630 2202
rect 5334 2148 5390 2150
rect 5414 2148 5470 2150
rect 5494 2148 5550 2150
rect 5574 2148 5630 2150
rect 7090 4936 7146 4992
rect 6446 4392 6502 4448
rect 7642 7520 7698 7576
rect 10001 25594 10057 25596
rect 10081 25594 10137 25596
rect 10161 25594 10217 25596
rect 10241 25594 10297 25596
rect 10001 25542 10027 25594
rect 10027 25542 10057 25594
rect 10081 25542 10091 25594
rect 10091 25542 10137 25594
rect 10161 25542 10207 25594
rect 10207 25542 10217 25594
rect 10241 25542 10271 25594
rect 10271 25542 10297 25594
rect 10001 25540 10057 25542
rect 10081 25540 10137 25542
rect 10161 25540 10217 25542
rect 10241 25540 10297 25542
rect 10001 24506 10057 24508
rect 10081 24506 10137 24508
rect 10161 24506 10217 24508
rect 10241 24506 10297 24508
rect 10001 24454 10027 24506
rect 10027 24454 10057 24506
rect 10081 24454 10091 24506
rect 10091 24454 10137 24506
rect 10161 24454 10207 24506
rect 10207 24454 10217 24506
rect 10241 24454 10271 24506
rect 10271 24454 10297 24506
rect 10001 24452 10057 24454
rect 10081 24452 10137 24454
rect 10161 24452 10217 24454
rect 10241 24452 10297 24454
rect 10678 23568 10734 23624
rect 10001 23418 10057 23420
rect 10081 23418 10137 23420
rect 10161 23418 10217 23420
rect 10241 23418 10297 23420
rect 10001 23366 10027 23418
rect 10027 23366 10057 23418
rect 10081 23366 10091 23418
rect 10091 23366 10137 23418
rect 10161 23366 10207 23418
rect 10207 23366 10217 23418
rect 10241 23366 10271 23418
rect 10271 23366 10297 23418
rect 10001 23364 10057 23366
rect 10081 23364 10137 23366
rect 10161 23364 10217 23366
rect 10241 23364 10297 23366
rect 10586 22480 10642 22536
rect 10001 22330 10057 22332
rect 10081 22330 10137 22332
rect 10161 22330 10217 22332
rect 10241 22330 10297 22332
rect 10001 22278 10027 22330
rect 10027 22278 10057 22330
rect 10081 22278 10091 22330
rect 10091 22278 10137 22330
rect 10161 22278 10207 22330
rect 10207 22278 10217 22330
rect 10241 22278 10271 22330
rect 10271 22278 10297 22330
rect 10001 22276 10057 22278
rect 10081 22276 10137 22278
rect 10161 22276 10217 22278
rect 10241 22276 10297 22278
rect 8470 7792 8526 7848
rect 7734 6568 7790 6624
rect 7826 5636 7882 5672
rect 7826 5616 7828 5636
rect 7828 5616 7880 5636
rect 7880 5616 7882 5636
rect 8010 4972 8012 4992
rect 8012 4972 8064 4992
rect 8064 4972 8066 4992
rect 8010 4936 8066 4972
rect 8286 3984 8342 4040
rect 8378 3848 8434 3904
rect 7734 3712 7790 3768
rect 7182 2916 7238 2952
rect 7182 2896 7184 2916
rect 7184 2896 7236 2916
rect 7236 2896 7238 2916
rect 9206 7420 9208 7440
rect 9208 7420 9260 7440
rect 9260 7420 9262 7440
rect 9206 7384 9262 7420
rect 10001 21242 10057 21244
rect 10081 21242 10137 21244
rect 10161 21242 10217 21244
rect 10241 21242 10297 21244
rect 10001 21190 10027 21242
rect 10027 21190 10057 21242
rect 10081 21190 10091 21242
rect 10091 21190 10137 21242
rect 10161 21190 10207 21242
rect 10207 21190 10217 21242
rect 10241 21190 10271 21242
rect 10271 21190 10297 21242
rect 10001 21188 10057 21190
rect 10081 21188 10137 21190
rect 10161 21188 10217 21190
rect 10241 21188 10297 21190
rect 9666 20984 9722 21040
rect 10001 20154 10057 20156
rect 10081 20154 10137 20156
rect 10161 20154 10217 20156
rect 10241 20154 10297 20156
rect 10001 20102 10027 20154
rect 10027 20102 10057 20154
rect 10081 20102 10091 20154
rect 10091 20102 10137 20154
rect 10161 20102 10207 20154
rect 10207 20102 10217 20154
rect 10241 20102 10271 20154
rect 10271 20102 10297 20154
rect 10001 20100 10057 20102
rect 10081 20100 10137 20102
rect 10161 20100 10217 20102
rect 10241 20100 10297 20102
rect 10001 19066 10057 19068
rect 10081 19066 10137 19068
rect 10161 19066 10217 19068
rect 10241 19066 10297 19068
rect 10001 19014 10027 19066
rect 10027 19014 10057 19066
rect 10081 19014 10091 19066
rect 10091 19014 10137 19066
rect 10161 19014 10207 19066
rect 10207 19014 10217 19066
rect 10241 19014 10271 19066
rect 10271 19014 10297 19066
rect 10001 19012 10057 19014
rect 10081 19012 10137 19014
rect 10161 19012 10217 19014
rect 10241 19012 10297 19014
rect 10001 17978 10057 17980
rect 10081 17978 10137 17980
rect 10161 17978 10217 17980
rect 10241 17978 10297 17980
rect 10001 17926 10027 17978
rect 10027 17926 10057 17978
rect 10081 17926 10091 17978
rect 10091 17926 10137 17978
rect 10161 17926 10207 17978
rect 10207 17926 10217 17978
rect 10241 17926 10271 17978
rect 10271 17926 10297 17978
rect 10001 17924 10057 17926
rect 10081 17924 10137 17926
rect 10161 17924 10217 17926
rect 10241 17924 10297 17926
rect 9850 16940 9852 16960
rect 9852 16940 9904 16960
rect 9904 16940 9906 16960
rect 9850 16904 9906 16940
rect 10001 16890 10057 16892
rect 10081 16890 10137 16892
rect 10161 16890 10217 16892
rect 10241 16890 10297 16892
rect 10001 16838 10027 16890
rect 10027 16838 10057 16890
rect 10081 16838 10091 16890
rect 10091 16838 10137 16890
rect 10161 16838 10207 16890
rect 10207 16838 10217 16890
rect 10241 16838 10271 16890
rect 10271 16838 10297 16890
rect 10001 16836 10057 16838
rect 10081 16836 10137 16838
rect 10161 16836 10217 16838
rect 10241 16836 10297 16838
rect 10001 15802 10057 15804
rect 10081 15802 10137 15804
rect 10161 15802 10217 15804
rect 10241 15802 10297 15804
rect 10001 15750 10027 15802
rect 10027 15750 10057 15802
rect 10081 15750 10091 15802
rect 10091 15750 10137 15802
rect 10161 15750 10207 15802
rect 10207 15750 10217 15802
rect 10241 15750 10271 15802
rect 10271 15750 10297 15802
rect 10001 15748 10057 15750
rect 10081 15748 10137 15750
rect 10161 15748 10217 15750
rect 10241 15748 10297 15750
rect 10001 14714 10057 14716
rect 10081 14714 10137 14716
rect 10161 14714 10217 14716
rect 10241 14714 10297 14716
rect 10001 14662 10027 14714
rect 10027 14662 10057 14714
rect 10081 14662 10091 14714
rect 10091 14662 10137 14714
rect 10161 14662 10207 14714
rect 10207 14662 10217 14714
rect 10241 14662 10271 14714
rect 10271 14662 10297 14714
rect 10001 14660 10057 14662
rect 10081 14660 10137 14662
rect 10161 14660 10217 14662
rect 10241 14660 10297 14662
rect 10001 13626 10057 13628
rect 10081 13626 10137 13628
rect 10161 13626 10217 13628
rect 10241 13626 10297 13628
rect 10001 13574 10027 13626
rect 10027 13574 10057 13626
rect 10081 13574 10091 13626
rect 10091 13574 10137 13626
rect 10161 13574 10207 13626
rect 10207 13574 10217 13626
rect 10241 13574 10271 13626
rect 10271 13574 10297 13626
rect 10001 13572 10057 13574
rect 10081 13572 10137 13574
rect 10161 13572 10217 13574
rect 10241 13572 10297 13574
rect 10001 12538 10057 12540
rect 10081 12538 10137 12540
rect 10161 12538 10217 12540
rect 10241 12538 10297 12540
rect 10001 12486 10027 12538
rect 10027 12486 10057 12538
rect 10081 12486 10091 12538
rect 10091 12486 10137 12538
rect 10161 12486 10207 12538
rect 10207 12486 10217 12538
rect 10241 12486 10271 12538
rect 10271 12486 10297 12538
rect 10001 12484 10057 12486
rect 10081 12484 10137 12486
rect 10161 12484 10217 12486
rect 10241 12484 10297 12486
rect 10001 11450 10057 11452
rect 10081 11450 10137 11452
rect 10161 11450 10217 11452
rect 10241 11450 10297 11452
rect 10001 11398 10027 11450
rect 10027 11398 10057 11450
rect 10081 11398 10091 11450
rect 10091 11398 10137 11450
rect 10161 11398 10207 11450
rect 10207 11398 10217 11450
rect 10241 11398 10271 11450
rect 10271 11398 10297 11450
rect 10001 11396 10057 11398
rect 10081 11396 10137 11398
rect 10161 11396 10217 11398
rect 10241 11396 10297 11398
rect 10001 10362 10057 10364
rect 10081 10362 10137 10364
rect 10161 10362 10217 10364
rect 10241 10362 10297 10364
rect 10001 10310 10027 10362
rect 10027 10310 10057 10362
rect 10081 10310 10091 10362
rect 10091 10310 10137 10362
rect 10161 10310 10207 10362
rect 10207 10310 10217 10362
rect 10241 10310 10271 10362
rect 10271 10310 10297 10362
rect 10001 10308 10057 10310
rect 10081 10308 10137 10310
rect 10161 10308 10217 10310
rect 10241 10308 10297 10310
rect 10001 9274 10057 9276
rect 10081 9274 10137 9276
rect 10161 9274 10217 9276
rect 10241 9274 10297 9276
rect 10001 9222 10027 9274
rect 10027 9222 10057 9274
rect 10081 9222 10091 9274
rect 10091 9222 10137 9274
rect 10161 9222 10207 9274
rect 10207 9222 10217 9274
rect 10241 9222 10271 9274
rect 10271 9222 10297 9274
rect 10001 9220 10057 9222
rect 10081 9220 10137 9222
rect 10161 9220 10217 9222
rect 10241 9220 10297 9222
rect 12242 21392 12298 21448
rect 11138 19760 11194 19816
rect 10001 8186 10057 8188
rect 10081 8186 10137 8188
rect 10161 8186 10217 8188
rect 10241 8186 10297 8188
rect 10001 8134 10027 8186
rect 10027 8134 10057 8186
rect 10081 8134 10091 8186
rect 10091 8134 10137 8186
rect 10161 8134 10207 8186
rect 10207 8134 10217 8186
rect 10241 8134 10271 8186
rect 10271 8134 10297 8186
rect 10001 8132 10057 8134
rect 10081 8132 10137 8134
rect 10161 8132 10217 8134
rect 10241 8132 10297 8134
rect 11874 8880 11930 8936
rect 10310 7268 10366 7304
rect 10310 7248 10312 7268
rect 10312 7248 10364 7268
rect 10364 7248 10366 7268
rect 10001 7098 10057 7100
rect 10081 7098 10137 7100
rect 10161 7098 10217 7100
rect 10241 7098 10297 7100
rect 10001 7046 10027 7098
rect 10027 7046 10057 7098
rect 10081 7046 10091 7098
rect 10091 7046 10137 7098
rect 10161 7046 10207 7098
rect 10207 7046 10217 7098
rect 10241 7046 10271 7098
rect 10271 7046 10297 7098
rect 10001 7044 10057 7046
rect 10081 7044 10137 7046
rect 10161 7044 10217 7046
rect 10241 7044 10297 7046
rect 10770 6704 10826 6760
rect 10001 6010 10057 6012
rect 10081 6010 10137 6012
rect 10161 6010 10217 6012
rect 10241 6010 10297 6012
rect 10001 5958 10027 6010
rect 10027 5958 10057 6010
rect 10081 5958 10091 6010
rect 10091 5958 10137 6010
rect 10161 5958 10207 6010
rect 10207 5958 10217 6010
rect 10241 5958 10271 6010
rect 10271 5958 10297 6010
rect 10001 5956 10057 5958
rect 10081 5956 10137 5958
rect 10161 5956 10217 5958
rect 10241 5956 10297 5958
rect 8838 4528 8894 4584
rect 7826 2372 7882 2408
rect 7826 2352 7828 2372
rect 7828 2352 7880 2372
rect 7880 2352 7882 2372
rect 8286 2216 8342 2272
rect 8378 2080 8434 2136
rect 8194 1672 8250 1728
rect 11506 5616 11562 5672
rect 10954 5092 11010 5128
rect 10954 5072 10956 5092
rect 10956 5072 11008 5092
rect 11008 5072 11010 5092
rect 10001 4922 10057 4924
rect 10081 4922 10137 4924
rect 10161 4922 10217 4924
rect 10241 4922 10297 4924
rect 10001 4870 10027 4922
rect 10027 4870 10057 4922
rect 10081 4870 10091 4922
rect 10091 4870 10137 4922
rect 10161 4870 10207 4922
rect 10207 4870 10217 4922
rect 10241 4870 10271 4922
rect 10271 4870 10297 4922
rect 10001 4868 10057 4870
rect 10081 4868 10137 4870
rect 10161 4868 10217 4870
rect 10241 4868 10297 4870
rect 9758 4120 9814 4176
rect 8930 3712 8986 3768
rect 9022 3576 9078 3632
rect 8654 1944 8710 2000
rect 8562 1808 8618 1864
rect 8470 1536 8526 1592
rect 10402 3848 10458 3904
rect 10001 3834 10057 3836
rect 10081 3834 10137 3836
rect 10161 3834 10217 3836
rect 10241 3834 10297 3836
rect 10001 3782 10027 3834
rect 10027 3782 10057 3834
rect 10081 3782 10091 3834
rect 10091 3782 10137 3834
rect 10161 3782 10207 3834
rect 10207 3782 10217 3834
rect 10241 3782 10271 3834
rect 10271 3782 10297 3834
rect 10001 3780 10057 3782
rect 10081 3780 10137 3782
rect 10161 3780 10217 3782
rect 10241 3780 10297 3782
rect 9850 3304 9906 3360
rect 10001 2746 10057 2748
rect 10081 2746 10137 2748
rect 10161 2746 10217 2748
rect 10241 2746 10297 2748
rect 10001 2694 10027 2746
rect 10027 2694 10057 2746
rect 10081 2694 10091 2746
rect 10091 2694 10137 2746
rect 10161 2694 10207 2746
rect 10207 2694 10217 2746
rect 10241 2694 10271 2746
rect 10271 2694 10297 2746
rect 10001 2692 10057 2694
rect 10081 2692 10137 2694
rect 10161 2692 10217 2694
rect 10241 2692 10297 2694
rect 10494 2760 10550 2816
rect 10678 2644 10734 2680
rect 10678 2624 10680 2644
rect 10680 2624 10732 2644
rect 10732 2624 10734 2644
rect 11046 4664 11102 4720
rect 10310 2216 10366 2272
rect 10494 2080 10550 2136
rect 10402 1400 10458 1456
rect 11598 4140 11654 4176
rect 11598 4120 11600 4140
rect 11600 4120 11652 4140
rect 11652 4120 11654 4140
rect 11138 3712 11194 3768
rect 11874 4020 11876 4040
rect 11876 4020 11928 4040
rect 11928 4020 11930 4040
rect 11874 3984 11930 4020
rect 12426 21972 12428 21992
rect 12428 21972 12480 21992
rect 12480 21972 12482 21992
rect 12426 21936 12482 21972
rect 12334 20984 12390 21040
rect 12886 17060 12942 17096
rect 12886 17040 12888 17060
rect 12888 17040 12940 17060
rect 12940 17040 12942 17060
rect 14668 25050 14724 25052
rect 14748 25050 14804 25052
rect 14828 25050 14884 25052
rect 14908 25050 14964 25052
rect 14668 24998 14694 25050
rect 14694 24998 14724 25050
rect 14748 24998 14758 25050
rect 14758 24998 14804 25050
rect 14828 24998 14874 25050
rect 14874 24998 14884 25050
rect 14908 24998 14938 25050
rect 14938 24998 14964 25050
rect 14668 24996 14724 24998
rect 14748 24996 14804 24998
rect 14828 24996 14884 24998
rect 14908 24996 14964 24998
rect 14668 23962 14724 23964
rect 14748 23962 14804 23964
rect 14828 23962 14884 23964
rect 14908 23962 14964 23964
rect 14668 23910 14694 23962
rect 14694 23910 14724 23962
rect 14748 23910 14758 23962
rect 14758 23910 14804 23962
rect 14828 23910 14874 23962
rect 14874 23910 14884 23962
rect 14908 23910 14938 23962
rect 14938 23910 14964 23962
rect 14668 23908 14724 23910
rect 14748 23908 14804 23910
rect 14828 23908 14884 23910
rect 14908 23908 14964 23910
rect 23558 27104 23614 27160
rect 23466 26560 23522 26616
rect 19334 25594 19390 25596
rect 19414 25594 19470 25596
rect 19494 25594 19550 25596
rect 19574 25594 19630 25596
rect 19334 25542 19360 25594
rect 19360 25542 19390 25594
rect 19414 25542 19424 25594
rect 19424 25542 19470 25594
rect 19494 25542 19540 25594
rect 19540 25542 19550 25594
rect 19574 25542 19604 25594
rect 19604 25542 19630 25594
rect 19334 25540 19390 25542
rect 19414 25540 19470 25542
rect 19494 25540 19550 25542
rect 19574 25540 19630 25542
rect 19334 24506 19390 24508
rect 19414 24506 19470 24508
rect 19494 24506 19550 24508
rect 19574 24506 19630 24508
rect 19334 24454 19360 24506
rect 19360 24454 19390 24506
rect 19414 24454 19424 24506
rect 19424 24454 19470 24506
rect 19494 24454 19540 24506
rect 19540 24454 19550 24506
rect 19574 24454 19604 24506
rect 19604 24454 19630 24506
rect 19334 24452 19390 24454
rect 19414 24452 19470 24454
rect 19494 24452 19550 24454
rect 19574 24452 19630 24454
rect 19334 23418 19390 23420
rect 19414 23418 19470 23420
rect 19494 23418 19550 23420
rect 19574 23418 19630 23420
rect 19334 23366 19360 23418
rect 19360 23366 19390 23418
rect 19414 23366 19424 23418
rect 19424 23366 19470 23418
rect 19494 23366 19540 23418
rect 19540 23366 19550 23418
rect 19574 23366 19604 23418
rect 19604 23366 19630 23418
rect 19334 23364 19390 23366
rect 19414 23364 19470 23366
rect 19494 23364 19550 23366
rect 19574 23364 19630 23366
rect 19234 23160 19290 23216
rect 14668 22874 14724 22876
rect 14748 22874 14804 22876
rect 14828 22874 14884 22876
rect 14908 22874 14964 22876
rect 14668 22822 14694 22874
rect 14694 22822 14724 22874
rect 14748 22822 14758 22874
rect 14758 22822 14804 22874
rect 14828 22822 14874 22874
rect 14874 22822 14884 22874
rect 14908 22822 14938 22874
rect 14938 22822 14964 22874
rect 14668 22820 14724 22822
rect 14748 22820 14804 22822
rect 14828 22820 14884 22822
rect 14908 22820 14964 22822
rect 23190 22500 23246 22536
rect 23190 22480 23192 22500
rect 23192 22480 23244 22500
rect 23244 22480 23246 22500
rect 19334 22330 19390 22332
rect 19414 22330 19470 22332
rect 19494 22330 19550 22332
rect 19574 22330 19630 22332
rect 19334 22278 19360 22330
rect 19360 22278 19390 22330
rect 19414 22278 19424 22330
rect 19424 22278 19470 22330
rect 19494 22278 19540 22330
rect 19540 22278 19550 22330
rect 19574 22278 19604 22330
rect 19604 22278 19630 22330
rect 19334 22276 19390 22278
rect 19414 22276 19470 22278
rect 19494 22276 19550 22278
rect 19574 22276 19630 22278
rect 14668 21786 14724 21788
rect 14748 21786 14804 21788
rect 14828 21786 14884 21788
rect 14908 21786 14964 21788
rect 14668 21734 14694 21786
rect 14694 21734 14724 21786
rect 14748 21734 14758 21786
rect 14758 21734 14804 21786
rect 14828 21734 14874 21786
rect 14874 21734 14884 21786
rect 14908 21734 14938 21786
rect 14938 21734 14964 21786
rect 14668 21732 14724 21734
rect 14748 21732 14804 21734
rect 14828 21732 14884 21734
rect 14908 21732 14964 21734
rect 14726 21428 14728 21448
rect 14728 21428 14780 21448
rect 14780 21428 14782 21448
rect 14726 21392 14782 21428
rect 15002 21412 15058 21448
rect 15002 21392 15004 21412
rect 15004 21392 15056 21412
rect 15056 21392 15058 21412
rect 19334 21242 19390 21244
rect 19414 21242 19470 21244
rect 19494 21242 19550 21244
rect 19574 21242 19630 21244
rect 19334 21190 19360 21242
rect 19360 21190 19390 21242
rect 19414 21190 19424 21242
rect 19424 21190 19470 21242
rect 19494 21190 19540 21242
rect 19540 21190 19550 21242
rect 19574 21190 19604 21242
rect 19604 21190 19630 21242
rect 19334 21188 19390 21190
rect 19414 21188 19470 21190
rect 19494 21188 19550 21190
rect 19574 21188 19630 21190
rect 14668 20698 14724 20700
rect 14748 20698 14804 20700
rect 14828 20698 14884 20700
rect 14908 20698 14964 20700
rect 14668 20646 14694 20698
rect 14694 20646 14724 20698
rect 14748 20646 14758 20698
rect 14758 20646 14804 20698
rect 14828 20646 14874 20698
rect 14874 20646 14884 20698
rect 14908 20646 14938 20698
rect 14938 20646 14964 20698
rect 14668 20644 14724 20646
rect 14748 20644 14804 20646
rect 14828 20644 14884 20646
rect 14908 20644 14964 20646
rect 15646 20304 15702 20360
rect 23190 20340 23192 20360
rect 23192 20340 23244 20360
rect 23244 20340 23246 20360
rect 23190 20304 23246 20340
rect 14668 19610 14724 19612
rect 14748 19610 14804 19612
rect 14828 19610 14884 19612
rect 14908 19610 14964 19612
rect 14668 19558 14694 19610
rect 14694 19558 14724 19610
rect 14748 19558 14758 19610
rect 14758 19558 14804 19610
rect 14828 19558 14874 19610
rect 14874 19558 14884 19610
rect 14908 19558 14938 19610
rect 14938 19558 14964 19610
rect 14668 19556 14724 19558
rect 14748 19556 14804 19558
rect 14828 19556 14884 19558
rect 14908 19556 14964 19558
rect 14668 18522 14724 18524
rect 14748 18522 14804 18524
rect 14828 18522 14884 18524
rect 14908 18522 14964 18524
rect 14668 18470 14694 18522
rect 14694 18470 14724 18522
rect 14748 18470 14758 18522
rect 14758 18470 14804 18522
rect 14828 18470 14874 18522
rect 14874 18470 14884 18522
rect 14908 18470 14938 18522
rect 14938 18470 14964 18522
rect 14668 18468 14724 18470
rect 14748 18468 14804 18470
rect 14828 18468 14884 18470
rect 14908 18468 14964 18470
rect 14668 17434 14724 17436
rect 14748 17434 14804 17436
rect 14828 17434 14884 17436
rect 14908 17434 14964 17436
rect 14668 17382 14694 17434
rect 14694 17382 14724 17434
rect 14748 17382 14758 17434
rect 14758 17382 14804 17434
rect 14828 17382 14874 17434
rect 14874 17382 14884 17434
rect 14908 17382 14938 17434
rect 14938 17382 14964 17434
rect 14668 17380 14724 17382
rect 14748 17380 14804 17382
rect 14828 17380 14884 17382
rect 14908 17380 14964 17382
rect 13530 16496 13586 16552
rect 14668 16346 14724 16348
rect 14748 16346 14804 16348
rect 14828 16346 14884 16348
rect 14908 16346 14964 16348
rect 14668 16294 14694 16346
rect 14694 16294 14724 16346
rect 14748 16294 14758 16346
rect 14758 16294 14804 16346
rect 14828 16294 14874 16346
rect 14874 16294 14884 16346
rect 14908 16294 14938 16346
rect 14938 16294 14964 16346
rect 14668 16292 14724 16294
rect 14748 16292 14804 16294
rect 14828 16292 14884 16294
rect 14908 16292 14964 16294
rect 12426 15816 12482 15872
rect 15002 15852 15004 15872
rect 15004 15852 15056 15872
rect 15056 15852 15058 15872
rect 15002 15816 15058 15852
rect 12334 3712 12390 3768
rect 11874 2916 11930 2952
rect 11874 2896 11876 2916
rect 11876 2896 11928 2916
rect 11928 2896 11930 2916
rect 14668 15258 14724 15260
rect 14748 15258 14804 15260
rect 14828 15258 14884 15260
rect 14908 15258 14964 15260
rect 14668 15206 14694 15258
rect 14694 15206 14724 15258
rect 14748 15206 14758 15258
rect 14758 15206 14804 15258
rect 14828 15206 14874 15258
rect 14874 15206 14884 15258
rect 14908 15206 14938 15258
rect 14938 15206 14964 15258
rect 14668 15204 14724 15206
rect 14748 15204 14804 15206
rect 14828 15204 14884 15206
rect 14908 15204 14964 15206
rect 13162 14864 13218 14920
rect 13070 9288 13126 9344
rect 12610 9016 12666 9072
rect 15186 14456 15242 14512
rect 14668 14170 14724 14172
rect 14748 14170 14804 14172
rect 14828 14170 14884 14172
rect 14908 14170 14964 14172
rect 14668 14118 14694 14170
rect 14694 14118 14724 14170
rect 14748 14118 14758 14170
rect 14758 14118 14804 14170
rect 14828 14118 14874 14170
rect 14874 14118 14884 14170
rect 14908 14118 14938 14170
rect 14938 14118 14964 14170
rect 14668 14116 14724 14118
rect 14748 14116 14804 14118
rect 14828 14116 14884 14118
rect 14908 14116 14964 14118
rect 15002 13232 15058 13288
rect 14668 13082 14724 13084
rect 14748 13082 14804 13084
rect 14828 13082 14884 13084
rect 14908 13082 14964 13084
rect 14668 13030 14694 13082
rect 14694 13030 14724 13082
rect 14748 13030 14758 13082
rect 14758 13030 14804 13082
rect 14828 13030 14874 13082
rect 14874 13030 14884 13082
rect 14908 13030 14938 13082
rect 14938 13030 14964 13082
rect 14668 13028 14724 13030
rect 14748 13028 14804 13030
rect 14828 13028 14884 13030
rect 14908 13028 14964 13030
rect 14668 11994 14724 11996
rect 14748 11994 14804 11996
rect 14828 11994 14884 11996
rect 14908 11994 14964 11996
rect 14668 11942 14694 11994
rect 14694 11942 14724 11994
rect 14748 11942 14758 11994
rect 14758 11942 14804 11994
rect 14828 11942 14874 11994
rect 14874 11942 14884 11994
rect 14908 11942 14938 11994
rect 14938 11942 14964 11994
rect 14668 11940 14724 11942
rect 14748 11940 14804 11942
rect 14828 11940 14884 11942
rect 14908 11940 14964 11942
rect 13622 11600 13678 11656
rect 14450 11328 14506 11384
rect 15002 11328 15058 11384
rect 13346 8356 13402 8392
rect 13346 8336 13348 8356
rect 13348 8336 13400 8356
rect 13400 8336 13402 8356
rect 12794 3848 12850 3904
rect 12886 2916 12942 2952
rect 12886 2896 12888 2916
rect 12888 2896 12940 2916
rect 12940 2896 12942 2916
rect 12610 2624 12666 2680
rect 13622 6604 13624 6624
rect 13624 6604 13676 6624
rect 13676 6604 13678 6624
rect 13622 6568 13678 6604
rect 13346 3440 13402 3496
rect 13070 2624 13126 2680
rect 14358 8064 14414 8120
rect 14358 7792 14414 7848
rect 13898 4936 13954 4992
rect 14668 10906 14724 10908
rect 14748 10906 14804 10908
rect 14828 10906 14884 10908
rect 14908 10906 14964 10908
rect 14668 10854 14694 10906
rect 14694 10854 14724 10906
rect 14748 10854 14758 10906
rect 14758 10854 14804 10906
rect 14828 10854 14874 10906
rect 14874 10854 14884 10906
rect 14908 10854 14938 10906
rect 14938 10854 14964 10906
rect 14668 10852 14724 10854
rect 14748 10852 14804 10854
rect 14828 10852 14884 10854
rect 14908 10852 14964 10854
rect 14668 9818 14724 9820
rect 14748 9818 14804 9820
rect 14828 9818 14884 9820
rect 14908 9818 14964 9820
rect 14668 9766 14694 9818
rect 14694 9766 14724 9818
rect 14748 9766 14758 9818
rect 14758 9766 14804 9818
rect 14828 9766 14874 9818
rect 14874 9766 14884 9818
rect 14908 9766 14938 9818
rect 14938 9766 14964 9818
rect 14668 9764 14724 9766
rect 14748 9764 14804 9766
rect 14828 9764 14884 9766
rect 14908 9764 14964 9766
rect 14668 8730 14724 8732
rect 14748 8730 14804 8732
rect 14828 8730 14884 8732
rect 14908 8730 14964 8732
rect 14668 8678 14694 8730
rect 14694 8678 14724 8730
rect 14748 8678 14758 8730
rect 14758 8678 14804 8730
rect 14828 8678 14874 8730
rect 14874 8678 14884 8730
rect 14908 8678 14938 8730
rect 14938 8678 14964 8730
rect 14668 8676 14724 8678
rect 14748 8676 14804 8678
rect 14828 8676 14884 8678
rect 14908 8676 14964 8678
rect 14668 7642 14724 7644
rect 14748 7642 14804 7644
rect 14828 7642 14884 7644
rect 14908 7642 14964 7644
rect 14668 7590 14694 7642
rect 14694 7590 14724 7642
rect 14748 7590 14758 7642
rect 14758 7590 14804 7642
rect 14828 7590 14874 7642
rect 14874 7590 14884 7642
rect 14908 7590 14938 7642
rect 14938 7590 14964 7642
rect 14668 7588 14724 7590
rect 14748 7588 14804 7590
rect 14828 7588 14884 7590
rect 14908 7588 14964 7590
rect 15278 11212 15334 11248
rect 15278 11192 15280 11212
rect 15280 11192 15332 11212
rect 15332 11192 15334 11212
rect 15370 9036 15426 9072
rect 15370 9016 15372 9036
rect 15372 9016 15424 9036
rect 15424 9016 15426 9036
rect 15370 6840 15426 6896
rect 14668 6554 14724 6556
rect 14748 6554 14804 6556
rect 14828 6554 14884 6556
rect 14908 6554 14964 6556
rect 14668 6502 14694 6554
rect 14694 6502 14724 6554
rect 14748 6502 14758 6554
rect 14758 6502 14804 6554
rect 14828 6502 14874 6554
rect 14874 6502 14884 6554
rect 14908 6502 14938 6554
rect 14938 6502 14964 6554
rect 14668 6500 14724 6502
rect 14748 6500 14804 6502
rect 14828 6500 14884 6502
rect 14908 6500 14964 6502
rect 15554 6432 15610 6488
rect 15002 5772 15058 5808
rect 15002 5752 15004 5772
rect 15004 5752 15056 5772
rect 15056 5752 15058 5772
rect 14668 5466 14724 5468
rect 14748 5466 14804 5468
rect 14828 5466 14884 5468
rect 14908 5466 14964 5468
rect 14668 5414 14694 5466
rect 14694 5414 14724 5466
rect 14748 5414 14758 5466
rect 14758 5414 14804 5466
rect 14828 5414 14874 5466
rect 14874 5414 14884 5466
rect 14908 5414 14938 5466
rect 14938 5414 14964 5466
rect 14668 5412 14724 5414
rect 14748 5412 14804 5414
rect 14828 5412 14884 5414
rect 14908 5412 14964 5414
rect 13622 1400 13678 1456
rect 14358 4800 14414 4856
rect 21442 20168 21498 20224
rect 19334 20154 19390 20156
rect 19414 20154 19470 20156
rect 19494 20154 19550 20156
rect 19574 20154 19630 20156
rect 19334 20102 19360 20154
rect 19360 20102 19390 20154
rect 19414 20102 19424 20154
rect 19424 20102 19470 20154
rect 19494 20102 19540 20154
rect 19540 20102 19550 20154
rect 19574 20102 19604 20154
rect 19604 20102 19630 20154
rect 19334 20100 19390 20102
rect 19414 20100 19470 20102
rect 19494 20100 19550 20102
rect 19574 20100 19630 20102
rect 19334 19066 19390 19068
rect 19414 19066 19470 19068
rect 19494 19066 19550 19068
rect 19574 19066 19630 19068
rect 19334 19014 19360 19066
rect 19360 19014 19390 19066
rect 19414 19014 19424 19066
rect 19424 19014 19470 19066
rect 19494 19014 19540 19066
rect 19540 19014 19550 19066
rect 19574 19014 19604 19066
rect 19604 19014 19630 19066
rect 19334 19012 19390 19014
rect 19414 19012 19470 19014
rect 19494 19012 19550 19014
rect 19574 19012 19630 19014
rect 15738 18828 15794 18864
rect 15738 18808 15740 18828
rect 15740 18808 15792 18828
rect 15792 18808 15794 18828
rect 19334 17978 19390 17980
rect 19414 17978 19470 17980
rect 19494 17978 19550 17980
rect 19574 17978 19630 17980
rect 19334 17926 19360 17978
rect 19360 17926 19390 17978
rect 19414 17926 19424 17978
rect 19424 17926 19470 17978
rect 19494 17926 19540 17978
rect 19540 17926 19550 17978
rect 19574 17926 19604 17978
rect 19604 17926 19630 17978
rect 19334 17924 19390 17926
rect 19414 17924 19470 17926
rect 19494 17924 19550 17926
rect 19574 17924 19630 17926
rect 16014 17604 16070 17640
rect 16014 17584 16016 17604
rect 16016 17584 16068 17604
rect 16068 17584 16070 17604
rect 16106 17312 16162 17368
rect 15922 11756 15978 11792
rect 15922 11736 15924 11756
rect 15924 11736 15976 11756
rect 15976 11736 15978 11756
rect 15738 10104 15794 10160
rect 14358 4392 14414 4448
rect 14668 4378 14724 4380
rect 14748 4378 14804 4380
rect 14828 4378 14884 4380
rect 14908 4378 14964 4380
rect 14668 4326 14694 4378
rect 14694 4326 14724 4378
rect 14748 4326 14758 4378
rect 14758 4326 14804 4378
rect 14828 4326 14874 4378
rect 14874 4326 14884 4378
rect 14908 4326 14938 4378
rect 14938 4326 14964 4378
rect 14668 4324 14724 4326
rect 14748 4324 14804 4326
rect 14828 4324 14884 4326
rect 14908 4324 14964 4326
rect 15278 4392 15334 4448
rect 15370 3596 15426 3632
rect 15370 3576 15372 3596
rect 15372 3576 15424 3596
rect 15424 3576 15426 3596
rect 14542 3440 14598 3496
rect 14668 3290 14724 3292
rect 14748 3290 14804 3292
rect 14828 3290 14884 3292
rect 14908 3290 14964 3292
rect 14668 3238 14694 3290
rect 14694 3238 14724 3290
rect 14748 3238 14758 3290
rect 14758 3238 14804 3290
rect 14828 3238 14874 3290
rect 14874 3238 14884 3290
rect 14908 3238 14938 3290
rect 14938 3238 14964 3290
rect 14668 3236 14724 3238
rect 14748 3236 14804 3238
rect 14828 3236 14884 3238
rect 14908 3236 14964 3238
rect 15002 2896 15058 2952
rect 14668 2202 14724 2204
rect 14748 2202 14804 2204
rect 14828 2202 14884 2204
rect 14908 2202 14964 2204
rect 14668 2150 14694 2202
rect 14694 2150 14724 2202
rect 14748 2150 14758 2202
rect 14758 2150 14804 2202
rect 14828 2150 14874 2202
rect 14874 2150 14884 2202
rect 14908 2150 14938 2202
rect 14938 2150 14964 2202
rect 14668 2148 14724 2150
rect 14748 2148 14804 2150
rect 14828 2148 14884 2150
rect 14908 2148 14964 2150
rect 15922 6296 15978 6352
rect 15830 6196 15832 6216
rect 15832 6196 15884 6216
rect 15884 6196 15886 6216
rect 15830 6160 15886 6196
rect 19334 16890 19390 16892
rect 19414 16890 19470 16892
rect 19494 16890 19550 16892
rect 19574 16890 19630 16892
rect 19334 16838 19360 16890
rect 19360 16838 19390 16890
rect 19414 16838 19424 16890
rect 19424 16838 19470 16890
rect 19494 16838 19540 16890
rect 19540 16838 19550 16890
rect 19574 16838 19604 16890
rect 19604 16838 19630 16890
rect 19334 16836 19390 16838
rect 19414 16836 19470 16838
rect 19494 16836 19550 16838
rect 19574 16836 19630 16838
rect 18222 16632 18278 16688
rect 18590 13932 18646 13968
rect 18590 13912 18592 13932
rect 18592 13912 18644 13932
rect 18644 13912 18646 13932
rect 16658 12824 16714 12880
rect 16198 11056 16254 11112
rect 18590 12708 18646 12744
rect 18590 12688 18592 12708
rect 18592 12688 18644 12708
rect 18644 12688 18646 12708
rect 16842 10920 16898 10976
rect 16474 7384 16530 7440
rect 16198 5480 16254 5536
rect 16106 4800 16162 4856
rect 16382 5072 16438 5128
rect 16290 4256 16346 4312
rect 16382 3188 16438 3224
rect 16382 3168 16384 3188
rect 16384 3168 16436 3188
rect 16436 3168 16438 3188
rect 18314 11076 18370 11112
rect 18314 11056 18316 11076
rect 18316 11056 18368 11076
rect 18368 11056 18370 11076
rect 17486 9444 17542 9480
rect 17486 9424 17488 9444
rect 17488 9424 17540 9444
rect 17540 9424 17542 9444
rect 17854 9560 17910 9616
rect 17854 9424 17910 9480
rect 17946 8744 18002 8800
rect 17854 8064 17910 8120
rect 17118 6704 17174 6760
rect 17026 5208 17082 5264
rect 16934 5072 16990 5128
rect 16842 4936 16898 4992
rect 16934 4120 16990 4176
rect 17302 6704 17358 6760
rect 17302 5364 17358 5400
rect 17302 5344 17304 5364
rect 17304 5344 17356 5364
rect 17356 5344 17358 5364
rect 17210 4392 17266 4448
rect 17118 3712 17174 3768
rect 16750 2896 16806 2952
rect 16566 2644 16622 2680
rect 16566 2624 16568 2644
rect 16568 2624 16620 2644
rect 16620 2624 16622 2644
rect 18222 7656 18278 7712
rect 18314 7404 18370 7440
rect 18314 7384 18316 7404
rect 18316 7384 18368 7404
rect 18368 7384 18370 7404
rect 18498 7248 18554 7304
rect 18038 5208 18094 5264
rect 17946 4256 18002 4312
rect 19334 15802 19390 15804
rect 19414 15802 19470 15804
rect 19494 15802 19550 15804
rect 19574 15802 19630 15804
rect 19334 15750 19360 15802
rect 19360 15750 19390 15802
rect 19414 15750 19424 15802
rect 19424 15750 19470 15802
rect 19494 15750 19540 15802
rect 19540 15750 19550 15802
rect 19574 15750 19604 15802
rect 19604 15750 19630 15802
rect 19334 15748 19390 15750
rect 19414 15748 19470 15750
rect 19494 15748 19550 15750
rect 19574 15748 19630 15750
rect 19334 14714 19390 14716
rect 19414 14714 19470 14716
rect 19494 14714 19550 14716
rect 19574 14714 19630 14716
rect 19334 14662 19360 14714
rect 19360 14662 19390 14714
rect 19414 14662 19424 14714
rect 19424 14662 19470 14714
rect 19494 14662 19540 14714
rect 19540 14662 19550 14714
rect 19574 14662 19604 14714
rect 19604 14662 19630 14714
rect 19334 14660 19390 14662
rect 19414 14660 19470 14662
rect 19494 14660 19550 14662
rect 19574 14660 19630 14662
rect 19334 13626 19390 13628
rect 19414 13626 19470 13628
rect 19494 13626 19550 13628
rect 19574 13626 19630 13628
rect 19334 13574 19360 13626
rect 19360 13574 19390 13626
rect 19414 13574 19424 13626
rect 19424 13574 19470 13626
rect 19494 13574 19540 13626
rect 19540 13574 19550 13626
rect 19574 13574 19604 13626
rect 19604 13574 19630 13626
rect 19334 13572 19390 13574
rect 19414 13572 19470 13574
rect 19494 13572 19550 13574
rect 19574 13572 19630 13574
rect 18958 13096 19014 13152
rect 18958 12688 19014 12744
rect 19334 12538 19390 12540
rect 19414 12538 19470 12540
rect 19494 12538 19550 12540
rect 19574 12538 19630 12540
rect 19334 12486 19360 12538
rect 19360 12486 19390 12538
rect 19414 12486 19424 12538
rect 19424 12486 19470 12538
rect 19494 12486 19540 12538
rect 19540 12486 19550 12538
rect 19574 12486 19604 12538
rect 19604 12486 19630 12538
rect 19334 12484 19390 12486
rect 19414 12484 19470 12486
rect 19494 12484 19550 12486
rect 19574 12484 19630 12486
rect 19334 11450 19390 11452
rect 19414 11450 19470 11452
rect 19494 11450 19550 11452
rect 19574 11450 19630 11452
rect 19334 11398 19360 11450
rect 19360 11398 19390 11450
rect 19414 11398 19424 11450
rect 19424 11398 19470 11450
rect 19494 11398 19540 11450
rect 19540 11398 19550 11450
rect 19574 11398 19604 11450
rect 19604 11398 19630 11450
rect 19334 11396 19390 11398
rect 19414 11396 19470 11398
rect 19494 11396 19550 11398
rect 19574 11396 19630 11398
rect 19334 10362 19390 10364
rect 19414 10362 19470 10364
rect 19494 10362 19550 10364
rect 19574 10362 19630 10364
rect 19334 10310 19360 10362
rect 19360 10310 19390 10362
rect 19414 10310 19424 10362
rect 19424 10310 19470 10362
rect 19494 10310 19540 10362
rect 19540 10310 19550 10362
rect 19574 10310 19604 10362
rect 19604 10310 19630 10362
rect 19334 10308 19390 10310
rect 19414 10308 19470 10310
rect 19494 10308 19550 10310
rect 19574 10308 19630 10310
rect 18866 9324 18868 9344
rect 18868 9324 18920 9344
rect 18920 9324 18922 9344
rect 18866 9288 18922 9324
rect 22454 17312 22510 17368
rect 21534 16496 21590 16552
rect 20522 13132 20524 13152
rect 20524 13132 20576 13152
rect 20576 13132 20578 13152
rect 20522 13096 20578 13132
rect 21074 12960 21130 13016
rect 20614 11600 20670 11656
rect 19334 9274 19390 9276
rect 19414 9274 19470 9276
rect 19494 9274 19550 9276
rect 19574 9274 19630 9276
rect 19334 9222 19360 9274
rect 19360 9222 19390 9274
rect 19414 9222 19424 9274
rect 19424 9222 19470 9274
rect 19494 9222 19540 9274
rect 19540 9222 19550 9274
rect 19574 9222 19604 9274
rect 19604 9222 19630 9274
rect 19334 9220 19390 9222
rect 19414 9220 19470 9222
rect 19494 9220 19550 9222
rect 19574 9220 19630 9222
rect 18958 8336 19014 8392
rect 19334 8186 19390 8188
rect 19414 8186 19470 8188
rect 19494 8186 19550 8188
rect 19574 8186 19630 8188
rect 19334 8134 19360 8186
rect 19360 8134 19390 8186
rect 19414 8134 19424 8186
rect 19424 8134 19470 8186
rect 19494 8134 19540 8186
rect 19540 8134 19550 8186
rect 19574 8134 19604 8186
rect 19604 8134 19630 8186
rect 19334 8132 19390 8134
rect 19414 8132 19470 8134
rect 19494 8132 19550 8134
rect 19574 8132 19630 8134
rect 18958 7792 19014 7848
rect 18774 6296 18830 6352
rect 17486 3032 17542 3088
rect 18130 4004 18186 4040
rect 18130 3984 18132 4004
rect 18132 3984 18184 4004
rect 18184 3984 18186 4004
rect 19334 7098 19390 7100
rect 19414 7098 19470 7100
rect 19494 7098 19550 7100
rect 19574 7098 19630 7100
rect 19334 7046 19360 7098
rect 19360 7046 19390 7098
rect 19414 7046 19424 7098
rect 19424 7046 19470 7098
rect 19494 7046 19540 7098
rect 19540 7046 19550 7098
rect 19574 7046 19604 7098
rect 19604 7046 19630 7098
rect 19334 7044 19390 7046
rect 19414 7044 19470 7046
rect 19494 7044 19550 7046
rect 19574 7044 19630 7046
rect 19334 6010 19390 6012
rect 19414 6010 19470 6012
rect 19494 6010 19550 6012
rect 19574 6010 19630 6012
rect 19334 5958 19360 6010
rect 19360 5958 19390 6010
rect 19414 5958 19424 6010
rect 19424 5958 19470 6010
rect 19494 5958 19540 6010
rect 19540 5958 19550 6010
rect 19574 5958 19604 6010
rect 19604 5958 19630 6010
rect 19334 5956 19390 5958
rect 19414 5956 19470 5958
rect 19494 5956 19550 5958
rect 19574 5956 19630 5958
rect 20614 8916 20616 8936
rect 20616 8916 20668 8936
rect 20668 8916 20670 8936
rect 20614 8880 20670 8916
rect 19786 7112 19842 7168
rect 19510 5616 19566 5672
rect 19694 5616 19750 5672
rect 19142 5480 19198 5536
rect 18866 4256 18922 4312
rect 18314 2508 18370 2544
rect 18314 2488 18316 2508
rect 18316 2488 18368 2508
rect 18368 2488 18370 2508
rect 18682 3476 18684 3496
rect 18684 3476 18736 3496
rect 18736 3476 18738 3496
rect 18682 3440 18738 3476
rect 19334 4922 19390 4924
rect 19414 4922 19470 4924
rect 19494 4922 19550 4924
rect 19574 4922 19630 4924
rect 19334 4870 19360 4922
rect 19360 4870 19390 4922
rect 19414 4870 19424 4922
rect 19424 4870 19470 4922
rect 19494 4870 19540 4922
rect 19540 4870 19550 4922
rect 19574 4870 19604 4922
rect 19604 4870 19630 4922
rect 19334 4868 19390 4870
rect 19414 4868 19470 4870
rect 19494 4868 19550 4870
rect 19574 4868 19630 4870
rect 20982 8356 21038 8392
rect 20982 8336 20984 8356
rect 20984 8336 21036 8356
rect 21036 8336 21038 8356
rect 19970 7404 20026 7440
rect 19970 7384 19972 7404
rect 19972 7384 20024 7404
rect 20024 7384 20026 7404
rect 19970 4800 20026 4856
rect 23098 14864 23154 14920
rect 21718 11736 21774 11792
rect 23190 13776 23246 13832
rect 24478 25336 24534 25392
rect 24001 25050 24057 25052
rect 24081 25050 24137 25052
rect 24161 25050 24217 25052
rect 24241 25050 24297 25052
rect 24001 24998 24027 25050
rect 24027 24998 24057 25050
rect 24081 24998 24091 25050
rect 24091 24998 24137 25050
rect 24161 24998 24207 25050
rect 24207 24998 24217 25050
rect 24241 24998 24271 25050
rect 24271 24998 24297 25050
rect 24001 24996 24057 24998
rect 24081 24996 24137 24998
rect 24161 24996 24217 24998
rect 24241 24996 24297 24998
rect 24386 24248 24442 24304
rect 24001 23962 24057 23964
rect 24081 23962 24137 23964
rect 24161 23962 24217 23964
rect 24241 23962 24297 23964
rect 24001 23910 24027 23962
rect 24027 23910 24057 23962
rect 24081 23910 24091 23962
rect 24091 23910 24137 23962
rect 24161 23910 24207 23962
rect 24207 23910 24217 23962
rect 24241 23910 24271 23962
rect 24271 23910 24297 23962
rect 24001 23908 24057 23910
rect 24081 23908 24137 23910
rect 24161 23908 24217 23910
rect 24241 23908 24297 23910
rect 23742 23704 23798 23760
rect 24001 22874 24057 22876
rect 24081 22874 24137 22876
rect 24161 22874 24217 22876
rect 24241 22874 24297 22876
rect 24001 22822 24027 22874
rect 24027 22822 24057 22874
rect 24081 22822 24091 22874
rect 24091 22822 24137 22874
rect 24161 22822 24207 22874
rect 24207 22822 24217 22874
rect 24241 22822 24271 22874
rect 24271 22822 24297 22874
rect 24001 22820 24057 22822
rect 24081 22820 24137 22822
rect 24161 22820 24217 22822
rect 24241 22820 24297 22822
rect 25122 26016 25178 26072
rect 24478 23160 24534 23216
rect 24478 22616 24534 22672
rect 24386 22380 24388 22400
rect 24388 22380 24440 22400
rect 24440 22380 24442 22400
rect 24386 22344 24442 22380
rect 24001 21786 24057 21788
rect 24081 21786 24137 21788
rect 24161 21786 24217 21788
rect 24241 21786 24297 21788
rect 24001 21734 24027 21786
rect 24027 21734 24057 21786
rect 24081 21734 24091 21786
rect 24091 21734 24137 21786
rect 24161 21734 24207 21786
rect 24207 21734 24217 21786
rect 24241 21734 24271 21786
rect 24271 21734 24297 21786
rect 24001 21732 24057 21734
rect 24081 21732 24137 21734
rect 24161 21732 24217 21734
rect 24241 21732 24297 21734
rect 23558 21528 23614 21584
rect 24754 22480 24810 22536
rect 24662 21936 24718 21992
rect 24110 21428 24112 21448
rect 24112 21428 24164 21448
rect 24164 21428 24166 21448
rect 24110 21392 24166 21428
rect 24386 21392 24442 21448
rect 24001 20698 24057 20700
rect 24081 20698 24137 20700
rect 24161 20698 24217 20700
rect 24241 20698 24297 20700
rect 24001 20646 24027 20698
rect 24027 20646 24057 20698
rect 24081 20646 24091 20698
rect 24091 20646 24137 20698
rect 24161 20646 24207 20698
rect 24207 20646 24217 20698
rect 24241 20646 24271 20698
rect 24271 20646 24297 20698
rect 24001 20644 24057 20646
rect 24081 20644 24137 20646
rect 24161 20644 24217 20646
rect 24241 20644 24297 20646
rect 24478 20848 24534 20904
rect 24001 19610 24057 19612
rect 24081 19610 24137 19612
rect 24161 19610 24217 19612
rect 24241 19610 24297 19612
rect 24001 19558 24027 19610
rect 24027 19558 24057 19610
rect 24081 19558 24091 19610
rect 24091 19558 24137 19610
rect 24161 19558 24207 19610
rect 24207 19558 24217 19610
rect 24241 19558 24271 19610
rect 24271 19558 24297 19610
rect 24001 19556 24057 19558
rect 24081 19556 24137 19558
rect 24161 19556 24217 19558
rect 24241 19556 24297 19558
rect 23834 19352 23890 19408
rect 23834 19080 23890 19136
rect 23834 17584 23890 17640
rect 23834 17176 23890 17232
rect 23742 15000 23798 15056
rect 22730 12416 22786 12472
rect 22822 12280 22878 12336
rect 23006 12416 23062 12472
rect 23374 12724 23376 12744
rect 23376 12724 23428 12744
rect 23428 12724 23430 12744
rect 23374 12688 23430 12724
rect 22362 11056 22418 11112
rect 22822 11056 22878 11112
rect 20890 6452 20946 6488
rect 20890 6432 20892 6452
rect 20892 6432 20944 6452
rect 20944 6432 20946 6452
rect 20154 4392 20210 4448
rect 19878 4120 19934 4176
rect 20062 3884 20064 3904
rect 20064 3884 20116 3904
rect 20116 3884 20118 3904
rect 19334 3834 19390 3836
rect 19414 3834 19470 3836
rect 19494 3834 19550 3836
rect 19574 3834 19630 3836
rect 19334 3782 19360 3834
rect 19360 3782 19390 3834
rect 19414 3782 19424 3834
rect 19424 3782 19470 3834
rect 19494 3782 19540 3834
rect 19540 3782 19550 3834
rect 19574 3782 19604 3834
rect 19604 3782 19630 3834
rect 19334 3780 19390 3782
rect 19414 3780 19470 3782
rect 19494 3780 19550 3782
rect 19574 3780 19630 3782
rect 19694 3576 19750 3632
rect 19234 3168 19290 3224
rect 19142 2760 19198 2816
rect 19334 2746 19390 2748
rect 19414 2746 19470 2748
rect 19494 2746 19550 2748
rect 19574 2746 19630 2748
rect 19334 2694 19360 2746
rect 19360 2694 19390 2746
rect 19414 2694 19424 2746
rect 19424 2694 19470 2746
rect 19494 2694 19540 2746
rect 19540 2694 19550 2746
rect 19574 2694 19604 2746
rect 19604 2694 19630 2746
rect 19334 2692 19390 2694
rect 19414 2692 19470 2694
rect 19494 2692 19550 2694
rect 19574 2692 19630 2694
rect 20062 3848 20118 3884
rect 19970 3340 19972 3360
rect 19972 3340 20024 3360
rect 20024 3340 20026 3360
rect 19970 3304 20026 3340
rect 20614 3984 20670 4040
rect 21534 7148 21536 7168
rect 21536 7148 21588 7168
rect 21588 7148 21590 7168
rect 21534 7112 21590 7148
rect 21994 7384 22050 7440
rect 21626 6840 21682 6896
rect 21534 6568 21590 6624
rect 21442 4120 21498 4176
rect 20890 3440 20946 3496
rect 20706 3032 20762 3088
rect 20798 2624 20854 2680
rect 20154 1808 20210 1864
rect 20246 1536 20302 1592
rect 21534 3712 21590 3768
rect 21718 6452 21774 6488
rect 21718 6432 21720 6452
rect 21720 6432 21772 6452
rect 21772 6432 21774 6452
rect 22362 6296 22418 6352
rect 22178 5888 22234 5944
rect 22086 4820 22142 4856
rect 22086 4800 22088 4820
rect 22088 4800 22140 4820
rect 22140 4800 22142 4820
rect 21994 4684 22050 4720
rect 21994 4664 21996 4684
rect 21996 4664 22048 4684
rect 22048 4664 22050 4684
rect 22546 5652 22548 5672
rect 22548 5652 22600 5672
rect 22600 5652 22602 5672
rect 22546 5616 22602 5652
rect 22730 5208 22786 5264
rect 21718 2508 21774 2544
rect 21718 2488 21720 2508
rect 21720 2488 21772 2508
rect 21772 2488 21774 2508
rect 21902 2488 21958 2544
rect 23190 9580 23246 9616
rect 23190 9560 23192 9580
rect 23192 9560 23244 9580
rect 23244 9560 23246 9580
rect 23466 8744 23522 8800
rect 23098 7948 23154 7984
rect 23098 7928 23100 7948
rect 23100 7928 23152 7948
rect 23152 7928 23154 7948
rect 23374 5752 23430 5808
rect 23282 5344 23338 5400
rect 23190 4256 23246 4312
rect 23742 12960 23798 13016
rect 24570 20204 24572 20224
rect 24572 20204 24624 20224
rect 24624 20204 24626 20224
rect 24570 20168 24626 20204
rect 24846 19624 24902 19680
rect 24110 18808 24166 18864
rect 24386 18536 24442 18592
rect 24001 18522 24057 18524
rect 24081 18522 24137 18524
rect 24161 18522 24217 18524
rect 24241 18522 24297 18524
rect 24001 18470 24027 18522
rect 24027 18470 24057 18522
rect 24081 18470 24091 18522
rect 24091 18470 24137 18522
rect 24161 18470 24207 18522
rect 24207 18470 24217 18522
rect 24241 18470 24271 18522
rect 24271 18470 24297 18522
rect 24001 18468 24057 18470
rect 24081 18468 24137 18470
rect 24161 18468 24217 18470
rect 24241 18468 24297 18470
rect 24001 17434 24057 17436
rect 24081 17434 24137 17436
rect 24161 17434 24217 17436
rect 24241 17434 24297 17436
rect 24001 17382 24027 17434
rect 24027 17382 24057 17434
rect 24081 17382 24091 17434
rect 24091 17382 24137 17434
rect 24161 17382 24207 17434
rect 24207 17382 24217 17434
rect 24241 17382 24271 17434
rect 24271 17382 24297 17434
rect 24001 17380 24057 17382
rect 24081 17380 24137 17382
rect 24161 17380 24217 17382
rect 24241 17380 24297 17382
rect 24478 17992 24534 18048
rect 24662 17040 24718 17096
rect 24294 16632 24350 16688
rect 24478 16632 24534 16688
rect 24001 16346 24057 16348
rect 24081 16346 24137 16348
rect 24161 16346 24217 16348
rect 24241 16346 24297 16348
rect 24001 16294 24027 16346
rect 24027 16294 24057 16346
rect 24081 16294 24091 16346
rect 24091 16294 24137 16346
rect 24161 16294 24207 16346
rect 24207 16294 24217 16346
rect 24241 16294 24271 16346
rect 24271 16294 24297 16346
rect 24001 16292 24057 16294
rect 24081 16292 24137 16294
rect 24161 16292 24217 16294
rect 24241 16292 24297 16294
rect 24386 15680 24442 15736
rect 24001 15258 24057 15260
rect 24081 15258 24137 15260
rect 24161 15258 24217 15260
rect 24241 15258 24297 15260
rect 24001 15206 24027 15258
rect 24027 15206 24057 15258
rect 24081 15206 24091 15258
rect 24091 15206 24137 15258
rect 24161 15206 24207 15258
rect 24207 15206 24217 15258
rect 24241 15206 24271 15258
rect 24271 15206 24297 15258
rect 24001 15204 24057 15206
rect 24081 15204 24137 15206
rect 24161 15204 24217 15206
rect 24241 15204 24297 15206
rect 24662 16224 24718 16280
rect 24001 14170 24057 14172
rect 24081 14170 24137 14172
rect 24161 14170 24217 14172
rect 24241 14170 24297 14172
rect 24001 14118 24027 14170
rect 24027 14118 24057 14170
rect 24081 14118 24091 14170
rect 24091 14118 24137 14170
rect 24161 14118 24207 14170
rect 24207 14118 24217 14170
rect 24241 14118 24271 14170
rect 24271 14118 24297 14170
rect 24001 14116 24057 14118
rect 24081 14116 24137 14118
rect 24161 14116 24217 14118
rect 24241 14116 24297 14118
rect 24386 13912 24442 13968
rect 24846 13948 24848 13968
rect 24848 13948 24900 13968
rect 24900 13948 24902 13968
rect 24846 13912 24902 13948
rect 24001 13082 24057 13084
rect 24081 13082 24137 13084
rect 24161 13082 24217 13084
rect 24241 13082 24297 13084
rect 24001 13030 24027 13082
rect 24027 13030 24057 13082
rect 24081 13030 24091 13082
rect 24091 13030 24137 13082
rect 24161 13030 24207 13082
rect 24207 13030 24217 13082
rect 24241 13030 24271 13082
rect 24271 13030 24297 13082
rect 24001 13028 24057 13030
rect 24081 13028 24137 13030
rect 24161 13028 24217 13030
rect 24241 13028 24297 13030
rect 24294 12860 24296 12880
rect 24296 12860 24348 12880
rect 24348 12860 24350 12880
rect 24846 13232 24902 13288
rect 24294 12824 24350 12860
rect 24478 12824 24534 12880
rect 24001 11994 24057 11996
rect 24081 11994 24137 11996
rect 24161 11994 24217 11996
rect 24241 11994 24297 11996
rect 24001 11942 24027 11994
rect 24027 11942 24057 11994
rect 24081 11942 24091 11994
rect 24091 11942 24137 11994
rect 24161 11942 24207 11994
rect 24207 11942 24217 11994
rect 24241 11942 24271 11994
rect 24271 11942 24297 11994
rect 24001 11940 24057 11942
rect 24081 11940 24137 11942
rect 24161 11940 24217 11942
rect 24241 11940 24297 11942
rect 25950 22344 26006 22400
rect 25306 14592 25362 14648
rect 25398 13368 25454 13424
rect 24478 11736 24534 11792
rect 24001 10906 24057 10908
rect 24081 10906 24137 10908
rect 24161 10906 24217 10908
rect 24241 10906 24297 10908
rect 24001 10854 24027 10906
rect 24027 10854 24057 10906
rect 24081 10854 24091 10906
rect 24091 10854 24137 10906
rect 24161 10854 24207 10906
rect 24207 10854 24217 10906
rect 24241 10854 24271 10906
rect 24271 10854 24297 10906
rect 24001 10852 24057 10854
rect 24081 10852 24137 10854
rect 24161 10852 24217 10854
rect 24241 10852 24297 10854
rect 23834 10512 23890 10568
rect 23650 8200 23706 8256
rect 24386 9968 24442 10024
rect 24938 11192 24994 11248
rect 24001 9818 24057 9820
rect 24081 9818 24137 9820
rect 24161 9818 24217 9820
rect 24241 9818 24297 9820
rect 24001 9766 24027 9818
rect 24027 9766 24057 9818
rect 24081 9766 24091 9818
rect 24091 9766 24137 9818
rect 24161 9766 24207 9818
rect 24207 9766 24217 9818
rect 24241 9766 24271 9818
rect 24271 9766 24297 9818
rect 24001 9764 24057 9766
rect 24081 9764 24137 9766
rect 24161 9764 24217 9766
rect 24241 9764 24297 9766
rect 24001 8730 24057 8732
rect 24081 8730 24137 8732
rect 24161 8730 24217 8732
rect 24241 8730 24297 8732
rect 24001 8678 24027 8730
rect 24027 8678 24057 8730
rect 24081 8678 24091 8730
rect 24091 8678 24137 8730
rect 24161 8678 24207 8730
rect 24207 8678 24217 8730
rect 24241 8678 24271 8730
rect 24271 8678 24297 8730
rect 24001 8676 24057 8678
rect 24081 8676 24137 8678
rect 24161 8676 24217 8678
rect 24241 8676 24297 8678
rect 23190 3848 23246 3904
rect 24001 7642 24057 7644
rect 24081 7642 24137 7644
rect 24161 7642 24217 7644
rect 24241 7642 24297 7644
rect 24001 7590 24027 7642
rect 24027 7590 24057 7642
rect 24081 7590 24091 7642
rect 24091 7590 24137 7642
rect 24161 7590 24207 7642
rect 24207 7590 24217 7642
rect 24241 7590 24271 7642
rect 24271 7590 24297 7642
rect 24001 7588 24057 7590
rect 24081 7588 24137 7590
rect 24161 7588 24217 7590
rect 24241 7588 24297 7590
rect 23834 6432 23890 6488
rect 23834 5888 23890 5944
rect 23742 4936 23798 4992
rect 24001 6554 24057 6556
rect 24081 6554 24137 6556
rect 24161 6554 24217 6556
rect 24241 6554 24297 6556
rect 24001 6502 24027 6554
rect 24027 6502 24057 6554
rect 24081 6502 24091 6554
rect 24091 6502 24137 6554
rect 24161 6502 24207 6554
rect 24207 6502 24217 6554
rect 24241 6502 24271 6554
rect 24271 6502 24297 6554
rect 24001 6500 24057 6502
rect 24081 6500 24137 6502
rect 24161 6500 24217 6502
rect 24241 6500 24297 6502
rect 24001 5466 24057 5468
rect 24081 5466 24137 5468
rect 24161 5466 24217 5468
rect 24241 5466 24297 5468
rect 24001 5414 24027 5466
rect 24027 5414 24057 5466
rect 24081 5414 24091 5466
rect 24091 5414 24137 5466
rect 24161 5414 24207 5466
rect 24207 5414 24217 5466
rect 24241 5414 24271 5466
rect 24271 5414 24297 5466
rect 24001 5412 24057 5414
rect 24081 5412 24137 5414
rect 24161 5412 24217 5414
rect 24241 5412 24297 5414
rect 24478 8880 24534 8936
rect 24938 10104 24994 10160
rect 24386 4800 24442 4856
rect 24938 7812 24994 7848
rect 24938 7792 24940 7812
rect 24940 7792 24992 7812
rect 24992 7792 24994 7812
rect 25674 7656 25730 7712
rect 24754 4936 24810 4992
rect 24001 4378 24057 4380
rect 24081 4378 24137 4380
rect 24161 4378 24217 4380
rect 24241 4378 24297 4380
rect 24001 4326 24027 4378
rect 24027 4326 24057 4378
rect 24081 4326 24091 4378
rect 24091 4326 24137 4378
rect 24161 4326 24207 4378
rect 24207 4326 24217 4378
rect 24241 4326 24271 4378
rect 24271 4326 24297 4378
rect 24001 4324 24057 4326
rect 24081 4324 24137 4326
rect 24161 4324 24217 4326
rect 24241 4324 24297 4326
rect 24386 4256 24442 4312
rect 23466 3304 23522 3360
rect 23374 2896 23430 2952
rect 24001 3290 24057 3292
rect 24081 3290 24137 3292
rect 24161 3290 24217 3292
rect 24241 3290 24297 3292
rect 24001 3238 24027 3290
rect 24027 3238 24057 3290
rect 24081 3238 24091 3290
rect 24091 3238 24137 3290
rect 24161 3238 24207 3290
rect 24207 3238 24217 3290
rect 24241 3238 24271 3290
rect 24271 3238 24297 3290
rect 24001 3236 24057 3238
rect 24081 3236 24137 3238
rect 24161 3236 24217 3238
rect 24241 3236 24297 3238
rect 23926 3052 23982 3088
rect 23926 3032 23928 3052
rect 23928 3032 23980 3052
rect 23980 3032 23982 3052
rect 23650 1808 23706 1864
rect 23466 1400 23522 1456
rect 24202 2644 24258 2680
rect 24202 2624 24204 2644
rect 24204 2624 24256 2644
rect 24256 2624 24258 2644
rect 24110 2352 24166 2408
rect 24001 2202 24057 2204
rect 24081 2202 24137 2204
rect 24161 2202 24217 2204
rect 24241 2202 24297 2204
rect 24001 2150 24027 2202
rect 24027 2150 24057 2202
rect 24081 2150 24091 2202
rect 24091 2150 24137 2202
rect 24161 2150 24207 2202
rect 24207 2150 24217 2202
rect 24241 2150 24271 2202
rect 24271 2150 24297 2202
rect 24001 2148 24057 2150
rect 24081 2148 24137 2150
rect 24161 2148 24217 2150
rect 24241 2148 24297 2150
rect 24846 3440 24902 3496
rect 25030 3168 25086 3224
rect 24662 2896 24718 2952
rect 24570 1672 24626 1728
rect 24478 856 24534 912
rect 25122 2796 25124 2816
rect 25124 2796 25176 2816
rect 25176 2796 25178 2816
rect 25122 2760 25178 2796
rect 25306 3576 25362 3632
rect 25306 1944 25362 2000
rect 27238 2760 27294 2816
rect 23834 312 23890 368
<< metal3 >>
rect 23686 27644 23692 27708
rect 23756 27706 23762 27708
rect 27232 27706 27712 27736
rect 23756 27646 27712 27706
rect 23756 27644 23762 27646
rect 27232 27616 27712 27646
rect 23553 27162 23619 27165
rect 27232 27162 27712 27192
rect 23553 27160 27712 27162
rect 23553 27104 23558 27160
rect 23614 27104 27712 27160
rect 23553 27102 27712 27104
rect 23553 27099 23619 27102
rect 27232 27072 27712 27102
rect 23461 26618 23527 26621
rect 27232 26618 27712 26648
rect 23461 26616 27712 26618
rect 23461 26560 23466 26616
rect 23522 26560 27712 26616
rect 23461 26558 27712 26560
rect 23461 26555 23527 26558
rect 27232 26528 27712 26558
rect 25117 26074 25183 26077
rect 27232 26074 27712 26104
rect 25117 26072 27712 26074
rect 25117 26016 25122 26072
rect 25178 26016 27712 26072
rect 25117 26014 27712 26016
rect 25117 26011 25183 26014
rect 27232 25984 27712 26014
rect 9989 25600 10309 25601
rect 9989 25536 9997 25600
rect 10061 25536 10077 25600
rect 10141 25536 10157 25600
rect 10221 25536 10237 25600
rect 10301 25536 10309 25600
rect 9989 25535 10309 25536
rect 19322 25600 19642 25601
rect 19322 25536 19330 25600
rect 19394 25536 19410 25600
rect 19474 25536 19490 25600
rect 19554 25536 19570 25600
rect 19634 25536 19642 25600
rect 19322 25535 19642 25536
rect 24473 25394 24539 25397
rect 27232 25394 27712 25424
rect 24473 25392 27712 25394
rect 24473 25336 24478 25392
rect 24534 25336 27712 25392
rect 24473 25334 27712 25336
rect 24473 25331 24539 25334
rect 27232 25304 27712 25334
rect 5322 25056 5642 25057
rect 5322 24992 5330 25056
rect 5394 24992 5410 25056
rect 5474 24992 5490 25056
rect 5554 24992 5570 25056
rect 5634 24992 5642 25056
rect 5322 24991 5642 24992
rect 14656 25056 14976 25057
rect 14656 24992 14664 25056
rect 14728 24992 14744 25056
rect 14808 24992 14824 25056
rect 14888 24992 14904 25056
rect 14968 24992 14976 25056
rect 14656 24991 14976 24992
rect 23989 25056 24309 25057
rect 23989 24992 23997 25056
rect 24061 24992 24077 25056
rect 24141 24992 24157 25056
rect 24221 24992 24237 25056
rect 24301 24992 24309 25056
rect 23989 24991 24309 24992
rect 27232 24850 27712 24880
rect 27190 24760 27712 24850
rect 27190 24578 27250 24760
rect 26638 24518 27250 24578
rect 9989 24512 10309 24513
rect 9989 24448 9997 24512
rect 10061 24448 10077 24512
rect 10141 24448 10157 24512
rect 10221 24448 10237 24512
rect 10301 24448 10309 24512
rect 9989 24447 10309 24448
rect 19322 24512 19642 24513
rect 19322 24448 19330 24512
rect 19394 24448 19410 24512
rect 19474 24448 19490 24512
rect 19554 24448 19570 24512
rect 19634 24448 19642 24512
rect 19322 24447 19642 24448
rect 26638 24442 26698 24518
rect 21118 24382 26698 24442
rect 5322 23968 5642 23969
rect 5322 23904 5330 23968
rect 5394 23904 5410 23968
rect 5474 23904 5490 23968
rect 5554 23904 5570 23968
rect 5634 23904 5642 23968
rect 5322 23903 5642 23904
rect 14656 23968 14976 23969
rect 14656 23904 14664 23968
rect 14728 23904 14744 23968
rect 14808 23904 14824 23968
rect 14888 23904 14904 23968
rect 14968 23904 14976 23968
rect 14656 23903 14976 23904
rect 10673 23626 10739 23629
rect 21118 23626 21178 24382
rect 24381 24306 24447 24309
rect 27232 24306 27712 24336
rect 24381 24304 27712 24306
rect 24381 24248 24386 24304
rect 24442 24248 27712 24304
rect 24381 24246 27712 24248
rect 24381 24243 24447 24246
rect 27232 24216 27712 24246
rect 23989 23968 24309 23969
rect 23989 23904 23997 23968
rect 24061 23904 24077 23968
rect 24141 23904 24157 23968
rect 24221 23904 24237 23968
rect 24301 23904 24309 23968
rect 23989 23903 24309 23904
rect 23737 23762 23803 23765
rect 27232 23762 27712 23792
rect 23737 23760 27712 23762
rect 23737 23704 23742 23760
rect 23798 23704 27712 23760
rect 23737 23702 27712 23704
rect 23737 23699 23803 23702
rect 27232 23672 27712 23702
rect 10673 23624 21178 23626
rect 10673 23568 10678 23624
rect 10734 23568 21178 23624
rect 10673 23566 21178 23568
rect 10673 23563 10739 23566
rect 9989 23424 10309 23425
rect 9989 23360 9997 23424
rect 10061 23360 10077 23424
rect 10141 23360 10157 23424
rect 10221 23360 10237 23424
rect 10301 23360 10309 23424
rect 9989 23359 10309 23360
rect 19322 23424 19642 23425
rect 19322 23360 19330 23424
rect 19394 23360 19410 23424
rect 19474 23360 19490 23424
rect 19554 23360 19570 23424
rect 19634 23360 19642 23424
rect 19322 23359 19642 23360
rect 19229 23218 19295 23221
rect 24473 23218 24539 23221
rect 27232 23218 27712 23248
rect 19229 23216 24539 23218
rect 19229 23160 19234 23216
rect 19290 23160 24478 23216
rect 24534 23160 24539 23216
rect 19229 23158 24539 23160
rect 19229 23155 19295 23158
rect 24473 23155 24539 23158
rect 24614 23158 27712 23218
rect 5322 22880 5642 22881
rect 5322 22816 5330 22880
rect 5394 22816 5410 22880
rect 5474 22816 5490 22880
rect 5554 22816 5570 22880
rect 5634 22816 5642 22880
rect 5322 22815 5642 22816
rect 14656 22880 14976 22881
rect 14656 22816 14664 22880
rect 14728 22816 14744 22880
rect 14808 22816 14824 22880
rect 14888 22816 14904 22880
rect 14968 22816 14976 22880
rect 14656 22815 14976 22816
rect 23989 22880 24309 22881
rect 23989 22816 23997 22880
rect 24061 22816 24077 22880
rect 24141 22816 24157 22880
rect 24221 22816 24237 22880
rect 24301 22816 24309 22880
rect 23989 22815 24309 22816
rect 24473 22674 24539 22677
rect 24614 22674 24674 23158
rect 27232 23128 27712 23158
rect 24473 22672 24674 22674
rect 24473 22616 24478 22672
rect 24534 22616 24674 22672
rect 24473 22614 24674 22616
rect 24473 22611 24539 22614
rect 10581 22538 10647 22541
rect 23185 22538 23251 22541
rect 10581 22536 23251 22538
rect 10581 22480 10586 22536
rect 10642 22480 23190 22536
rect 23246 22480 23251 22536
rect 10581 22478 23251 22480
rect 10581 22475 10647 22478
rect 23185 22475 23251 22478
rect 24749 22538 24815 22541
rect 27232 22538 27712 22568
rect 24749 22536 27712 22538
rect 24749 22480 24754 22536
rect 24810 22480 27712 22536
rect 24749 22478 27712 22480
rect 24749 22475 24815 22478
rect 27232 22448 27712 22478
rect 24381 22402 24447 22405
rect 25945 22402 26011 22405
rect 24381 22400 26011 22402
rect 24381 22344 24386 22400
rect 24442 22344 25950 22400
rect 26006 22344 26011 22400
rect 24381 22342 26011 22344
rect 24381 22339 24447 22342
rect 25945 22339 26011 22342
rect 9989 22336 10309 22337
rect 9989 22272 9997 22336
rect 10061 22272 10077 22336
rect 10141 22272 10157 22336
rect 10221 22272 10237 22336
rect 10301 22272 10309 22336
rect 9989 22271 10309 22272
rect 19322 22336 19642 22337
rect 19322 22272 19330 22336
rect 19394 22272 19410 22336
rect 19474 22272 19490 22336
rect 19554 22272 19570 22336
rect 19634 22272 19642 22336
rect 19322 22271 19642 22272
rect 12421 21994 12487 21997
rect 24657 21994 24723 21997
rect 27232 21994 27712 22024
rect 12421 21992 24723 21994
rect 12421 21936 12426 21992
rect 12482 21936 24662 21992
rect 24718 21936 24723 21992
rect 12421 21934 24723 21936
rect 12421 21931 12487 21934
rect 24657 21931 24723 21934
rect 24798 21934 27712 21994
rect 5322 21792 5642 21793
rect 5322 21728 5330 21792
rect 5394 21728 5410 21792
rect 5474 21728 5490 21792
rect 5554 21728 5570 21792
rect 5634 21728 5642 21792
rect 5322 21727 5642 21728
rect 14656 21792 14976 21793
rect 14656 21728 14664 21792
rect 14728 21728 14744 21792
rect 14808 21728 14824 21792
rect 14888 21728 14904 21792
rect 14968 21728 14976 21792
rect 14656 21727 14976 21728
rect 23989 21792 24309 21793
rect 23989 21728 23997 21792
rect 24061 21728 24077 21792
rect 24141 21728 24157 21792
rect 24221 21728 24237 21792
rect 24301 21728 24309 21792
rect 23989 21727 24309 21728
rect 23553 21586 23619 21589
rect 24798 21586 24858 21934
rect 27232 21904 27712 21934
rect 23553 21584 24858 21586
rect 23553 21528 23558 21584
rect 23614 21528 24858 21584
rect 23553 21526 24858 21528
rect 23553 21523 23619 21526
rect 12237 21450 12303 21453
rect 14721 21450 14787 21453
rect 12237 21448 14787 21450
rect 12237 21392 12242 21448
rect 12298 21392 14726 21448
rect 14782 21392 14787 21448
rect 12237 21390 14787 21392
rect 12237 21387 12303 21390
rect 14721 21387 14787 21390
rect 14997 21450 15063 21453
rect 24105 21450 24171 21453
rect 14997 21448 24171 21450
rect 14997 21392 15002 21448
rect 15058 21392 24110 21448
rect 24166 21392 24171 21448
rect 14997 21390 24171 21392
rect 14997 21387 15063 21390
rect 24105 21387 24171 21390
rect 24381 21450 24447 21453
rect 27232 21450 27712 21480
rect 24381 21448 27712 21450
rect 24381 21392 24386 21448
rect 24442 21392 27712 21448
rect 24381 21390 27712 21392
rect 24381 21387 24447 21390
rect 27232 21360 27712 21390
rect 9989 21248 10309 21249
rect 9989 21184 9997 21248
rect 10061 21184 10077 21248
rect 10141 21184 10157 21248
rect 10221 21184 10237 21248
rect 10301 21184 10309 21248
rect 9989 21183 10309 21184
rect 19322 21248 19642 21249
rect 19322 21184 19330 21248
rect 19394 21184 19410 21248
rect 19474 21184 19490 21248
rect 19554 21184 19570 21248
rect 19634 21184 19642 21248
rect 19322 21183 19642 21184
rect 9661 21042 9727 21045
rect 12329 21042 12395 21045
rect 9661 21040 12395 21042
rect 9661 20984 9666 21040
rect 9722 20984 12334 21040
rect 12390 20984 12395 21040
rect 9661 20982 12395 20984
rect 9661 20979 9727 20982
rect 12329 20979 12395 20982
rect 24473 20906 24539 20909
rect 27232 20906 27712 20936
rect 24473 20904 27712 20906
rect 24473 20848 24478 20904
rect 24534 20848 27712 20904
rect 24473 20846 27712 20848
rect 24473 20843 24539 20846
rect 27232 20816 27712 20846
rect 5322 20704 5642 20705
rect 5322 20640 5330 20704
rect 5394 20640 5410 20704
rect 5474 20640 5490 20704
rect 5554 20640 5570 20704
rect 5634 20640 5642 20704
rect 5322 20639 5642 20640
rect 14656 20704 14976 20705
rect 14656 20640 14664 20704
rect 14728 20640 14744 20704
rect 14808 20640 14824 20704
rect 14888 20640 14904 20704
rect 14968 20640 14976 20704
rect 14656 20639 14976 20640
rect 23989 20704 24309 20705
rect 23989 20640 23997 20704
rect 24061 20640 24077 20704
rect 24141 20640 24157 20704
rect 24221 20640 24237 20704
rect 24301 20640 24309 20704
rect 23989 20639 24309 20640
rect 15641 20362 15707 20365
rect 23185 20362 23251 20365
rect 27232 20362 27712 20392
rect 15641 20360 23251 20362
rect 15641 20304 15646 20360
rect 15702 20304 23190 20360
rect 23246 20304 23251 20360
rect 15641 20302 23251 20304
rect 15641 20299 15707 20302
rect 23185 20299 23251 20302
rect 24752 20302 27712 20362
rect 21437 20226 21503 20229
rect 24565 20226 24631 20229
rect 21437 20224 24631 20226
rect 21437 20168 21442 20224
rect 21498 20168 24570 20224
rect 24626 20168 24631 20224
rect 21437 20166 24631 20168
rect 21437 20163 21503 20166
rect 24565 20163 24631 20166
rect 9989 20160 10309 20161
rect 9989 20096 9997 20160
rect 10061 20096 10077 20160
rect 10141 20096 10157 20160
rect 10221 20096 10237 20160
rect 10301 20096 10309 20160
rect 9989 20095 10309 20096
rect 19322 20160 19642 20161
rect 19322 20096 19330 20160
rect 19394 20096 19410 20160
rect 19474 20096 19490 20160
rect 19554 20096 19570 20160
rect 19634 20096 19642 20160
rect 19322 20095 19642 20096
rect 11133 19818 11199 19821
rect 24752 19818 24812 20302
rect 27232 20272 27712 20302
rect 11133 19816 24812 19818
rect 11133 19760 11138 19816
rect 11194 19760 24812 19816
rect 11133 19758 24812 19760
rect 11133 19755 11199 19758
rect 24841 19682 24907 19685
rect 27232 19682 27712 19712
rect 24841 19680 27712 19682
rect 24841 19624 24846 19680
rect 24902 19624 27712 19680
rect 24841 19622 27712 19624
rect 24841 19619 24907 19622
rect 5322 19616 5642 19617
rect 5322 19552 5330 19616
rect 5394 19552 5410 19616
rect 5474 19552 5490 19616
rect 5554 19552 5570 19616
rect 5634 19552 5642 19616
rect 5322 19551 5642 19552
rect 14656 19616 14976 19617
rect 14656 19552 14664 19616
rect 14728 19552 14744 19616
rect 14808 19552 14824 19616
rect 14888 19552 14904 19616
rect 14968 19552 14976 19616
rect 14656 19551 14976 19552
rect 23989 19616 24309 19617
rect 23989 19552 23997 19616
rect 24061 19552 24077 19616
rect 24141 19552 24157 19616
rect 24221 19552 24237 19616
rect 24301 19552 24309 19616
rect 27232 19592 27712 19622
rect 23989 19551 24309 19552
rect 23686 19348 23692 19412
rect 23756 19410 23762 19412
rect 23829 19410 23895 19413
rect 23756 19408 23895 19410
rect 23756 19352 23834 19408
rect 23890 19352 23895 19408
rect 23756 19350 23895 19352
rect 23756 19348 23762 19350
rect 23829 19347 23895 19350
rect 23829 19138 23895 19141
rect 27232 19138 27712 19168
rect 23829 19136 27712 19138
rect 23829 19080 23834 19136
rect 23890 19080 27712 19136
rect 23829 19078 27712 19080
rect 23829 19075 23895 19078
rect 9989 19072 10309 19073
rect 9989 19008 9997 19072
rect 10061 19008 10077 19072
rect 10141 19008 10157 19072
rect 10221 19008 10237 19072
rect 10301 19008 10309 19072
rect 9989 19007 10309 19008
rect 19322 19072 19642 19073
rect 19322 19008 19330 19072
rect 19394 19008 19410 19072
rect 19474 19008 19490 19072
rect 19554 19008 19570 19072
rect 19634 19008 19642 19072
rect 27232 19048 27712 19078
rect 19322 19007 19642 19008
rect 15733 18866 15799 18869
rect 24105 18866 24171 18869
rect 15733 18864 24171 18866
rect 15733 18808 15738 18864
rect 15794 18808 24110 18864
rect 24166 18808 24171 18864
rect 15733 18806 24171 18808
rect 15733 18803 15799 18806
rect 24105 18803 24171 18806
rect 24381 18594 24447 18597
rect 27232 18594 27712 18624
rect 24381 18592 27712 18594
rect 24381 18536 24386 18592
rect 24442 18536 27712 18592
rect 24381 18534 27712 18536
rect 24381 18531 24447 18534
rect 5322 18528 5642 18529
rect 5322 18464 5330 18528
rect 5394 18464 5410 18528
rect 5474 18464 5490 18528
rect 5554 18464 5570 18528
rect 5634 18464 5642 18528
rect 5322 18463 5642 18464
rect 14656 18528 14976 18529
rect 14656 18464 14664 18528
rect 14728 18464 14744 18528
rect 14808 18464 14824 18528
rect 14888 18464 14904 18528
rect 14968 18464 14976 18528
rect 14656 18463 14976 18464
rect 23989 18528 24309 18529
rect 23989 18464 23997 18528
rect 24061 18464 24077 18528
rect 24141 18464 24157 18528
rect 24221 18464 24237 18528
rect 24301 18464 24309 18528
rect 27232 18504 27712 18534
rect 23989 18463 24309 18464
rect 24473 18050 24539 18053
rect 27232 18050 27712 18080
rect 24473 18048 27712 18050
rect 24473 17992 24478 18048
rect 24534 17992 27712 18048
rect 24473 17990 27712 17992
rect 24473 17987 24539 17990
rect 9989 17984 10309 17985
rect 9989 17920 9997 17984
rect 10061 17920 10077 17984
rect 10141 17920 10157 17984
rect 10221 17920 10237 17984
rect 10301 17920 10309 17984
rect 9989 17919 10309 17920
rect 19322 17984 19642 17985
rect 19322 17920 19330 17984
rect 19394 17920 19410 17984
rect 19474 17920 19490 17984
rect 19554 17920 19570 17984
rect 19634 17920 19642 17984
rect 27232 17960 27712 17990
rect 19322 17919 19642 17920
rect 16009 17642 16075 17645
rect 23829 17642 23895 17645
rect 16009 17640 23895 17642
rect 16009 17584 16014 17640
rect 16070 17584 23834 17640
rect 23890 17584 23895 17640
rect 16009 17582 23895 17584
rect 16009 17579 16075 17582
rect 23829 17579 23895 17582
rect 27232 17506 27712 17536
rect 24384 17446 27712 17506
rect 5322 17440 5642 17441
rect 5322 17376 5330 17440
rect 5394 17376 5410 17440
rect 5474 17376 5490 17440
rect 5554 17376 5570 17440
rect 5634 17376 5642 17440
rect 5322 17375 5642 17376
rect 14656 17440 14976 17441
rect 14656 17376 14664 17440
rect 14728 17376 14744 17440
rect 14808 17376 14824 17440
rect 14888 17376 14904 17440
rect 14968 17376 14976 17440
rect 14656 17375 14976 17376
rect 23989 17440 24309 17441
rect 23989 17376 23997 17440
rect 24061 17376 24077 17440
rect 24141 17376 24157 17440
rect 24221 17376 24237 17440
rect 24301 17376 24309 17440
rect 23989 17375 24309 17376
rect 16101 17370 16167 17373
rect 22449 17370 22515 17373
rect 16101 17368 22515 17370
rect 16101 17312 16106 17368
rect 16162 17312 22454 17368
rect 22510 17312 22515 17368
rect 16101 17310 22515 17312
rect 16101 17307 16167 17310
rect 22449 17307 22515 17310
rect 23829 17234 23895 17237
rect 24384 17234 24444 17446
rect 27232 17416 27712 17446
rect 23829 17232 24444 17234
rect 23829 17176 23834 17232
rect 23890 17176 24444 17232
rect 23829 17174 24444 17176
rect 23829 17171 23895 17174
rect 12881 17098 12947 17101
rect 24657 17098 24723 17101
rect 12881 17096 24723 17098
rect 12881 17040 12886 17096
rect 12942 17040 24662 17096
rect 24718 17040 24723 17096
rect 12881 17038 24723 17040
rect 12881 17035 12947 17038
rect 24657 17035 24723 17038
rect 7545 16962 7611 16965
rect 9845 16962 9911 16965
rect 7545 16960 9911 16962
rect 7545 16904 7550 16960
rect 7606 16904 9850 16960
rect 9906 16904 9911 16960
rect 7545 16902 9911 16904
rect 7545 16899 7611 16902
rect 9845 16899 9911 16902
rect 9989 16896 10309 16897
rect 9989 16832 9997 16896
rect 10061 16832 10077 16896
rect 10141 16832 10157 16896
rect 10221 16832 10237 16896
rect 10301 16832 10309 16896
rect 9989 16831 10309 16832
rect 19322 16896 19642 16897
rect 19322 16832 19330 16896
rect 19394 16832 19410 16896
rect 19474 16832 19490 16896
rect 19554 16832 19570 16896
rect 19634 16832 19642 16896
rect 19322 16831 19642 16832
rect 27232 16826 27712 16856
rect 24752 16766 27712 16826
rect 18217 16690 18283 16693
rect 24289 16690 24355 16693
rect 18217 16688 24355 16690
rect 18217 16632 18222 16688
rect 18278 16632 24294 16688
rect 24350 16632 24355 16688
rect 18217 16630 24355 16632
rect 18217 16627 18283 16630
rect 24289 16627 24355 16630
rect 24473 16690 24539 16693
rect 24752 16690 24812 16766
rect 27232 16736 27712 16766
rect 24473 16688 24812 16690
rect 24473 16632 24478 16688
rect 24534 16632 24812 16688
rect 24473 16630 24812 16632
rect 24473 16627 24539 16630
rect 13525 16554 13591 16557
rect 21529 16554 21595 16557
rect 13525 16552 21595 16554
rect 13525 16496 13530 16552
rect 13586 16496 21534 16552
rect 21590 16496 21595 16552
rect 13525 16494 21595 16496
rect 13525 16491 13591 16494
rect 21529 16491 21595 16494
rect 5322 16352 5642 16353
rect 5322 16288 5330 16352
rect 5394 16288 5410 16352
rect 5474 16288 5490 16352
rect 5554 16288 5570 16352
rect 5634 16288 5642 16352
rect 5322 16287 5642 16288
rect 14656 16352 14976 16353
rect 14656 16288 14664 16352
rect 14728 16288 14744 16352
rect 14808 16288 14824 16352
rect 14888 16288 14904 16352
rect 14968 16288 14976 16352
rect 14656 16287 14976 16288
rect 23989 16352 24309 16353
rect 23989 16288 23997 16352
rect 24061 16288 24077 16352
rect 24141 16288 24157 16352
rect 24221 16288 24237 16352
rect 24301 16288 24309 16352
rect 23989 16287 24309 16288
rect 24657 16282 24723 16285
rect 27232 16282 27712 16312
rect 24657 16280 27712 16282
rect 24657 16224 24662 16280
rect 24718 16224 27712 16280
rect 24657 16222 27712 16224
rect 24657 16219 24723 16222
rect 27232 16192 27712 16222
rect 12421 15874 12487 15877
rect 14997 15874 15063 15877
rect 12421 15872 15063 15874
rect 12421 15816 12426 15872
rect 12482 15816 15002 15872
rect 15058 15816 15063 15872
rect 12421 15814 15063 15816
rect 12421 15811 12487 15814
rect 14997 15811 15063 15814
rect 9989 15808 10309 15809
rect 9989 15744 9997 15808
rect 10061 15744 10077 15808
rect 10141 15744 10157 15808
rect 10221 15744 10237 15808
rect 10301 15744 10309 15808
rect 9989 15743 10309 15744
rect 19322 15808 19642 15809
rect 19322 15744 19330 15808
rect 19394 15744 19410 15808
rect 19474 15744 19490 15808
rect 19554 15744 19570 15808
rect 19634 15744 19642 15808
rect 19322 15743 19642 15744
rect 24381 15738 24447 15741
rect 27232 15738 27712 15768
rect 24381 15736 27712 15738
rect 24381 15680 24386 15736
rect 24442 15680 27712 15736
rect 24381 15678 27712 15680
rect 24381 15675 24447 15678
rect 27232 15648 27712 15678
rect 5322 15264 5642 15265
rect 5322 15200 5330 15264
rect 5394 15200 5410 15264
rect 5474 15200 5490 15264
rect 5554 15200 5570 15264
rect 5634 15200 5642 15264
rect 5322 15199 5642 15200
rect 14656 15264 14976 15265
rect 14656 15200 14664 15264
rect 14728 15200 14744 15264
rect 14808 15200 14824 15264
rect 14888 15200 14904 15264
rect 14968 15200 14976 15264
rect 14656 15199 14976 15200
rect 23989 15264 24309 15265
rect 23989 15200 23997 15264
rect 24061 15200 24077 15264
rect 24141 15200 24157 15264
rect 24221 15200 24237 15264
rect 24301 15200 24309 15264
rect 23989 15199 24309 15200
rect 27232 15194 27712 15224
rect 24384 15134 27712 15194
rect 23737 15058 23803 15061
rect 24384 15058 24444 15134
rect 27232 15104 27712 15134
rect 23737 15056 24444 15058
rect 23737 15000 23742 15056
rect 23798 15000 24444 15056
rect 23737 14998 24444 15000
rect 23737 14995 23803 14998
rect 13157 14922 13223 14925
rect 23093 14922 23159 14925
rect 13157 14920 23159 14922
rect 13157 14864 13162 14920
rect 13218 14864 23098 14920
rect 23154 14864 23159 14920
rect 13157 14862 23159 14864
rect 13157 14859 13223 14862
rect 23093 14859 23159 14862
rect 9989 14720 10309 14721
rect 9989 14656 9997 14720
rect 10061 14656 10077 14720
rect 10141 14656 10157 14720
rect 10221 14656 10237 14720
rect 10301 14656 10309 14720
rect 9989 14655 10309 14656
rect 19322 14720 19642 14721
rect 19322 14656 19330 14720
rect 19394 14656 19410 14720
rect 19474 14656 19490 14720
rect 19554 14656 19570 14720
rect 19634 14656 19642 14720
rect 19322 14655 19642 14656
rect 25301 14650 25367 14653
rect 27232 14650 27712 14680
rect 25301 14648 27712 14650
rect 25301 14592 25306 14648
rect 25362 14592 27712 14648
rect 25301 14590 27712 14592
rect 25301 14587 25367 14590
rect 27232 14560 27712 14590
rect 3773 14514 3839 14517
rect 15181 14514 15247 14517
rect 3773 14512 15247 14514
rect 3773 14456 3778 14512
rect 3834 14456 15186 14512
rect 15242 14456 15247 14512
rect 3773 14454 15247 14456
rect 3773 14451 3839 14454
rect 15181 14451 15247 14454
rect 5322 14176 5642 14177
rect 5322 14112 5330 14176
rect 5394 14112 5410 14176
rect 5474 14112 5490 14176
rect 5554 14112 5570 14176
rect 5634 14112 5642 14176
rect 5322 14111 5642 14112
rect 14656 14176 14976 14177
rect 14656 14112 14664 14176
rect 14728 14112 14744 14176
rect 14808 14112 14824 14176
rect 14888 14112 14904 14176
rect 14968 14112 14976 14176
rect 14656 14111 14976 14112
rect 23989 14176 24309 14177
rect 23989 14112 23997 14176
rect 24061 14112 24077 14176
rect 24141 14112 24157 14176
rect 24221 14112 24237 14176
rect 24301 14112 24309 14176
rect 23989 14111 24309 14112
rect 18585 13970 18651 13973
rect 24381 13970 24447 13973
rect 24841 13970 24907 13973
rect 27232 13970 27712 14000
rect 18585 13968 24907 13970
rect 18585 13912 18590 13968
rect 18646 13912 24386 13968
rect 24442 13912 24846 13968
rect 24902 13912 24907 13968
rect 18585 13910 24907 13912
rect 18585 13907 18651 13910
rect 24381 13907 24447 13910
rect 24841 13907 24907 13910
rect 24982 13910 27712 13970
rect 23185 13834 23251 13837
rect 24982 13834 25042 13910
rect 27232 13880 27712 13910
rect 23185 13832 25042 13834
rect 23185 13776 23190 13832
rect 23246 13776 25042 13832
rect 23185 13774 25042 13776
rect 23185 13771 23251 13774
rect 9989 13632 10309 13633
rect 9989 13568 9997 13632
rect 10061 13568 10077 13632
rect 10141 13568 10157 13632
rect 10221 13568 10237 13632
rect 10301 13568 10309 13632
rect 9989 13567 10309 13568
rect 19322 13632 19642 13633
rect 19322 13568 19330 13632
rect 19394 13568 19410 13632
rect 19474 13568 19490 13632
rect 19554 13568 19570 13632
rect 19634 13568 19642 13632
rect 19322 13567 19642 13568
rect 25393 13426 25459 13429
rect 27232 13426 27712 13456
rect 25393 13424 27712 13426
rect 25393 13368 25398 13424
rect 25454 13368 27712 13424
rect 25393 13366 27712 13368
rect 25393 13363 25459 13366
rect 27232 13336 27712 13366
rect 14997 13290 15063 13293
rect 24841 13290 24907 13293
rect 14997 13288 24907 13290
rect 14997 13232 15002 13288
rect 15058 13232 24846 13288
rect 24902 13232 24907 13288
rect 14997 13230 24907 13232
rect 14997 13227 15063 13230
rect 24841 13227 24907 13230
rect 18953 13154 19019 13157
rect 20517 13154 20583 13157
rect 18953 13152 20583 13154
rect 18953 13096 18958 13152
rect 19014 13096 20522 13152
rect 20578 13096 20583 13152
rect 18953 13094 20583 13096
rect 18953 13091 19019 13094
rect 20517 13091 20583 13094
rect 5322 13088 5642 13089
rect 5322 13024 5330 13088
rect 5394 13024 5410 13088
rect 5474 13024 5490 13088
rect 5554 13024 5570 13088
rect 5634 13024 5642 13088
rect 5322 13023 5642 13024
rect 14656 13088 14976 13089
rect 14656 13024 14664 13088
rect 14728 13024 14744 13088
rect 14808 13024 14824 13088
rect 14888 13024 14904 13088
rect 14968 13024 14976 13088
rect 14656 13023 14976 13024
rect 23989 13088 24309 13089
rect 23989 13024 23997 13088
rect 24061 13024 24077 13088
rect 24141 13024 24157 13088
rect 24221 13024 24237 13088
rect 24301 13024 24309 13088
rect 23989 13023 24309 13024
rect 21069 13018 21135 13021
rect 23737 13018 23803 13021
rect 21069 13016 23803 13018
rect 21069 12960 21074 13016
rect 21130 12960 23742 13016
rect 23798 12960 23803 13016
rect 21069 12958 23803 12960
rect 21069 12955 21135 12958
rect 23737 12955 23803 12958
rect 16653 12882 16719 12885
rect 24289 12882 24355 12885
rect 16653 12880 24355 12882
rect 16653 12824 16658 12880
rect 16714 12824 24294 12880
rect 24350 12824 24355 12880
rect 16653 12822 24355 12824
rect 16653 12819 16719 12822
rect 24289 12819 24355 12822
rect 24473 12882 24539 12885
rect 27232 12882 27712 12912
rect 24473 12880 27712 12882
rect 24473 12824 24478 12880
rect 24534 12824 27712 12880
rect 24473 12822 27712 12824
rect 24473 12819 24539 12822
rect 27232 12792 27712 12822
rect 3865 12746 3931 12749
rect 18585 12746 18651 12749
rect 3865 12744 18651 12746
rect 3865 12688 3870 12744
rect 3926 12688 18590 12744
rect 18646 12688 18651 12744
rect 3865 12686 18651 12688
rect 3865 12683 3931 12686
rect 18585 12683 18651 12686
rect 18953 12746 19019 12749
rect 23369 12746 23435 12749
rect 18953 12744 23435 12746
rect 18953 12688 18958 12744
rect 19014 12688 23374 12744
rect 23430 12688 23435 12744
rect 18953 12686 23435 12688
rect 18953 12683 19019 12686
rect 23369 12683 23435 12686
rect 9989 12544 10309 12545
rect 9989 12480 9997 12544
rect 10061 12480 10077 12544
rect 10141 12480 10157 12544
rect 10221 12480 10237 12544
rect 10301 12480 10309 12544
rect 9989 12479 10309 12480
rect 19322 12544 19642 12545
rect 19322 12480 19330 12544
rect 19394 12480 19410 12544
rect 19474 12480 19490 12544
rect 19554 12480 19570 12544
rect 19634 12480 19642 12544
rect 19322 12479 19642 12480
rect 22725 12474 22791 12477
rect 23001 12474 23067 12477
rect 22725 12472 23067 12474
rect 22725 12416 22730 12472
rect 22786 12416 23006 12472
rect 23062 12416 23067 12472
rect 22725 12414 23067 12416
rect 22725 12411 22791 12414
rect 23001 12411 23067 12414
rect 22817 12338 22883 12341
rect 27232 12338 27712 12368
rect 22817 12336 27712 12338
rect 22817 12280 22822 12336
rect 22878 12280 27712 12336
rect 22817 12278 27712 12280
rect 22817 12275 22883 12278
rect 27232 12248 27712 12278
rect 5322 12000 5642 12001
rect 5322 11936 5330 12000
rect 5394 11936 5410 12000
rect 5474 11936 5490 12000
rect 5554 11936 5570 12000
rect 5634 11936 5642 12000
rect 5322 11935 5642 11936
rect 14656 12000 14976 12001
rect 14656 11936 14664 12000
rect 14728 11936 14744 12000
rect 14808 11936 14824 12000
rect 14888 11936 14904 12000
rect 14968 11936 14976 12000
rect 14656 11935 14976 11936
rect 23989 12000 24309 12001
rect 23989 11936 23997 12000
rect 24061 11936 24077 12000
rect 24141 11936 24157 12000
rect 24221 11936 24237 12000
rect 24301 11936 24309 12000
rect 23989 11935 24309 11936
rect 15917 11794 15983 11797
rect 21713 11794 21779 11797
rect 15917 11792 21779 11794
rect 15917 11736 15922 11792
rect 15978 11736 21718 11792
rect 21774 11736 21779 11792
rect 15917 11734 21779 11736
rect 15917 11731 15983 11734
rect 21713 11731 21779 11734
rect 24473 11794 24539 11797
rect 27232 11794 27712 11824
rect 24473 11792 27712 11794
rect 24473 11736 24478 11792
rect 24534 11736 27712 11792
rect 24473 11734 27712 11736
rect 24473 11731 24539 11734
rect 27232 11704 27712 11734
rect 13617 11658 13683 11661
rect 20609 11658 20675 11661
rect 13617 11656 20675 11658
rect 13617 11600 13622 11656
rect 13678 11600 20614 11656
rect 20670 11600 20675 11656
rect 13617 11598 20675 11600
rect 13617 11595 13683 11598
rect 20609 11595 20675 11598
rect 9989 11456 10309 11457
rect 9989 11392 9997 11456
rect 10061 11392 10077 11456
rect 10141 11392 10157 11456
rect 10221 11392 10237 11456
rect 10301 11392 10309 11456
rect 9989 11391 10309 11392
rect 19322 11456 19642 11457
rect 19322 11392 19330 11456
rect 19394 11392 19410 11456
rect 19474 11392 19490 11456
rect 19554 11392 19570 11456
rect 19634 11392 19642 11456
rect 19322 11391 19642 11392
rect 14445 11386 14511 11389
rect 14997 11386 15063 11389
rect 14445 11384 15063 11386
rect 14445 11328 14450 11384
rect 14506 11328 15002 11384
rect 15058 11328 15063 11384
rect 14445 11326 15063 11328
rect 14445 11323 14511 11326
rect 14997 11323 15063 11326
rect 15273 11250 15339 11253
rect 24933 11250 24999 11253
rect 15273 11248 24999 11250
rect 15273 11192 15278 11248
rect 15334 11192 24938 11248
rect 24994 11192 24999 11248
rect 15273 11190 24999 11192
rect 15273 11187 15339 11190
rect 24933 11187 24999 11190
rect 16193 11114 16259 11117
rect 18309 11114 18375 11117
rect 22357 11114 22423 11117
rect 16193 11112 18375 11114
rect 16193 11056 16198 11112
rect 16254 11056 18314 11112
rect 18370 11056 18375 11112
rect 16193 11054 18375 11056
rect 16193 11051 16259 11054
rect 18309 11051 18375 11054
rect 18542 11112 22423 11114
rect 18542 11056 22362 11112
rect 22418 11056 22423 11112
rect 18542 11054 22423 11056
rect 16837 10978 16903 10981
rect 18542 10978 18602 11054
rect 22357 11051 22423 11054
rect 22817 11114 22883 11117
rect 27232 11114 27712 11144
rect 22817 11112 27712 11114
rect 22817 11056 22822 11112
rect 22878 11056 27712 11112
rect 22817 11054 27712 11056
rect 22817 11051 22883 11054
rect 27232 11024 27712 11054
rect 16837 10976 18602 10978
rect 16837 10920 16842 10976
rect 16898 10920 18602 10976
rect 16837 10918 18602 10920
rect 16837 10915 16903 10918
rect 5322 10912 5642 10913
rect 5322 10848 5330 10912
rect 5394 10848 5410 10912
rect 5474 10848 5490 10912
rect 5554 10848 5570 10912
rect 5634 10848 5642 10912
rect 5322 10847 5642 10848
rect 14656 10912 14976 10913
rect 14656 10848 14664 10912
rect 14728 10848 14744 10912
rect 14808 10848 14824 10912
rect 14888 10848 14904 10912
rect 14968 10848 14976 10912
rect 14656 10847 14976 10848
rect 23989 10912 24309 10913
rect 23989 10848 23997 10912
rect 24061 10848 24077 10912
rect 24141 10848 24157 10912
rect 24221 10848 24237 10912
rect 24301 10848 24309 10912
rect 23989 10847 24309 10848
rect 23829 10570 23895 10573
rect 27232 10570 27712 10600
rect 23829 10568 27712 10570
rect 23829 10512 23834 10568
rect 23890 10512 27712 10568
rect 23829 10510 27712 10512
rect 23829 10507 23895 10510
rect 27232 10480 27712 10510
rect 9989 10368 10309 10369
rect 9989 10304 9997 10368
rect 10061 10304 10077 10368
rect 10141 10304 10157 10368
rect 10221 10304 10237 10368
rect 10301 10304 10309 10368
rect 9989 10303 10309 10304
rect 19322 10368 19642 10369
rect 19322 10304 19330 10368
rect 19394 10304 19410 10368
rect 19474 10304 19490 10368
rect 19554 10304 19570 10368
rect 19634 10304 19642 10368
rect 19322 10303 19642 10304
rect 15733 10162 15799 10165
rect 24933 10162 24999 10165
rect 15733 10160 24999 10162
rect 15733 10104 15738 10160
rect 15794 10104 24938 10160
rect 24994 10104 24999 10160
rect 15733 10102 24999 10104
rect 15733 10099 15799 10102
rect 24933 10099 24999 10102
rect 24381 10026 24447 10029
rect 27232 10026 27712 10056
rect 24381 10024 27712 10026
rect 24381 9968 24386 10024
rect 24442 9968 27712 10024
rect 24381 9966 27712 9968
rect 24381 9963 24447 9966
rect 27232 9936 27712 9966
rect 5322 9824 5642 9825
rect 5322 9760 5330 9824
rect 5394 9760 5410 9824
rect 5474 9760 5490 9824
rect 5554 9760 5570 9824
rect 5634 9760 5642 9824
rect 5322 9759 5642 9760
rect 14656 9824 14976 9825
rect 14656 9760 14664 9824
rect 14728 9760 14744 9824
rect 14808 9760 14824 9824
rect 14888 9760 14904 9824
rect 14968 9760 14976 9824
rect 14656 9759 14976 9760
rect 23989 9824 24309 9825
rect 23989 9760 23997 9824
rect 24061 9760 24077 9824
rect 24141 9760 24157 9824
rect 24221 9760 24237 9824
rect 24301 9760 24309 9824
rect 23989 9759 24309 9760
rect 17849 9618 17915 9621
rect 23185 9618 23251 9621
rect 17849 9616 23251 9618
rect 17849 9560 17854 9616
rect 17910 9560 23190 9616
rect 23246 9560 23251 9616
rect 17849 9558 23251 9560
rect 17849 9555 17915 9558
rect 23185 9555 23251 9558
rect 5797 9482 5863 9485
rect 17481 9482 17547 9485
rect 5797 9480 17547 9482
rect 5797 9424 5802 9480
rect 5858 9424 17486 9480
rect 17542 9424 17547 9480
rect 5797 9422 17547 9424
rect 5797 9419 5863 9422
rect 17481 9419 17547 9422
rect 17849 9482 17915 9485
rect 27232 9482 27712 9512
rect 17849 9480 27712 9482
rect 17849 9424 17854 9480
rect 17910 9424 27712 9480
rect 17849 9422 27712 9424
rect 17849 9419 17915 9422
rect 27232 9392 27712 9422
rect 13065 9346 13131 9349
rect 18861 9346 18927 9349
rect 13065 9344 18927 9346
rect 13065 9288 13070 9344
rect 13126 9288 18866 9344
rect 18922 9288 18927 9344
rect 13065 9286 18927 9288
rect 13065 9283 13131 9286
rect 18861 9283 18927 9286
rect 9989 9280 10309 9281
rect 9989 9216 9997 9280
rect 10061 9216 10077 9280
rect 10141 9216 10157 9280
rect 10221 9216 10237 9280
rect 10301 9216 10309 9280
rect 9989 9215 10309 9216
rect 19322 9280 19642 9281
rect 19322 9216 19330 9280
rect 19394 9216 19410 9280
rect 19474 9216 19490 9280
rect 19554 9216 19570 9280
rect 19634 9216 19642 9280
rect 19322 9215 19642 9216
rect 12605 9074 12671 9077
rect 15365 9074 15431 9077
rect 12605 9072 15431 9074
rect 12605 9016 12610 9072
rect 12666 9016 15370 9072
rect 15426 9016 15431 9072
rect 12605 9014 15431 9016
rect 12605 9011 12671 9014
rect 15365 9011 15431 9014
rect 11869 8938 11935 8941
rect 20609 8938 20675 8941
rect 11869 8936 20675 8938
rect 11869 8880 11874 8936
rect 11930 8880 20614 8936
rect 20670 8880 20675 8936
rect 11869 8878 20675 8880
rect 11869 8875 11935 8878
rect 20609 8875 20675 8878
rect 24473 8938 24539 8941
rect 27232 8938 27712 8968
rect 24473 8936 27712 8938
rect 24473 8880 24478 8936
rect 24534 8880 27712 8936
rect 24473 8878 27712 8880
rect 24473 8875 24539 8878
rect 27232 8848 27712 8878
rect 17941 8802 18007 8805
rect 23461 8802 23527 8805
rect 17941 8800 23527 8802
rect 17941 8744 17946 8800
rect 18002 8744 23466 8800
rect 23522 8744 23527 8800
rect 17941 8742 23527 8744
rect 17941 8739 18007 8742
rect 23461 8739 23527 8742
rect 5322 8736 5642 8737
rect 5322 8672 5330 8736
rect 5394 8672 5410 8736
rect 5474 8672 5490 8736
rect 5554 8672 5570 8736
rect 5634 8672 5642 8736
rect 5322 8671 5642 8672
rect 14656 8736 14976 8737
rect 14656 8672 14664 8736
rect 14728 8672 14744 8736
rect 14808 8672 14824 8736
rect 14888 8672 14904 8736
rect 14968 8672 14976 8736
rect 14656 8671 14976 8672
rect 23989 8736 24309 8737
rect 23989 8672 23997 8736
rect 24061 8672 24077 8736
rect 24141 8672 24157 8736
rect 24221 8672 24237 8736
rect 24301 8672 24309 8736
rect 23989 8671 24309 8672
rect 1289 8394 1355 8397
rect 13341 8394 13407 8397
rect 1289 8392 13407 8394
rect 1289 8336 1294 8392
rect 1350 8336 13346 8392
rect 13402 8336 13407 8392
rect 1289 8334 13407 8336
rect 1289 8331 1355 8334
rect 13341 8331 13407 8334
rect 18953 8394 19019 8397
rect 20977 8394 21043 8397
rect 18953 8392 21043 8394
rect 18953 8336 18958 8392
rect 19014 8336 20982 8392
rect 21038 8336 21043 8392
rect 18953 8334 21043 8336
rect 18953 8331 19019 8334
rect 20977 8331 21043 8334
rect 23645 8258 23711 8261
rect 27232 8258 27712 8288
rect 23645 8256 27712 8258
rect 23645 8200 23650 8256
rect 23706 8200 27712 8256
rect 23645 8198 27712 8200
rect 23645 8195 23711 8198
rect 9989 8192 10309 8193
rect 9989 8128 9997 8192
rect 10061 8128 10077 8192
rect 10141 8128 10157 8192
rect 10221 8128 10237 8192
rect 10301 8128 10309 8192
rect 9989 8127 10309 8128
rect 19322 8192 19642 8193
rect 19322 8128 19330 8192
rect 19394 8128 19410 8192
rect 19474 8128 19490 8192
rect 19554 8128 19570 8192
rect 19634 8128 19642 8192
rect 27232 8168 27712 8198
rect 19322 8127 19642 8128
rect 14353 8122 14419 8125
rect 17849 8122 17915 8125
rect 14353 8120 17915 8122
rect 14353 8064 14358 8120
rect 14414 8064 17854 8120
rect 17910 8064 17915 8120
rect 14353 8062 17915 8064
rect 14353 8059 14419 8062
rect 17849 8059 17915 8062
rect 5061 7986 5127 7989
rect 23093 7986 23159 7989
rect 5061 7984 23159 7986
rect 5061 7928 5066 7984
rect 5122 7928 23098 7984
rect 23154 7928 23159 7984
rect 5061 7926 23159 7928
rect 5061 7923 5127 7926
rect 23093 7923 23159 7926
rect 8465 7850 8531 7853
rect 14353 7850 14419 7853
rect 18953 7850 19019 7853
rect 24933 7850 24999 7853
rect 8465 7848 14419 7850
rect 8465 7792 8470 7848
rect 8526 7792 14358 7848
rect 14414 7792 14419 7848
rect 8465 7790 14419 7792
rect 8465 7787 8531 7790
rect 14353 7787 14419 7790
rect 14494 7848 19019 7850
rect 14494 7792 18958 7848
rect 19014 7792 19019 7848
rect 14494 7790 19019 7792
rect 5322 7648 5642 7649
rect 5322 7584 5330 7648
rect 5394 7584 5410 7648
rect 5474 7584 5490 7648
rect 5554 7584 5570 7648
rect 5634 7584 5642 7648
rect 5322 7583 5642 7584
rect 7637 7578 7703 7581
rect 14494 7578 14554 7790
rect 18953 7787 19019 7790
rect 21992 7848 24999 7850
rect 21992 7792 24938 7848
rect 24994 7792 24999 7848
rect 21992 7790 24999 7792
rect 18217 7714 18283 7717
rect 21992 7714 22052 7790
rect 24933 7787 24999 7790
rect 18217 7712 22052 7714
rect 18217 7656 18222 7712
rect 18278 7656 22052 7712
rect 18217 7654 22052 7656
rect 25669 7714 25735 7717
rect 27232 7714 27712 7744
rect 25669 7712 27712 7714
rect 25669 7656 25674 7712
rect 25730 7656 27712 7712
rect 25669 7654 27712 7656
rect 18217 7651 18283 7654
rect 25669 7651 25735 7654
rect 14656 7648 14976 7649
rect 14656 7584 14664 7648
rect 14728 7584 14744 7648
rect 14808 7584 14824 7648
rect 14888 7584 14904 7648
rect 14968 7584 14976 7648
rect 14656 7583 14976 7584
rect 23989 7648 24309 7649
rect 23989 7584 23997 7648
rect 24061 7584 24077 7648
rect 24141 7584 24157 7648
rect 24221 7584 24237 7648
rect 24301 7584 24309 7648
rect 27232 7624 27712 7654
rect 23989 7583 24309 7584
rect 7637 7576 14554 7578
rect 7637 7520 7642 7576
rect 7698 7520 14554 7576
rect 7637 7518 14554 7520
rect 7637 7515 7703 7518
rect 9201 7442 9267 7445
rect 16469 7442 16535 7445
rect 18309 7442 18375 7445
rect 9201 7440 18375 7442
rect 9201 7384 9206 7440
rect 9262 7384 16474 7440
rect 16530 7384 18314 7440
rect 18370 7384 18375 7440
rect 9201 7382 18375 7384
rect 9201 7379 9267 7382
rect 16469 7379 16535 7382
rect 18309 7379 18375 7382
rect 19965 7442 20031 7445
rect 21989 7442 22055 7445
rect 19965 7440 22055 7442
rect 19965 7384 19970 7440
rect 20026 7384 21994 7440
rect 22050 7384 22055 7440
rect 19965 7382 22055 7384
rect 19965 7379 20031 7382
rect 21989 7379 22055 7382
rect 1933 7306 1999 7309
rect 10305 7306 10371 7309
rect 1933 7304 10371 7306
rect 1933 7248 1938 7304
rect 1994 7248 10310 7304
rect 10366 7248 10371 7304
rect 1933 7246 10371 7248
rect 1933 7243 1999 7246
rect 10305 7243 10371 7246
rect 18493 7306 18559 7309
rect 18493 7304 23248 7306
rect 18493 7248 18498 7304
rect 18554 7248 23248 7304
rect 18493 7246 23248 7248
rect 18493 7243 18559 7246
rect 19781 7170 19847 7173
rect 21529 7170 21595 7173
rect 19781 7168 21595 7170
rect 19781 7112 19786 7168
rect 19842 7112 21534 7168
rect 21590 7112 21595 7168
rect 19781 7110 21595 7112
rect 23188 7170 23248 7246
rect 27232 7170 27712 7200
rect 23188 7110 27712 7170
rect 19781 7107 19847 7110
rect 21529 7107 21595 7110
rect 9989 7104 10309 7105
rect 9989 7040 9997 7104
rect 10061 7040 10077 7104
rect 10141 7040 10157 7104
rect 10221 7040 10237 7104
rect 10301 7040 10309 7104
rect 9989 7039 10309 7040
rect 19322 7104 19642 7105
rect 19322 7040 19330 7104
rect 19394 7040 19410 7104
rect 19474 7040 19490 7104
rect 19554 7040 19570 7104
rect 19634 7040 19642 7104
rect 27232 7080 27712 7110
rect 19322 7039 19642 7040
rect 15365 6898 15431 6901
rect 21621 6898 21687 6901
rect 15365 6896 21687 6898
rect 15365 6840 15370 6896
rect 15426 6840 21626 6896
rect 21682 6840 21687 6896
rect 15365 6838 21687 6840
rect 15365 6835 15431 6838
rect 21621 6835 21687 6838
rect 10765 6762 10831 6765
rect 17113 6762 17179 6765
rect 10765 6760 17179 6762
rect 10765 6704 10770 6760
rect 10826 6704 17118 6760
rect 17174 6704 17179 6760
rect 10765 6702 17179 6704
rect 10765 6699 10831 6702
rect 17070 6699 17179 6702
rect 17297 6762 17363 6765
rect 17297 6760 24674 6762
rect 17297 6704 17302 6760
rect 17358 6704 24674 6760
rect 17297 6702 24674 6704
rect 17297 6699 17363 6702
rect 7729 6626 7795 6629
rect 13617 6626 13683 6629
rect 7729 6624 13683 6626
rect 7729 6568 7734 6624
rect 7790 6568 13622 6624
rect 13678 6568 13683 6624
rect 7729 6566 13683 6568
rect 17070 6626 17130 6699
rect 21529 6626 21595 6629
rect 17070 6624 21595 6626
rect 17070 6568 21534 6624
rect 21590 6568 21595 6624
rect 17070 6566 21595 6568
rect 24614 6626 24674 6702
rect 27232 6626 27712 6656
rect 24614 6566 27712 6626
rect 7729 6563 7795 6566
rect 13617 6563 13683 6566
rect 21529 6563 21595 6566
rect 5322 6560 5642 6561
rect 5322 6496 5330 6560
rect 5394 6496 5410 6560
rect 5474 6496 5490 6560
rect 5554 6496 5570 6560
rect 5634 6496 5642 6560
rect 5322 6495 5642 6496
rect 14656 6560 14976 6561
rect 14656 6496 14664 6560
rect 14728 6496 14744 6560
rect 14808 6496 14824 6560
rect 14888 6496 14904 6560
rect 14968 6496 14976 6560
rect 14656 6495 14976 6496
rect 23989 6560 24309 6561
rect 23989 6496 23997 6560
rect 24061 6496 24077 6560
rect 24141 6496 24157 6560
rect 24221 6496 24237 6560
rect 24301 6496 24309 6560
rect 27232 6536 27712 6566
rect 23989 6495 24309 6496
rect 15549 6490 15615 6493
rect 20885 6490 20951 6493
rect 15549 6488 20951 6490
rect 15549 6432 15554 6488
rect 15610 6432 20890 6488
rect 20946 6432 20951 6488
rect 15549 6430 20951 6432
rect 15549 6427 15615 6430
rect 20885 6427 20951 6430
rect 21713 6490 21779 6493
rect 23829 6490 23895 6493
rect 21713 6488 23895 6490
rect 21713 6432 21718 6488
rect 21774 6432 23834 6488
rect 23890 6432 23895 6488
rect 21713 6430 23895 6432
rect 21713 6427 21779 6430
rect 23829 6427 23895 6430
rect 645 6354 711 6357
rect 15917 6354 15983 6357
rect 645 6352 15983 6354
rect 645 6296 650 6352
rect 706 6296 15922 6352
rect 15978 6296 15983 6352
rect 645 6294 15983 6296
rect 645 6291 711 6294
rect 15917 6291 15983 6294
rect 18769 6354 18835 6357
rect 22357 6354 22423 6357
rect 18769 6352 22423 6354
rect 18769 6296 18774 6352
rect 18830 6296 22362 6352
rect 22418 6296 22423 6352
rect 18769 6294 22423 6296
rect 18769 6291 18835 6294
rect 22357 6291 22423 6294
rect 15825 6218 15891 6221
rect 15825 6216 23248 6218
rect 15825 6160 15830 6216
rect 15886 6160 23248 6216
rect 15825 6158 23248 6160
rect 15825 6155 15891 6158
rect 23188 6082 23248 6158
rect 27232 6082 27712 6112
rect 23188 6022 27712 6082
rect 9989 6016 10309 6017
rect 9989 5952 9997 6016
rect 10061 5952 10077 6016
rect 10141 5952 10157 6016
rect 10221 5952 10237 6016
rect 10301 5952 10309 6016
rect 9989 5951 10309 5952
rect 19322 6016 19642 6017
rect 19322 5952 19330 6016
rect 19394 5952 19410 6016
rect 19474 5952 19490 6016
rect 19554 5952 19570 6016
rect 19634 5952 19642 6016
rect 27232 5992 27712 6022
rect 19322 5951 19642 5952
rect 22173 5946 22239 5949
rect 23829 5946 23895 5949
rect 22173 5944 23895 5946
rect 22173 5888 22178 5944
rect 22234 5888 23834 5944
rect 23890 5888 23895 5944
rect 22173 5886 23895 5888
rect 22173 5883 22239 5886
rect 23829 5883 23895 5886
rect 14997 5810 15063 5813
rect 23369 5810 23435 5813
rect 14997 5808 23435 5810
rect 14997 5752 15002 5808
rect 15058 5752 23374 5808
rect 23430 5752 23435 5808
rect 14997 5750 23435 5752
rect 14997 5747 15063 5750
rect 23369 5747 23435 5750
rect 7821 5674 7887 5677
rect 11501 5674 11567 5677
rect 7821 5672 11567 5674
rect 7821 5616 7826 5672
rect 7882 5616 11506 5672
rect 11562 5616 11567 5672
rect 7821 5614 11567 5616
rect 7821 5611 7887 5614
rect 11501 5611 11567 5614
rect 19505 5674 19571 5677
rect 19689 5674 19755 5677
rect 22541 5674 22607 5677
rect 19505 5672 22607 5674
rect 19505 5616 19510 5672
rect 19566 5616 19694 5672
rect 19750 5616 22546 5672
rect 22602 5616 22607 5672
rect 19505 5614 22607 5616
rect 19505 5611 19571 5614
rect 19689 5611 19755 5614
rect 22541 5611 22607 5614
rect 16193 5538 16259 5541
rect 19137 5538 19203 5541
rect 16193 5536 19203 5538
rect 16193 5480 16198 5536
rect 16254 5480 19142 5536
rect 19198 5480 19203 5536
rect 16193 5478 19203 5480
rect 16193 5475 16259 5478
rect 19137 5475 19203 5478
rect 5322 5472 5642 5473
rect 5322 5408 5330 5472
rect 5394 5408 5410 5472
rect 5474 5408 5490 5472
rect 5554 5408 5570 5472
rect 5634 5408 5642 5472
rect 5322 5407 5642 5408
rect 14656 5472 14976 5473
rect 14656 5408 14664 5472
rect 14728 5408 14744 5472
rect 14808 5408 14824 5472
rect 14888 5408 14904 5472
rect 14968 5408 14976 5472
rect 14656 5407 14976 5408
rect 23989 5472 24309 5473
rect 23989 5408 23997 5472
rect 24061 5408 24077 5472
rect 24141 5408 24157 5472
rect 24221 5408 24237 5472
rect 24301 5408 24309 5472
rect 23989 5407 24309 5408
rect 17297 5402 17363 5405
rect 23277 5402 23343 5405
rect 27232 5402 27712 5432
rect 17297 5400 23343 5402
rect 17297 5344 17302 5400
rect 17358 5344 23282 5400
rect 23338 5344 23343 5400
rect 17297 5342 23343 5344
rect 17297 5339 17363 5342
rect 23277 5339 23343 5342
rect 24614 5342 27712 5402
rect 4509 5266 4575 5269
rect 17021 5266 17087 5269
rect 4509 5264 17087 5266
rect 4509 5208 4514 5264
rect 4570 5208 17026 5264
rect 17082 5208 17087 5264
rect 4509 5206 17087 5208
rect 4509 5203 4575 5206
rect 17021 5203 17087 5206
rect 18033 5266 18099 5269
rect 22725 5266 22791 5269
rect 18033 5264 22791 5266
rect 18033 5208 18038 5264
rect 18094 5208 22730 5264
rect 22786 5208 22791 5264
rect 18033 5206 22791 5208
rect 18033 5203 18099 5206
rect 22725 5203 22791 5206
rect 10949 5130 11015 5133
rect 16377 5130 16443 5133
rect 10949 5128 16443 5130
rect 10949 5072 10954 5128
rect 11010 5072 16382 5128
rect 16438 5072 16443 5128
rect 10949 5070 16443 5072
rect 10949 5067 11015 5070
rect 16377 5067 16443 5070
rect 16929 5130 16995 5133
rect 24614 5130 24674 5342
rect 27232 5312 27712 5342
rect 16929 5128 24674 5130
rect 16929 5072 16934 5128
rect 16990 5072 24674 5128
rect 16929 5070 24674 5072
rect 16929 5067 16995 5070
rect 7085 4994 7151 4997
rect 8005 4994 8071 4997
rect 7085 4992 8071 4994
rect 7085 4936 7090 4992
rect 7146 4936 8010 4992
rect 8066 4936 8071 4992
rect 7085 4934 8071 4936
rect 7085 4931 7151 4934
rect 8005 4931 8071 4934
rect 13893 4994 13959 4997
rect 16837 4994 16903 4997
rect 13893 4992 16903 4994
rect 13893 4936 13898 4992
rect 13954 4936 16842 4992
rect 16898 4936 16903 4992
rect 13893 4934 16903 4936
rect 13893 4931 13959 4934
rect 16837 4931 16903 4934
rect 23737 4994 23803 4997
rect 24749 4994 24815 4997
rect 23737 4992 24815 4994
rect 23737 4936 23742 4992
rect 23798 4936 24754 4992
rect 24810 4936 24815 4992
rect 23737 4934 24815 4936
rect 23737 4931 23803 4934
rect 24749 4931 24815 4934
rect 9989 4928 10309 4929
rect 9989 4864 9997 4928
rect 10061 4864 10077 4928
rect 10141 4864 10157 4928
rect 10221 4864 10237 4928
rect 10301 4864 10309 4928
rect 9989 4863 10309 4864
rect 19322 4928 19642 4929
rect 19322 4864 19330 4928
rect 19394 4864 19410 4928
rect 19474 4864 19490 4928
rect 19554 4864 19570 4928
rect 19634 4864 19642 4928
rect 19322 4863 19642 4864
rect 14353 4858 14419 4861
rect 16101 4858 16167 4861
rect 14353 4856 16167 4858
rect 14353 4800 14358 4856
rect 14414 4800 16106 4856
rect 16162 4800 16167 4856
rect 14353 4798 16167 4800
rect 14353 4795 14419 4798
rect 16101 4795 16167 4798
rect 19965 4858 20031 4861
rect 22081 4858 22147 4861
rect 24381 4858 24447 4861
rect 27232 4858 27712 4888
rect 19965 4856 24447 4858
rect 19965 4800 19970 4856
rect 20026 4800 22086 4856
rect 22142 4800 24386 4856
rect 24442 4800 24447 4856
rect 19965 4798 24447 4800
rect 19965 4795 20031 4798
rect 22081 4795 22147 4798
rect 24381 4795 24447 4798
rect 24614 4798 27712 4858
rect 11041 4722 11107 4725
rect 21989 4722 22055 4725
rect 11041 4720 22055 4722
rect 11041 4664 11046 4720
rect 11102 4664 21994 4720
rect 22050 4664 22055 4720
rect 11041 4662 22055 4664
rect 11041 4659 11107 4662
rect 21989 4659 22055 4662
rect 8833 4586 8899 4589
rect 24614 4586 24674 4798
rect 27232 4768 27712 4798
rect 8833 4584 24674 4586
rect 8833 4528 8838 4584
rect 8894 4528 24674 4584
rect 8833 4526 24674 4528
rect 8833 4523 8899 4526
rect 5061 4450 5127 4453
rect 3086 4448 5127 4450
rect 3086 4392 5066 4448
rect 5122 4392 5127 4448
rect 3086 4390 5127 4392
rect 1 4178 67 4181
rect 3086 4178 3146 4390
rect 5061 4387 5127 4390
rect 6441 4450 6507 4453
rect 14353 4450 14419 4453
rect 6441 4448 14419 4450
rect 6441 4392 6446 4448
rect 6502 4392 14358 4448
rect 14414 4392 14419 4448
rect 6441 4390 14419 4392
rect 6441 4387 6507 4390
rect 14353 4387 14419 4390
rect 15273 4450 15339 4453
rect 17205 4450 17271 4453
rect 20149 4450 20215 4453
rect 15273 4448 20215 4450
rect 15273 4392 15278 4448
rect 15334 4392 17210 4448
rect 17266 4392 20154 4448
rect 20210 4392 20215 4448
rect 15273 4390 20215 4392
rect 15273 4387 15339 4390
rect 17205 4387 17271 4390
rect 20149 4387 20215 4390
rect 5322 4384 5642 4385
rect 5322 4320 5330 4384
rect 5394 4320 5410 4384
rect 5474 4320 5490 4384
rect 5554 4320 5570 4384
rect 5634 4320 5642 4384
rect 5322 4319 5642 4320
rect 14656 4384 14976 4385
rect 14656 4320 14664 4384
rect 14728 4320 14744 4384
rect 14808 4320 14824 4384
rect 14888 4320 14904 4384
rect 14968 4320 14976 4384
rect 14656 4319 14976 4320
rect 23989 4384 24309 4385
rect 23989 4320 23997 4384
rect 24061 4320 24077 4384
rect 24141 4320 24157 4384
rect 24221 4320 24237 4384
rect 24301 4320 24309 4384
rect 23989 4319 24309 4320
rect 16285 4314 16351 4317
rect 17941 4314 18007 4317
rect 16285 4312 18007 4314
rect 16285 4256 16290 4312
rect 16346 4256 17946 4312
rect 18002 4256 18007 4312
rect 16285 4254 18007 4256
rect 16285 4251 16351 4254
rect 17941 4251 18007 4254
rect 18861 4314 18927 4317
rect 23185 4314 23251 4317
rect 18861 4312 23251 4314
rect 18861 4256 18866 4312
rect 18922 4256 23190 4312
rect 23246 4256 23251 4312
rect 18861 4254 23251 4256
rect 18861 4251 18927 4254
rect 23185 4251 23251 4254
rect 24381 4314 24447 4317
rect 27232 4314 27712 4344
rect 24381 4312 27712 4314
rect 24381 4256 24386 4312
rect 24442 4256 27712 4312
rect 24381 4254 27712 4256
rect 24381 4251 24447 4254
rect 27232 4224 27712 4254
rect 1 4176 3146 4178
rect 1 4120 6 4176
rect 62 4120 3146 4176
rect 1 4118 3146 4120
rect 3221 4178 3287 4181
rect 9753 4178 9819 4181
rect 3221 4176 9819 4178
rect 3221 4120 3226 4176
rect 3282 4120 9758 4176
rect 9814 4120 9819 4176
rect 3221 4118 9819 4120
rect 1 4115 67 4118
rect 3221 4115 3287 4118
rect 9753 4115 9819 4118
rect 11593 4178 11659 4181
rect 16929 4178 16995 4181
rect 11593 4176 16995 4178
rect 11593 4120 11598 4176
rect 11654 4120 16934 4176
rect 16990 4120 16995 4176
rect 11593 4118 16995 4120
rect 11593 4115 11659 4118
rect 16929 4115 16995 4118
rect 19873 4178 19939 4181
rect 21437 4178 21503 4181
rect 19873 4176 21503 4178
rect 19873 4120 19878 4176
rect 19934 4120 21442 4176
rect 21498 4120 21503 4176
rect 19873 4118 21503 4120
rect 19873 4115 19939 4118
rect 21437 4115 21503 4118
rect 8281 4042 8347 4045
rect 11869 4042 11935 4045
rect 8281 4040 11935 4042
rect 8281 3984 8286 4040
rect 8342 3984 11874 4040
rect 11930 3984 11935 4040
rect 8281 3982 11935 3984
rect 8281 3979 8347 3982
rect 11869 3979 11935 3982
rect 18125 4042 18191 4045
rect 20609 4042 20675 4045
rect 18125 4040 20675 4042
rect 18125 3984 18130 4040
rect 18186 3984 20614 4040
rect 20670 3984 20675 4040
rect 18125 3982 20675 3984
rect 18125 3979 18191 3982
rect 20609 3979 20675 3982
rect 2577 3906 2643 3909
rect 8373 3906 8439 3909
rect 2577 3904 8439 3906
rect 2577 3848 2582 3904
rect 2638 3848 8378 3904
rect 8434 3848 8439 3904
rect 2577 3846 8439 3848
rect 2577 3843 2643 3846
rect 8373 3843 8439 3846
rect 10397 3906 10463 3909
rect 12789 3906 12855 3909
rect 10397 3904 12855 3906
rect 10397 3848 10402 3904
rect 10458 3848 12794 3904
rect 12850 3848 12855 3904
rect 10397 3846 12855 3848
rect 10397 3843 10463 3846
rect 12789 3843 12855 3846
rect 20057 3906 20123 3909
rect 23185 3906 23251 3909
rect 20057 3904 23251 3906
rect 20057 3848 20062 3904
rect 20118 3848 23190 3904
rect 23246 3848 23251 3904
rect 20057 3846 23251 3848
rect 20057 3843 20123 3846
rect 23185 3843 23251 3846
rect 9989 3840 10309 3841
rect 9989 3776 9997 3840
rect 10061 3776 10077 3840
rect 10141 3776 10157 3840
rect 10221 3776 10237 3840
rect 10301 3776 10309 3840
rect 9989 3775 10309 3776
rect 19322 3840 19642 3841
rect 19322 3776 19330 3840
rect 19394 3776 19410 3840
rect 19474 3776 19490 3840
rect 19554 3776 19570 3840
rect 19634 3776 19642 3840
rect 19322 3775 19642 3776
rect 7729 3770 7795 3773
rect 8925 3770 8991 3773
rect 7729 3768 8991 3770
rect 7729 3712 7734 3768
rect 7790 3712 8930 3768
rect 8986 3712 8991 3768
rect 7729 3710 8991 3712
rect 7729 3707 7795 3710
rect 8925 3707 8991 3710
rect 11133 3770 11199 3773
rect 11542 3770 11548 3772
rect 11133 3768 11548 3770
rect 11133 3712 11138 3768
rect 11194 3712 11548 3768
rect 11133 3710 11548 3712
rect 11133 3707 11199 3710
rect 11542 3708 11548 3710
rect 11612 3708 11618 3772
rect 12329 3770 12395 3773
rect 17113 3770 17179 3773
rect 12329 3768 17179 3770
rect 12329 3712 12334 3768
rect 12390 3712 17118 3768
rect 17174 3712 17179 3768
rect 12329 3710 17179 3712
rect 12329 3707 12395 3710
rect 17113 3707 17179 3710
rect 21529 3770 21595 3773
rect 27232 3770 27712 3800
rect 21529 3768 27712 3770
rect 21529 3712 21534 3768
rect 21590 3712 27712 3768
rect 21529 3710 27712 3712
rect 21529 3707 21595 3710
rect 27232 3680 27712 3710
rect 9017 3634 9083 3637
rect 15365 3634 15431 3637
rect 9017 3632 15431 3634
rect 9017 3576 9022 3632
rect 9078 3576 15370 3632
rect 15426 3576 15431 3632
rect 9017 3574 15431 3576
rect 9017 3571 9083 3574
rect 15365 3571 15431 3574
rect 19689 3634 19755 3637
rect 25301 3634 25367 3637
rect 19689 3632 25367 3634
rect 19689 3576 19694 3632
rect 19750 3576 25306 3632
rect 25362 3576 25367 3632
rect 19689 3574 25367 3576
rect 19689 3571 19755 3574
rect 25301 3571 25367 3574
rect 3957 3498 4023 3501
rect 13341 3498 13407 3501
rect 3957 3496 13407 3498
rect 3957 3440 3962 3496
rect 4018 3440 13346 3496
rect 13402 3440 13407 3496
rect 3957 3438 13407 3440
rect 3957 3435 4023 3438
rect 13341 3435 13407 3438
rect 14537 3498 14603 3501
rect 18677 3498 18743 3501
rect 14537 3496 18743 3498
rect 14537 3440 14542 3496
rect 14598 3440 18682 3496
rect 18738 3440 18743 3496
rect 14537 3438 18743 3440
rect 14537 3435 14603 3438
rect 18677 3435 18743 3438
rect 20885 3498 20951 3501
rect 24841 3498 24907 3501
rect 20885 3496 24907 3498
rect 20885 3440 20890 3496
rect 20946 3440 24846 3496
rect 24902 3440 24907 3496
rect 20885 3438 24907 3440
rect 20885 3435 20951 3438
rect 24841 3435 24907 3438
rect 9845 3362 9911 3365
rect 19965 3362 20031 3365
rect 23461 3362 23527 3365
rect 9845 3360 14554 3362
rect 9845 3304 9850 3360
rect 9906 3304 14554 3360
rect 9845 3302 14554 3304
rect 9845 3299 9911 3302
rect 5322 3296 5642 3297
rect 5322 3232 5330 3296
rect 5394 3232 5410 3296
rect 5474 3232 5490 3296
rect 5554 3232 5570 3296
rect 5634 3232 5642 3296
rect 5322 3231 5642 3232
rect 14494 3090 14554 3302
rect 19965 3360 23527 3362
rect 19965 3304 19970 3360
rect 20026 3304 23466 3360
rect 23522 3304 23527 3360
rect 19965 3302 23527 3304
rect 19965 3299 20031 3302
rect 23461 3299 23527 3302
rect 14656 3296 14976 3297
rect 14656 3232 14664 3296
rect 14728 3232 14744 3296
rect 14808 3232 14824 3296
rect 14888 3232 14904 3296
rect 14968 3232 14976 3296
rect 14656 3231 14976 3232
rect 23989 3296 24309 3297
rect 23989 3232 23997 3296
rect 24061 3232 24077 3296
rect 24141 3232 24157 3296
rect 24221 3232 24237 3296
rect 24301 3232 24309 3296
rect 23989 3231 24309 3232
rect 16377 3226 16443 3229
rect 19229 3226 19295 3229
rect 16377 3224 19295 3226
rect 16377 3168 16382 3224
rect 16438 3168 19234 3224
rect 19290 3168 19295 3224
rect 16377 3166 19295 3168
rect 16377 3163 16443 3166
rect 19229 3163 19295 3166
rect 25025 3226 25091 3229
rect 27232 3226 27712 3256
rect 25025 3224 27712 3226
rect 25025 3168 25030 3224
rect 25086 3168 27712 3224
rect 25025 3166 27712 3168
rect 25025 3163 25091 3166
rect 27232 3136 27712 3166
rect 17481 3090 17547 3093
rect 14494 3088 17547 3090
rect 14494 3032 17486 3088
rect 17542 3032 17547 3088
rect 14494 3030 17547 3032
rect 17481 3027 17547 3030
rect 20701 3090 20767 3093
rect 23921 3090 23987 3093
rect 20701 3088 23987 3090
rect 20701 3032 20706 3088
rect 20762 3032 23926 3088
rect 23982 3032 23987 3088
rect 20701 3030 23987 3032
rect 20701 3027 20767 3030
rect 23921 3027 23987 3030
rect 7177 2954 7243 2957
rect 11869 2954 11935 2957
rect 7177 2952 11935 2954
rect 7177 2896 7182 2952
rect 7238 2896 11874 2952
rect 11930 2896 11935 2952
rect 7177 2894 11935 2896
rect 7177 2891 7243 2894
rect 11869 2891 11935 2894
rect 12881 2954 12947 2957
rect 14997 2954 15063 2957
rect 12881 2952 15063 2954
rect 12881 2896 12886 2952
rect 12942 2896 15002 2952
rect 15058 2896 15063 2952
rect 12881 2894 15063 2896
rect 12881 2891 12947 2894
rect 14997 2891 15063 2894
rect 16745 2954 16811 2957
rect 23369 2954 23435 2957
rect 24657 2956 24723 2957
rect 24606 2954 24612 2956
rect 16745 2952 23435 2954
rect 16745 2896 16750 2952
rect 16806 2896 23374 2952
rect 23430 2896 23435 2952
rect 16745 2894 23435 2896
rect 24566 2894 24612 2954
rect 24676 2952 24723 2956
rect 24718 2896 24723 2952
rect 16745 2891 16811 2894
rect 23369 2891 23435 2894
rect 24606 2892 24612 2894
rect 24676 2892 24723 2896
rect 24657 2891 24723 2892
rect 10489 2818 10555 2821
rect 19137 2818 19203 2821
rect 10489 2816 19203 2818
rect 10489 2760 10494 2816
rect 10550 2760 19142 2816
rect 19198 2760 19203 2816
rect 10489 2758 19203 2760
rect 10489 2755 10555 2758
rect 19137 2755 19203 2758
rect 25117 2818 25183 2821
rect 27233 2818 27299 2821
rect 25117 2816 27299 2818
rect 25117 2760 25122 2816
rect 25178 2760 27238 2816
rect 27294 2760 27299 2816
rect 25117 2758 27299 2760
rect 25117 2755 25183 2758
rect 27233 2755 27299 2758
rect 9989 2752 10309 2753
rect 9989 2688 9997 2752
rect 10061 2688 10077 2752
rect 10141 2688 10157 2752
rect 10221 2688 10237 2752
rect 10301 2688 10309 2752
rect 9989 2687 10309 2688
rect 19322 2752 19642 2753
rect 19322 2688 19330 2752
rect 19394 2688 19410 2752
rect 19474 2688 19490 2752
rect 19554 2688 19570 2752
rect 19634 2688 19642 2752
rect 19322 2687 19642 2688
rect 10673 2682 10739 2685
rect 12605 2682 12671 2685
rect 10673 2680 12671 2682
rect 10673 2624 10678 2680
rect 10734 2624 12610 2680
rect 12666 2624 12671 2680
rect 10673 2622 12671 2624
rect 10673 2619 10739 2622
rect 12605 2619 12671 2622
rect 13065 2682 13131 2685
rect 16561 2682 16627 2685
rect 13065 2680 16627 2682
rect 13065 2624 13070 2680
rect 13126 2624 16566 2680
rect 16622 2624 16627 2680
rect 13065 2622 16627 2624
rect 13065 2619 13131 2622
rect 16561 2619 16627 2622
rect 20793 2682 20859 2685
rect 24197 2682 24263 2685
rect 20793 2680 24263 2682
rect 20793 2624 20798 2680
rect 20854 2624 24202 2680
rect 24258 2624 24263 2680
rect 20793 2622 24263 2624
rect 20793 2619 20859 2622
rect 24197 2619 24263 2622
rect 18309 2546 18375 2549
rect 21713 2546 21779 2549
rect 18309 2544 21779 2546
rect 18309 2488 18314 2544
rect 18370 2488 21718 2544
rect 21774 2488 21779 2544
rect 18309 2486 21779 2488
rect 18309 2483 18375 2486
rect 21713 2483 21779 2486
rect 21897 2546 21963 2549
rect 27232 2546 27712 2576
rect 21897 2544 27712 2546
rect 21897 2488 21902 2544
rect 21958 2488 27712 2544
rect 21897 2486 27712 2488
rect 21897 2483 21963 2486
rect 27232 2456 27712 2486
rect 7821 2410 7887 2413
rect 24105 2410 24171 2413
rect 7821 2408 24171 2410
rect 7821 2352 7826 2408
rect 7882 2352 24110 2408
rect 24166 2352 24171 2408
rect 7821 2350 24171 2352
rect 7821 2347 7887 2350
rect 24105 2347 24171 2350
rect 8281 2274 8347 2277
rect 10305 2274 10371 2277
rect 8281 2272 10371 2274
rect 8281 2216 8286 2272
rect 8342 2216 10310 2272
rect 10366 2216 10371 2272
rect 8281 2214 10371 2216
rect 8281 2211 8347 2214
rect 10305 2211 10371 2214
rect 5322 2208 5642 2209
rect 5322 2144 5330 2208
rect 5394 2144 5410 2208
rect 5474 2144 5490 2208
rect 5554 2144 5570 2208
rect 5634 2144 5642 2208
rect 5322 2143 5642 2144
rect 14656 2208 14976 2209
rect 14656 2144 14664 2208
rect 14728 2144 14744 2208
rect 14808 2144 14824 2208
rect 14888 2144 14904 2208
rect 14968 2144 14976 2208
rect 14656 2143 14976 2144
rect 23989 2208 24309 2209
rect 23989 2144 23997 2208
rect 24061 2144 24077 2208
rect 24141 2144 24157 2208
rect 24221 2144 24237 2208
rect 24301 2144 24309 2208
rect 23989 2143 24309 2144
rect 8373 2138 8439 2141
rect 10489 2138 10555 2141
rect 8373 2136 10555 2138
rect 8373 2080 8378 2136
rect 8434 2080 10494 2136
rect 10550 2080 10555 2136
rect 8373 2078 10555 2080
rect 8373 2075 8439 2078
rect 10489 2075 10555 2078
rect 8649 2002 8715 2005
rect 25301 2002 25367 2005
rect 27232 2002 27712 2032
rect 8649 2000 25367 2002
rect 8649 1944 8654 2000
rect 8710 1944 25306 2000
rect 25362 1944 25367 2000
rect 8649 1942 25367 1944
rect 8649 1939 8715 1942
rect 25301 1939 25367 1942
rect 25534 1942 27712 2002
rect 8557 1866 8623 1869
rect 20149 1866 20215 1869
rect 8557 1864 20215 1866
rect 8557 1808 8562 1864
rect 8618 1808 20154 1864
rect 20210 1808 20215 1864
rect 8557 1806 20215 1808
rect 8557 1803 8623 1806
rect 20149 1803 20215 1806
rect 23645 1866 23711 1869
rect 25534 1866 25594 1942
rect 27232 1912 27712 1942
rect 23645 1864 25594 1866
rect 23645 1808 23650 1864
rect 23706 1808 25594 1864
rect 23645 1806 25594 1808
rect 23645 1803 23711 1806
rect 8189 1730 8255 1733
rect 24565 1730 24631 1733
rect 8189 1728 24631 1730
rect 8189 1672 8194 1728
rect 8250 1672 24570 1728
rect 24626 1672 24631 1728
rect 8189 1670 24631 1672
rect 8189 1667 8255 1670
rect 24565 1667 24631 1670
rect 8465 1594 8531 1597
rect 20241 1594 20307 1597
rect 8465 1592 20307 1594
rect 8465 1536 8470 1592
rect 8526 1536 20246 1592
rect 20302 1536 20307 1592
rect 8465 1534 20307 1536
rect 8465 1531 8531 1534
rect 20241 1531 20307 1534
rect 10397 1458 10463 1461
rect 13617 1458 13683 1461
rect 10397 1456 13683 1458
rect 10397 1400 10402 1456
rect 10458 1400 13622 1456
rect 13678 1400 13683 1456
rect 10397 1398 13683 1400
rect 10397 1395 10463 1398
rect 13617 1395 13683 1398
rect 23461 1458 23527 1461
rect 27232 1458 27712 1488
rect 23461 1456 27712 1458
rect 23461 1400 23466 1456
rect 23522 1400 27712 1456
rect 23461 1398 27712 1400
rect 23461 1395 23527 1398
rect 27232 1368 27712 1398
rect 24473 914 24539 917
rect 27232 914 27712 944
rect 24473 912 27712 914
rect 24473 856 24478 912
rect 24534 856 27712 912
rect 24473 854 27712 856
rect 24473 851 24539 854
rect 27232 824 27712 854
rect 23829 370 23895 373
rect 27232 370 27712 400
rect 23829 368 27712 370
rect 23829 312 23834 368
rect 23890 312 27712 368
rect 23829 310 27712 312
rect 23829 307 23895 310
rect 27232 280 27712 310
<< via3 >>
rect 23692 27644 23756 27708
rect 9997 25596 10061 25600
rect 9997 25540 10001 25596
rect 10001 25540 10057 25596
rect 10057 25540 10061 25596
rect 9997 25536 10061 25540
rect 10077 25596 10141 25600
rect 10077 25540 10081 25596
rect 10081 25540 10137 25596
rect 10137 25540 10141 25596
rect 10077 25536 10141 25540
rect 10157 25596 10221 25600
rect 10157 25540 10161 25596
rect 10161 25540 10217 25596
rect 10217 25540 10221 25596
rect 10157 25536 10221 25540
rect 10237 25596 10301 25600
rect 10237 25540 10241 25596
rect 10241 25540 10297 25596
rect 10297 25540 10301 25596
rect 10237 25536 10301 25540
rect 19330 25596 19394 25600
rect 19330 25540 19334 25596
rect 19334 25540 19390 25596
rect 19390 25540 19394 25596
rect 19330 25536 19394 25540
rect 19410 25596 19474 25600
rect 19410 25540 19414 25596
rect 19414 25540 19470 25596
rect 19470 25540 19474 25596
rect 19410 25536 19474 25540
rect 19490 25596 19554 25600
rect 19490 25540 19494 25596
rect 19494 25540 19550 25596
rect 19550 25540 19554 25596
rect 19490 25536 19554 25540
rect 19570 25596 19634 25600
rect 19570 25540 19574 25596
rect 19574 25540 19630 25596
rect 19630 25540 19634 25596
rect 19570 25536 19634 25540
rect 5330 25052 5394 25056
rect 5330 24996 5334 25052
rect 5334 24996 5390 25052
rect 5390 24996 5394 25052
rect 5330 24992 5394 24996
rect 5410 25052 5474 25056
rect 5410 24996 5414 25052
rect 5414 24996 5470 25052
rect 5470 24996 5474 25052
rect 5410 24992 5474 24996
rect 5490 25052 5554 25056
rect 5490 24996 5494 25052
rect 5494 24996 5550 25052
rect 5550 24996 5554 25052
rect 5490 24992 5554 24996
rect 5570 25052 5634 25056
rect 5570 24996 5574 25052
rect 5574 24996 5630 25052
rect 5630 24996 5634 25052
rect 5570 24992 5634 24996
rect 14664 25052 14728 25056
rect 14664 24996 14668 25052
rect 14668 24996 14724 25052
rect 14724 24996 14728 25052
rect 14664 24992 14728 24996
rect 14744 25052 14808 25056
rect 14744 24996 14748 25052
rect 14748 24996 14804 25052
rect 14804 24996 14808 25052
rect 14744 24992 14808 24996
rect 14824 25052 14888 25056
rect 14824 24996 14828 25052
rect 14828 24996 14884 25052
rect 14884 24996 14888 25052
rect 14824 24992 14888 24996
rect 14904 25052 14968 25056
rect 14904 24996 14908 25052
rect 14908 24996 14964 25052
rect 14964 24996 14968 25052
rect 14904 24992 14968 24996
rect 23997 25052 24061 25056
rect 23997 24996 24001 25052
rect 24001 24996 24057 25052
rect 24057 24996 24061 25052
rect 23997 24992 24061 24996
rect 24077 25052 24141 25056
rect 24077 24996 24081 25052
rect 24081 24996 24137 25052
rect 24137 24996 24141 25052
rect 24077 24992 24141 24996
rect 24157 25052 24221 25056
rect 24157 24996 24161 25052
rect 24161 24996 24217 25052
rect 24217 24996 24221 25052
rect 24157 24992 24221 24996
rect 24237 25052 24301 25056
rect 24237 24996 24241 25052
rect 24241 24996 24297 25052
rect 24297 24996 24301 25052
rect 24237 24992 24301 24996
rect 9997 24508 10061 24512
rect 9997 24452 10001 24508
rect 10001 24452 10057 24508
rect 10057 24452 10061 24508
rect 9997 24448 10061 24452
rect 10077 24508 10141 24512
rect 10077 24452 10081 24508
rect 10081 24452 10137 24508
rect 10137 24452 10141 24508
rect 10077 24448 10141 24452
rect 10157 24508 10221 24512
rect 10157 24452 10161 24508
rect 10161 24452 10217 24508
rect 10217 24452 10221 24508
rect 10157 24448 10221 24452
rect 10237 24508 10301 24512
rect 10237 24452 10241 24508
rect 10241 24452 10297 24508
rect 10297 24452 10301 24508
rect 10237 24448 10301 24452
rect 19330 24508 19394 24512
rect 19330 24452 19334 24508
rect 19334 24452 19390 24508
rect 19390 24452 19394 24508
rect 19330 24448 19394 24452
rect 19410 24508 19474 24512
rect 19410 24452 19414 24508
rect 19414 24452 19470 24508
rect 19470 24452 19474 24508
rect 19410 24448 19474 24452
rect 19490 24508 19554 24512
rect 19490 24452 19494 24508
rect 19494 24452 19550 24508
rect 19550 24452 19554 24508
rect 19490 24448 19554 24452
rect 19570 24508 19634 24512
rect 19570 24452 19574 24508
rect 19574 24452 19630 24508
rect 19630 24452 19634 24508
rect 19570 24448 19634 24452
rect 5330 23964 5394 23968
rect 5330 23908 5334 23964
rect 5334 23908 5390 23964
rect 5390 23908 5394 23964
rect 5330 23904 5394 23908
rect 5410 23964 5474 23968
rect 5410 23908 5414 23964
rect 5414 23908 5470 23964
rect 5470 23908 5474 23964
rect 5410 23904 5474 23908
rect 5490 23964 5554 23968
rect 5490 23908 5494 23964
rect 5494 23908 5550 23964
rect 5550 23908 5554 23964
rect 5490 23904 5554 23908
rect 5570 23964 5634 23968
rect 5570 23908 5574 23964
rect 5574 23908 5630 23964
rect 5630 23908 5634 23964
rect 5570 23904 5634 23908
rect 14664 23964 14728 23968
rect 14664 23908 14668 23964
rect 14668 23908 14724 23964
rect 14724 23908 14728 23964
rect 14664 23904 14728 23908
rect 14744 23964 14808 23968
rect 14744 23908 14748 23964
rect 14748 23908 14804 23964
rect 14804 23908 14808 23964
rect 14744 23904 14808 23908
rect 14824 23964 14888 23968
rect 14824 23908 14828 23964
rect 14828 23908 14884 23964
rect 14884 23908 14888 23964
rect 14824 23904 14888 23908
rect 14904 23964 14968 23968
rect 14904 23908 14908 23964
rect 14908 23908 14964 23964
rect 14964 23908 14968 23964
rect 14904 23904 14968 23908
rect 23997 23964 24061 23968
rect 23997 23908 24001 23964
rect 24001 23908 24057 23964
rect 24057 23908 24061 23964
rect 23997 23904 24061 23908
rect 24077 23964 24141 23968
rect 24077 23908 24081 23964
rect 24081 23908 24137 23964
rect 24137 23908 24141 23964
rect 24077 23904 24141 23908
rect 24157 23964 24221 23968
rect 24157 23908 24161 23964
rect 24161 23908 24217 23964
rect 24217 23908 24221 23964
rect 24157 23904 24221 23908
rect 24237 23964 24301 23968
rect 24237 23908 24241 23964
rect 24241 23908 24297 23964
rect 24297 23908 24301 23964
rect 24237 23904 24301 23908
rect 9997 23420 10061 23424
rect 9997 23364 10001 23420
rect 10001 23364 10057 23420
rect 10057 23364 10061 23420
rect 9997 23360 10061 23364
rect 10077 23420 10141 23424
rect 10077 23364 10081 23420
rect 10081 23364 10137 23420
rect 10137 23364 10141 23420
rect 10077 23360 10141 23364
rect 10157 23420 10221 23424
rect 10157 23364 10161 23420
rect 10161 23364 10217 23420
rect 10217 23364 10221 23420
rect 10157 23360 10221 23364
rect 10237 23420 10301 23424
rect 10237 23364 10241 23420
rect 10241 23364 10297 23420
rect 10297 23364 10301 23420
rect 10237 23360 10301 23364
rect 19330 23420 19394 23424
rect 19330 23364 19334 23420
rect 19334 23364 19390 23420
rect 19390 23364 19394 23420
rect 19330 23360 19394 23364
rect 19410 23420 19474 23424
rect 19410 23364 19414 23420
rect 19414 23364 19470 23420
rect 19470 23364 19474 23420
rect 19410 23360 19474 23364
rect 19490 23420 19554 23424
rect 19490 23364 19494 23420
rect 19494 23364 19550 23420
rect 19550 23364 19554 23420
rect 19490 23360 19554 23364
rect 19570 23420 19634 23424
rect 19570 23364 19574 23420
rect 19574 23364 19630 23420
rect 19630 23364 19634 23420
rect 19570 23360 19634 23364
rect 5330 22876 5394 22880
rect 5330 22820 5334 22876
rect 5334 22820 5390 22876
rect 5390 22820 5394 22876
rect 5330 22816 5394 22820
rect 5410 22876 5474 22880
rect 5410 22820 5414 22876
rect 5414 22820 5470 22876
rect 5470 22820 5474 22876
rect 5410 22816 5474 22820
rect 5490 22876 5554 22880
rect 5490 22820 5494 22876
rect 5494 22820 5550 22876
rect 5550 22820 5554 22876
rect 5490 22816 5554 22820
rect 5570 22876 5634 22880
rect 5570 22820 5574 22876
rect 5574 22820 5630 22876
rect 5630 22820 5634 22876
rect 5570 22816 5634 22820
rect 14664 22876 14728 22880
rect 14664 22820 14668 22876
rect 14668 22820 14724 22876
rect 14724 22820 14728 22876
rect 14664 22816 14728 22820
rect 14744 22876 14808 22880
rect 14744 22820 14748 22876
rect 14748 22820 14804 22876
rect 14804 22820 14808 22876
rect 14744 22816 14808 22820
rect 14824 22876 14888 22880
rect 14824 22820 14828 22876
rect 14828 22820 14884 22876
rect 14884 22820 14888 22876
rect 14824 22816 14888 22820
rect 14904 22876 14968 22880
rect 14904 22820 14908 22876
rect 14908 22820 14964 22876
rect 14964 22820 14968 22876
rect 14904 22816 14968 22820
rect 23997 22876 24061 22880
rect 23997 22820 24001 22876
rect 24001 22820 24057 22876
rect 24057 22820 24061 22876
rect 23997 22816 24061 22820
rect 24077 22876 24141 22880
rect 24077 22820 24081 22876
rect 24081 22820 24137 22876
rect 24137 22820 24141 22876
rect 24077 22816 24141 22820
rect 24157 22876 24221 22880
rect 24157 22820 24161 22876
rect 24161 22820 24217 22876
rect 24217 22820 24221 22876
rect 24157 22816 24221 22820
rect 24237 22876 24301 22880
rect 24237 22820 24241 22876
rect 24241 22820 24297 22876
rect 24297 22820 24301 22876
rect 24237 22816 24301 22820
rect 9997 22332 10061 22336
rect 9997 22276 10001 22332
rect 10001 22276 10057 22332
rect 10057 22276 10061 22332
rect 9997 22272 10061 22276
rect 10077 22332 10141 22336
rect 10077 22276 10081 22332
rect 10081 22276 10137 22332
rect 10137 22276 10141 22332
rect 10077 22272 10141 22276
rect 10157 22332 10221 22336
rect 10157 22276 10161 22332
rect 10161 22276 10217 22332
rect 10217 22276 10221 22332
rect 10157 22272 10221 22276
rect 10237 22332 10301 22336
rect 10237 22276 10241 22332
rect 10241 22276 10297 22332
rect 10297 22276 10301 22332
rect 10237 22272 10301 22276
rect 19330 22332 19394 22336
rect 19330 22276 19334 22332
rect 19334 22276 19390 22332
rect 19390 22276 19394 22332
rect 19330 22272 19394 22276
rect 19410 22332 19474 22336
rect 19410 22276 19414 22332
rect 19414 22276 19470 22332
rect 19470 22276 19474 22332
rect 19410 22272 19474 22276
rect 19490 22332 19554 22336
rect 19490 22276 19494 22332
rect 19494 22276 19550 22332
rect 19550 22276 19554 22332
rect 19490 22272 19554 22276
rect 19570 22332 19634 22336
rect 19570 22276 19574 22332
rect 19574 22276 19630 22332
rect 19630 22276 19634 22332
rect 19570 22272 19634 22276
rect 5330 21788 5394 21792
rect 5330 21732 5334 21788
rect 5334 21732 5390 21788
rect 5390 21732 5394 21788
rect 5330 21728 5394 21732
rect 5410 21788 5474 21792
rect 5410 21732 5414 21788
rect 5414 21732 5470 21788
rect 5470 21732 5474 21788
rect 5410 21728 5474 21732
rect 5490 21788 5554 21792
rect 5490 21732 5494 21788
rect 5494 21732 5550 21788
rect 5550 21732 5554 21788
rect 5490 21728 5554 21732
rect 5570 21788 5634 21792
rect 5570 21732 5574 21788
rect 5574 21732 5630 21788
rect 5630 21732 5634 21788
rect 5570 21728 5634 21732
rect 14664 21788 14728 21792
rect 14664 21732 14668 21788
rect 14668 21732 14724 21788
rect 14724 21732 14728 21788
rect 14664 21728 14728 21732
rect 14744 21788 14808 21792
rect 14744 21732 14748 21788
rect 14748 21732 14804 21788
rect 14804 21732 14808 21788
rect 14744 21728 14808 21732
rect 14824 21788 14888 21792
rect 14824 21732 14828 21788
rect 14828 21732 14884 21788
rect 14884 21732 14888 21788
rect 14824 21728 14888 21732
rect 14904 21788 14968 21792
rect 14904 21732 14908 21788
rect 14908 21732 14964 21788
rect 14964 21732 14968 21788
rect 14904 21728 14968 21732
rect 23997 21788 24061 21792
rect 23997 21732 24001 21788
rect 24001 21732 24057 21788
rect 24057 21732 24061 21788
rect 23997 21728 24061 21732
rect 24077 21788 24141 21792
rect 24077 21732 24081 21788
rect 24081 21732 24137 21788
rect 24137 21732 24141 21788
rect 24077 21728 24141 21732
rect 24157 21788 24221 21792
rect 24157 21732 24161 21788
rect 24161 21732 24217 21788
rect 24217 21732 24221 21788
rect 24157 21728 24221 21732
rect 24237 21788 24301 21792
rect 24237 21732 24241 21788
rect 24241 21732 24297 21788
rect 24297 21732 24301 21788
rect 24237 21728 24301 21732
rect 9997 21244 10061 21248
rect 9997 21188 10001 21244
rect 10001 21188 10057 21244
rect 10057 21188 10061 21244
rect 9997 21184 10061 21188
rect 10077 21244 10141 21248
rect 10077 21188 10081 21244
rect 10081 21188 10137 21244
rect 10137 21188 10141 21244
rect 10077 21184 10141 21188
rect 10157 21244 10221 21248
rect 10157 21188 10161 21244
rect 10161 21188 10217 21244
rect 10217 21188 10221 21244
rect 10157 21184 10221 21188
rect 10237 21244 10301 21248
rect 10237 21188 10241 21244
rect 10241 21188 10297 21244
rect 10297 21188 10301 21244
rect 10237 21184 10301 21188
rect 19330 21244 19394 21248
rect 19330 21188 19334 21244
rect 19334 21188 19390 21244
rect 19390 21188 19394 21244
rect 19330 21184 19394 21188
rect 19410 21244 19474 21248
rect 19410 21188 19414 21244
rect 19414 21188 19470 21244
rect 19470 21188 19474 21244
rect 19410 21184 19474 21188
rect 19490 21244 19554 21248
rect 19490 21188 19494 21244
rect 19494 21188 19550 21244
rect 19550 21188 19554 21244
rect 19490 21184 19554 21188
rect 19570 21244 19634 21248
rect 19570 21188 19574 21244
rect 19574 21188 19630 21244
rect 19630 21188 19634 21244
rect 19570 21184 19634 21188
rect 5330 20700 5394 20704
rect 5330 20644 5334 20700
rect 5334 20644 5390 20700
rect 5390 20644 5394 20700
rect 5330 20640 5394 20644
rect 5410 20700 5474 20704
rect 5410 20644 5414 20700
rect 5414 20644 5470 20700
rect 5470 20644 5474 20700
rect 5410 20640 5474 20644
rect 5490 20700 5554 20704
rect 5490 20644 5494 20700
rect 5494 20644 5550 20700
rect 5550 20644 5554 20700
rect 5490 20640 5554 20644
rect 5570 20700 5634 20704
rect 5570 20644 5574 20700
rect 5574 20644 5630 20700
rect 5630 20644 5634 20700
rect 5570 20640 5634 20644
rect 14664 20700 14728 20704
rect 14664 20644 14668 20700
rect 14668 20644 14724 20700
rect 14724 20644 14728 20700
rect 14664 20640 14728 20644
rect 14744 20700 14808 20704
rect 14744 20644 14748 20700
rect 14748 20644 14804 20700
rect 14804 20644 14808 20700
rect 14744 20640 14808 20644
rect 14824 20700 14888 20704
rect 14824 20644 14828 20700
rect 14828 20644 14884 20700
rect 14884 20644 14888 20700
rect 14824 20640 14888 20644
rect 14904 20700 14968 20704
rect 14904 20644 14908 20700
rect 14908 20644 14964 20700
rect 14964 20644 14968 20700
rect 14904 20640 14968 20644
rect 23997 20700 24061 20704
rect 23997 20644 24001 20700
rect 24001 20644 24057 20700
rect 24057 20644 24061 20700
rect 23997 20640 24061 20644
rect 24077 20700 24141 20704
rect 24077 20644 24081 20700
rect 24081 20644 24137 20700
rect 24137 20644 24141 20700
rect 24077 20640 24141 20644
rect 24157 20700 24221 20704
rect 24157 20644 24161 20700
rect 24161 20644 24217 20700
rect 24217 20644 24221 20700
rect 24157 20640 24221 20644
rect 24237 20700 24301 20704
rect 24237 20644 24241 20700
rect 24241 20644 24297 20700
rect 24297 20644 24301 20700
rect 24237 20640 24301 20644
rect 9997 20156 10061 20160
rect 9997 20100 10001 20156
rect 10001 20100 10057 20156
rect 10057 20100 10061 20156
rect 9997 20096 10061 20100
rect 10077 20156 10141 20160
rect 10077 20100 10081 20156
rect 10081 20100 10137 20156
rect 10137 20100 10141 20156
rect 10077 20096 10141 20100
rect 10157 20156 10221 20160
rect 10157 20100 10161 20156
rect 10161 20100 10217 20156
rect 10217 20100 10221 20156
rect 10157 20096 10221 20100
rect 10237 20156 10301 20160
rect 10237 20100 10241 20156
rect 10241 20100 10297 20156
rect 10297 20100 10301 20156
rect 10237 20096 10301 20100
rect 19330 20156 19394 20160
rect 19330 20100 19334 20156
rect 19334 20100 19390 20156
rect 19390 20100 19394 20156
rect 19330 20096 19394 20100
rect 19410 20156 19474 20160
rect 19410 20100 19414 20156
rect 19414 20100 19470 20156
rect 19470 20100 19474 20156
rect 19410 20096 19474 20100
rect 19490 20156 19554 20160
rect 19490 20100 19494 20156
rect 19494 20100 19550 20156
rect 19550 20100 19554 20156
rect 19490 20096 19554 20100
rect 19570 20156 19634 20160
rect 19570 20100 19574 20156
rect 19574 20100 19630 20156
rect 19630 20100 19634 20156
rect 19570 20096 19634 20100
rect 5330 19612 5394 19616
rect 5330 19556 5334 19612
rect 5334 19556 5390 19612
rect 5390 19556 5394 19612
rect 5330 19552 5394 19556
rect 5410 19612 5474 19616
rect 5410 19556 5414 19612
rect 5414 19556 5470 19612
rect 5470 19556 5474 19612
rect 5410 19552 5474 19556
rect 5490 19612 5554 19616
rect 5490 19556 5494 19612
rect 5494 19556 5550 19612
rect 5550 19556 5554 19612
rect 5490 19552 5554 19556
rect 5570 19612 5634 19616
rect 5570 19556 5574 19612
rect 5574 19556 5630 19612
rect 5630 19556 5634 19612
rect 5570 19552 5634 19556
rect 14664 19612 14728 19616
rect 14664 19556 14668 19612
rect 14668 19556 14724 19612
rect 14724 19556 14728 19612
rect 14664 19552 14728 19556
rect 14744 19612 14808 19616
rect 14744 19556 14748 19612
rect 14748 19556 14804 19612
rect 14804 19556 14808 19612
rect 14744 19552 14808 19556
rect 14824 19612 14888 19616
rect 14824 19556 14828 19612
rect 14828 19556 14884 19612
rect 14884 19556 14888 19612
rect 14824 19552 14888 19556
rect 14904 19612 14968 19616
rect 14904 19556 14908 19612
rect 14908 19556 14964 19612
rect 14964 19556 14968 19612
rect 14904 19552 14968 19556
rect 23997 19612 24061 19616
rect 23997 19556 24001 19612
rect 24001 19556 24057 19612
rect 24057 19556 24061 19612
rect 23997 19552 24061 19556
rect 24077 19612 24141 19616
rect 24077 19556 24081 19612
rect 24081 19556 24137 19612
rect 24137 19556 24141 19612
rect 24077 19552 24141 19556
rect 24157 19612 24221 19616
rect 24157 19556 24161 19612
rect 24161 19556 24217 19612
rect 24217 19556 24221 19612
rect 24157 19552 24221 19556
rect 24237 19612 24301 19616
rect 24237 19556 24241 19612
rect 24241 19556 24297 19612
rect 24297 19556 24301 19612
rect 24237 19552 24301 19556
rect 23692 19348 23756 19412
rect 9997 19068 10061 19072
rect 9997 19012 10001 19068
rect 10001 19012 10057 19068
rect 10057 19012 10061 19068
rect 9997 19008 10061 19012
rect 10077 19068 10141 19072
rect 10077 19012 10081 19068
rect 10081 19012 10137 19068
rect 10137 19012 10141 19068
rect 10077 19008 10141 19012
rect 10157 19068 10221 19072
rect 10157 19012 10161 19068
rect 10161 19012 10217 19068
rect 10217 19012 10221 19068
rect 10157 19008 10221 19012
rect 10237 19068 10301 19072
rect 10237 19012 10241 19068
rect 10241 19012 10297 19068
rect 10297 19012 10301 19068
rect 10237 19008 10301 19012
rect 19330 19068 19394 19072
rect 19330 19012 19334 19068
rect 19334 19012 19390 19068
rect 19390 19012 19394 19068
rect 19330 19008 19394 19012
rect 19410 19068 19474 19072
rect 19410 19012 19414 19068
rect 19414 19012 19470 19068
rect 19470 19012 19474 19068
rect 19410 19008 19474 19012
rect 19490 19068 19554 19072
rect 19490 19012 19494 19068
rect 19494 19012 19550 19068
rect 19550 19012 19554 19068
rect 19490 19008 19554 19012
rect 19570 19068 19634 19072
rect 19570 19012 19574 19068
rect 19574 19012 19630 19068
rect 19630 19012 19634 19068
rect 19570 19008 19634 19012
rect 5330 18524 5394 18528
rect 5330 18468 5334 18524
rect 5334 18468 5390 18524
rect 5390 18468 5394 18524
rect 5330 18464 5394 18468
rect 5410 18524 5474 18528
rect 5410 18468 5414 18524
rect 5414 18468 5470 18524
rect 5470 18468 5474 18524
rect 5410 18464 5474 18468
rect 5490 18524 5554 18528
rect 5490 18468 5494 18524
rect 5494 18468 5550 18524
rect 5550 18468 5554 18524
rect 5490 18464 5554 18468
rect 5570 18524 5634 18528
rect 5570 18468 5574 18524
rect 5574 18468 5630 18524
rect 5630 18468 5634 18524
rect 5570 18464 5634 18468
rect 14664 18524 14728 18528
rect 14664 18468 14668 18524
rect 14668 18468 14724 18524
rect 14724 18468 14728 18524
rect 14664 18464 14728 18468
rect 14744 18524 14808 18528
rect 14744 18468 14748 18524
rect 14748 18468 14804 18524
rect 14804 18468 14808 18524
rect 14744 18464 14808 18468
rect 14824 18524 14888 18528
rect 14824 18468 14828 18524
rect 14828 18468 14884 18524
rect 14884 18468 14888 18524
rect 14824 18464 14888 18468
rect 14904 18524 14968 18528
rect 14904 18468 14908 18524
rect 14908 18468 14964 18524
rect 14964 18468 14968 18524
rect 14904 18464 14968 18468
rect 23997 18524 24061 18528
rect 23997 18468 24001 18524
rect 24001 18468 24057 18524
rect 24057 18468 24061 18524
rect 23997 18464 24061 18468
rect 24077 18524 24141 18528
rect 24077 18468 24081 18524
rect 24081 18468 24137 18524
rect 24137 18468 24141 18524
rect 24077 18464 24141 18468
rect 24157 18524 24221 18528
rect 24157 18468 24161 18524
rect 24161 18468 24217 18524
rect 24217 18468 24221 18524
rect 24157 18464 24221 18468
rect 24237 18524 24301 18528
rect 24237 18468 24241 18524
rect 24241 18468 24297 18524
rect 24297 18468 24301 18524
rect 24237 18464 24301 18468
rect 9997 17980 10061 17984
rect 9997 17924 10001 17980
rect 10001 17924 10057 17980
rect 10057 17924 10061 17980
rect 9997 17920 10061 17924
rect 10077 17980 10141 17984
rect 10077 17924 10081 17980
rect 10081 17924 10137 17980
rect 10137 17924 10141 17980
rect 10077 17920 10141 17924
rect 10157 17980 10221 17984
rect 10157 17924 10161 17980
rect 10161 17924 10217 17980
rect 10217 17924 10221 17980
rect 10157 17920 10221 17924
rect 10237 17980 10301 17984
rect 10237 17924 10241 17980
rect 10241 17924 10297 17980
rect 10297 17924 10301 17980
rect 10237 17920 10301 17924
rect 19330 17980 19394 17984
rect 19330 17924 19334 17980
rect 19334 17924 19390 17980
rect 19390 17924 19394 17980
rect 19330 17920 19394 17924
rect 19410 17980 19474 17984
rect 19410 17924 19414 17980
rect 19414 17924 19470 17980
rect 19470 17924 19474 17980
rect 19410 17920 19474 17924
rect 19490 17980 19554 17984
rect 19490 17924 19494 17980
rect 19494 17924 19550 17980
rect 19550 17924 19554 17980
rect 19490 17920 19554 17924
rect 19570 17980 19634 17984
rect 19570 17924 19574 17980
rect 19574 17924 19630 17980
rect 19630 17924 19634 17980
rect 19570 17920 19634 17924
rect 5330 17436 5394 17440
rect 5330 17380 5334 17436
rect 5334 17380 5390 17436
rect 5390 17380 5394 17436
rect 5330 17376 5394 17380
rect 5410 17436 5474 17440
rect 5410 17380 5414 17436
rect 5414 17380 5470 17436
rect 5470 17380 5474 17436
rect 5410 17376 5474 17380
rect 5490 17436 5554 17440
rect 5490 17380 5494 17436
rect 5494 17380 5550 17436
rect 5550 17380 5554 17436
rect 5490 17376 5554 17380
rect 5570 17436 5634 17440
rect 5570 17380 5574 17436
rect 5574 17380 5630 17436
rect 5630 17380 5634 17436
rect 5570 17376 5634 17380
rect 14664 17436 14728 17440
rect 14664 17380 14668 17436
rect 14668 17380 14724 17436
rect 14724 17380 14728 17436
rect 14664 17376 14728 17380
rect 14744 17436 14808 17440
rect 14744 17380 14748 17436
rect 14748 17380 14804 17436
rect 14804 17380 14808 17436
rect 14744 17376 14808 17380
rect 14824 17436 14888 17440
rect 14824 17380 14828 17436
rect 14828 17380 14884 17436
rect 14884 17380 14888 17436
rect 14824 17376 14888 17380
rect 14904 17436 14968 17440
rect 14904 17380 14908 17436
rect 14908 17380 14964 17436
rect 14964 17380 14968 17436
rect 14904 17376 14968 17380
rect 23997 17436 24061 17440
rect 23997 17380 24001 17436
rect 24001 17380 24057 17436
rect 24057 17380 24061 17436
rect 23997 17376 24061 17380
rect 24077 17436 24141 17440
rect 24077 17380 24081 17436
rect 24081 17380 24137 17436
rect 24137 17380 24141 17436
rect 24077 17376 24141 17380
rect 24157 17436 24221 17440
rect 24157 17380 24161 17436
rect 24161 17380 24217 17436
rect 24217 17380 24221 17436
rect 24157 17376 24221 17380
rect 24237 17436 24301 17440
rect 24237 17380 24241 17436
rect 24241 17380 24297 17436
rect 24297 17380 24301 17436
rect 24237 17376 24301 17380
rect 9997 16892 10061 16896
rect 9997 16836 10001 16892
rect 10001 16836 10057 16892
rect 10057 16836 10061 16892
rect 9997 16832 10061 16836
rect 10077 16892 10141 16896
rect 10077 16836 10081 16892
rect 10081 16836 10137 16892
rect 10137 16836 10141 16892
rect 10077 16832 10141 16836
rect 10157 16892 10221 16896
rect 10157 16836 10161 16892
rect 10161 16836 10217 16892
rect 10217 16836 10221 16892
rect 10157 16832 10221 16836
rect 10237 16892 10301 16896
rect 10237 16836 10241 16892
rect 10241 16836 10297 16892
rect 10297 16836 10301 16892
rect 10237 16832 10301 16836
rect 19330 16892 19394 16896
rect 19330 16836 19334 16892
rect 19334 16836 19390 16892
rect 19390 16836 19394 16892
rect 19330 16832 19394 16836
rect 19410 16892 19474 16896
rect 19410 16836 19414 16892
rect 19414 16836 19470 16892
rect 19470 16836 19474 16892
rect 19410 16832 19474 16836
rect 19490 16892 19554 16896
rect 19490 16836 19494 16892
rect 19494 16836 19550 16892
rect 19550 16836 19554 16892
rect 19490 16832 19554 16836
rect 19570 16892 19634 16896
rect 19570 16836 19574 16892
rect 19574 16836 19630 16892
rect 19630 16836 19634 16892
rect 19570 16832 19634 16836
rect 5330 16348 5394 16352
rect 5330 16292 5334 16348
rect 5334 16292 5390 16348
rect 5390 16292 5394 16348
rect 5330 16288 5394 16292
rect 5410 16348 5474 16352
rect 5410 16292 5414 16348
rect 5414 16292 5470 16348
rect 5470 16292 5474 16348
rect 5410 16288 5474 16292
rect 5490 16348 5554 16352
rect 5490 16292 5494 16348
rect 5494 16292 5550 16348
rect 5550 16292 5554 16348
rect 5490 16288 5554 16292
rect 5570 16348 5634 16352
rect 5570 16292 5574 16348
rect 5574 16292 5630 16348
rect 5630 16292 5634 16348
rect 5570 16288 5634 16292
rect 14664 16348 14728 16352
rect 14664 16292 14668 16348
rect 14668 16292 14724 16348
rect 14724 16292 14728 16348
rect 14664 16288 14728 16292
rect 14744 16348 14808 16352
rect 14744 16292 14748 16348
rect 14748 16292 14804 16348
rect 14804 16292 14808 16348
rect 14744 16288 14808 16292
rect 14824 16348 14888 16352
rect 14824 16292 14828 16348
rect 14828 16292 14884 16348
rect 14884 16292 14888 16348
rect 14824 16288 14888 16292
rect 14904 16348 14968 16352
rect 14904 16292 14908 16348
rect 14908 16292 14964 16348
rect 14964 16292 14968 16348
rect 14904 16288 14968 16292
rect 23997 16348 24061 16352
rect 23997 16292 24001 16348
rect 24001 16292 24057 16348
rect 24057 16292 24061 16348
rect 23997 16288 24061 16292
rect 24077 16348 24141 16352
rect 24077 16292 24081 16348
rect 24081 16292 24137 16348
rect 24137 16292 24141 16348
rect 24077 16288 24141 16292
rect 24157 16348 24221 16352
rect 24157 16292 24161 16348
rect 24161 16292 24217 16348
rect 24217 16292 24221 16348
rect 24157 16288 24221 16292
rect 24237 16348 24301 16352
rect 24237 16292 24241 16348
rect 24241 16292 24297 16348
rect 24297 16292 24301 16348
rect 24237 16288 24301 16292
rect 9997 15804 10061 15808
rect 9997 15748 10001 15804
rect 10001 15748 10057 15804
rect 10057 15748 10061 15804
rect 9997 15744 10061 15748
rect 10077 15804 10141 15808
rect 10077 15748 10081 15804
rect 10081 15748 10137 15804
rect 10137 15748 10141 15804
rect 10077 15744 10141 15748
rect 10157 15804 10221 15808
rect 10157 15748 10161 15804
rect 10161 15748 10217 15804
rect 10217 15748 10221 15804
rect 10157 15744 10221 15748
rect 10237 15804 10301 15808
rect 10237 15748 10241 15804
rect 10241 15748 10297 15804
rect 10297 15748 10301 15804
rect 10237 15744 10301 15748
rect 19330 15804 19394 15808
rect 19330 15748 19334 15804
rect 19334 15748 19390 15804
rect 19390 15748 19394 15804
rect 19330 15744 19394 15748
rect 19410 15804 19474 15808
rect 19410 15748 19414 15804
rect 19414 15748 19470 15804
rect 19470 15748 19474 15804
rect 19410 15744 19474 15748
rect 19490 15804 19554 15808
rect 19490 15748 19494 15804
rect 19494 15748 19550 15804
rect 19550 15748 19554 15804
rect 19490 15744 19554 15748
rect 19570 15804 19634 15808
rect 19570 15748 19574 15804
rect 19574 15748 19630 15804
rect 19630 15748 19634 15804
rect 19570 15744 19634 15748
rect 5330 15260 5394 15264
rect 5330 15204 5334 15260
rect 5334 15204 5390 15260
rect 5390 15204 5394 15260
rect 5330 15200 5394 15204
rect 5410 15260 5474 15264
rect 5410 15204 5414 15260
rect 5414 15204 5470 15260
rect 5470 15204 5474 15260
rect 5410 15200 5474 15204
rect 5490 15260 5554 15264
rect 5490 15204 5494 15260
rect 5494 15204 5550 15260
rect 5550 15204 5554 15260
rect 5490 15200 5554 15204
rect 5570 15260 5634 15264
rect 5570 15204 5574 15260
rect 5574 15204 5630 15260
rect 5630 15204 5634 15260
rect 5570 15200 5634 15204
rect 14664 15260 14728 15264
rect 14664 15204 14668 15260
rect 14668 15204 14724 15260
rect 14724 15204 14728 15260
rect 14664 15200 14728 15204
rect 14744 15260 14808 15264
rect 14744 15204 14748 15260
rect 14748 15204 14804 15260
rect 14804 15204 14808 15260
rect 14744 15200 14808 15204
rect 14824 15260 14888 15264
rect 14824 15204 14828 15260
rect 14828 15204 14884 15260
rect 14884 15204 14888 15260
rect 14824 15200 14888 15204
rect 14904 15260 14968 15264
rect 14904 15204 14908 15260
rect 14908 15204 14964 15260
rect 14964 15204 14968 15260
rect 14904 15200 14968 15204
rect 23997 15260 24061 15264
rect 23997 15204 24001 15260
rect 24001 15204 24057 15260
rect 24057 15204 24061 15260
rect 23997 15200 24061 15204
rect 24077 15260 24141 15264
rect 24077 15204 24081 15260
rect 24081 15204 24137 15260
rect 24137 15204 24141 15260
rect 24077 15200 24141 15204
rect 24157 15260 24221 15264
rect 24157 15204 24161 15260
rect 24161 15204 24217 15260
rect 24217 15204 24221 15260
rect 24157 15200 24221 15204
rect 24237 15260 24301 15264
rect 24237 15204 24241 15260
rect 24241 15204 24297 15260
rect 24297 15204 24301 15260
rect 24237 15200 24301 15204
rect 9997 14716 10061 14720
rect 9997 14660 10001 14716
rect 10001 14660 10057 14716
rect 10057 14660 10061 14716
rect 9997 14656 10061 14660
rect 10077 14716 10141 14720
rect 10077 14660 10081 14716
rect 10081 14660 10137 14716
rect 10137 14660 10141 14716
rect 10077 14656 10141 14660
rect 10157 14716 10221 14720
rect 10157 14660 10161 14716
rect 10161 14660 10217 14716
rect 10217 14660 10221 14716
rect 10157 14656 10221 14660
rect 10237 14716 10301 14720
rect 10237 14660 10241 14716
rect 10241 14660 10297 14716
rect 10297 14660 10301 14716
rect 10237 14656 10301 14660
rect 19330 14716 19394 14720
rect 19330 14660 19334 14716
rect 19334 14660 19390 14716
rect 19390 14660 19394 14716
rect 19330 14656 19394 14660
rect 19410 14716 19474 14720
rect 19410 14660 19414 14716
rect 19414 14660 19470 14716
rect 19470 14660 19474 14716
rect 19410 14656 19474 14660
rect 19490 14716 19554 14720
rect 19490 14660 19494 14716
rect 19494 14660 19550 14716
rect 19550 14660 19554 14716
rect 19490 14656 19554 14660
rect 19570 14716 19634 14720
rect 19570 14660 19574 14716
rect 19574 14660 19630 14716
rect 19630 14660 19634 14716
rect 19570 14656 19634 14660
rect 5330 14172 5394 14176
rect 5330 14116 5334 14172
rect 5334 14116 5390 14172
rect 5390 14116 5394 14172
rect 5330 14112 5394 14116
rect 5410 14172 5474 14176
rect 5410 14116 5414 14172
rect 5414 14116 5470 14172
rect 5470 14116 5474 14172
rect 5410 14112 5474 14116
rect 5490 14172 5554 14176
rect 5490 14116 5494 14172
rect 5494 14116 5550 14172
rect 5550 14116 5554 14172
rect 5490 14112 5554 14116
rect 5570 14172 5634 14176
rect 5570 14116 5574 14172
rect 5574 14116 5630 14172
rect 5630 14116 5634 14172
rect 5570 14112 5634 14116
rect 14664 14172 14728 14176
rect 14664 14116 14668 14172
rect 14668 14116 14724 14172
rect 14724 14116 14728 14172
rect 14664 14112 14728 14116
rect 14744 14172 14808 14176
rect 14744 14116 14748 14172
rect 14748 14116 14804 14172
rect 14804 14116 14808 14172
rect 14744 14112 14808 14116
rect 14824 14172 14888 14176
rect 14824 14116 14828 14172
rect 14828 14116 14884 14172
rect 14884 14116 14888 14172
rect 14824 14112 14888 14116
rect 14904 14172 14968 14176
rect 14904 14116 14908 14172
rect 14908 14116 14964 14172
rect 14964 14116 14968 14172
rect 14904 14112 14968 14116
rect 23997 14172 24061 14176
rect 23997 14116 24001 14172
rect 24001 14116 24057 14172
rect 24057 14116 24061 14172
rect 23997 14112 24061 14116
rect 24077 14172 24141 14176
rect 24077 14116 24081 14172
rect 24081 14116 24137 14172
rect 24137 14116 24141 14172
rect 24077 14112 24141 14116
rect 24157 14172 24221 14176
rect 24157 14116 24161 14172
rect 24161 14116 24217 14172
rect 24217 14116 24221 14172
rect 24157 14112 24221 14116
rect 24237 14172 24301 14176
rect 24237 14116 24241 14172
rect 24241 14116 24297 14172
rect 24297 14116 24301 14172
rect 24237 14112 24301 14116
rect 9997 13628 10061 13632
rect 9997 13572 10001 13628
rect 10001 13572 10057 13628
rect 10057 13572 10061 13628
rect 9997 13568 10061 13572
rect 10077 13628 10141 13632
rect 10077 13572 10081 13628
rect 10081 13572 10137 13628
rect 10137 13572 10141 13628
rect 10077 13568 10141 13572
rect 10157 13628 10221 13632
rect 10157 13572 10161 13628
rect 10161 13572 10217 13628
rect 10217 13572 10221 13628
rect 10157 13568 10221 13572
rect 10237 13628 10301 13632
rect 10237 13572 10241 13628
rect 10241 13572 10297 13628
rect 10297 13572 10301 13628
rect 10237 13568 10301 13572
rect 19330 13628 19394 13632
rect 19330 13572 19334 13628
rect 19334 13572 19390 13628
rect 19390 13572 19394 13628
rect 19330 13568 19394 13572
rect 19410 13628 19474 13632
rect 19410 13572 19414 13628
rect 19414 13572 19470 13628
rect 19470 13572 19474 13628
rect 19410 13568 19474 13572
rect 19490 13628 19554 13632
rect 19490 13572 19494 13628
rect 19494 13572 19550 13628
rect 19550 13572 19554 13628
rect 19490 13568 19554 13572
rect 19570 13628 19634 13632
rect 19570 13572 19574 13628
rect 19574 13572 19630 13628
rect 19630 13572 19634 13628
rect 19570 13568 19634 13572
rect 5330 13084 5394 13088
rect 5330 13028 5334 13084
rect 5334 13028 5390 13084
rect 5390 13028 5394 13084
rect 5330 13024 5394 13028
rect 5410 13084 5474 13088
rect 5410 13028 5414 13084
rect 5414 13028 5470 13084
rect 5470 13028 5474 13084
rect 5410 13024 5474 13028
rect 5490 13084 5554 13088
rect 5490 13028 5494 13084
rect 5494 13028 5550 13084
rect 5550 13028 5554 13084
rect 5490 13024 5554 13028
rect 5570 13084 5634 13088
rect 5570 13028 5574 13084
rect 5574 13028 5630 13084
rect 5630 13028 5634 13084
rect 5570 13024 5634 13028
rect 14664 13084 14728 13088
rect 14664 13028 14668 13084
rect 14668 13028 14724 13084
rect 14724 13028 14728 13084
rect 14664 13024 14728 13028
rect 14744 13084 14808 13088
rect 14744 13028 14748 13084
rect 14748 13028 14804 13084
rect 14804 13028 14808 13084
rect 14744 13024 14808 13028
rect 14824 13084 14888 13088
rect 14824 13028 14828 13084
rect 14828 13028 14884 13084
rect 14884 13028 14888 13084
rect 14824 13024 14888 13028
rect 14904 13084 14968 13088
rect 14904 13028 14908 13084
rect 14908 13028 14964 13084
rect 14964 13028 14968 13084
rect 14904 13024 14968 13028
rect 23997 13084 24061 13088
rect 23997 13028 24001 13084
rect 24001 13028 24057 13084
rect 24057 13028 24061 13084
rect 23997 13024 24061 13028
rect 24077 13084 24141 13088
rect 24077 13028 24081 13084
rect 24081 13028 24137 13084
rect 24137 13028 24141 13084
rect 24077 13024 24141 13028
rect 24157 13084 24221 13088
rect 24157 13028 24161 13084
rect 24161 13028 24217 13084
rect 24217 13028 24221 13084
rect 24157 13024 24221 13028
rect 24237 13084 24301 13088
rect 24237 13028 24241 13084
rect 24241 13028 24297 13084
rect 24297 13028 24301 13084
rect 24237 13024 24301 13028
rect 9997 12540 10061 12544
rect 9997 12484 10001 12540
rect 10001 12484 10057 12540
rect 10057 12484 10061 12540
rect 9997 12480 10061 12484
rect 10077 12540 10141 12544
rect 10077 12484 10081 12540
rect 10081 12484 10137 12540
rect 10137 12484 10141 12540
rect 10077 12480 10141 12484
rect 10157 12540 10221 12544
rect 10157 12484 10161 12540
rect 10161 12484 10217 12540
rect 10217 12484 10221 12540
rect 10157 12480 10221 12484
rect 10237 12540 10301 12544
rect 10237 12484 10241 12540
rect 10241 12484 10297 12540
rect 10297 12484 10301 12540
rect 10237 12480 10301 12484
rect 19330 12540 19394 12544
rect 19330 12484 19334 12540
rect 19334 12484 19390 12540
rect 19390 12484 19394 12540
rect 19330 12480 19394 12484
rect 19410 12540 19474 12544
rect 19410 12484 19414 12540
rect 19414 12484 19470 12540
rect 19470 12484 19474 12540
rect 19410 12480 19474 12484
rect 19490 12540 19554 12544
rect 19490 12484 19494 12540
rect 19494 12484 19550 12540
rect 19550 12484 19554 12540
rect 19490 12480 19554 12484
rect 19570 12540 19634 12544
rect 19570 12484 19574 12540
rect 19574 12484 19630 12540
rect 19630 12484 19634 12540
rect 19570 12480 19634 12484
rect 5330 11996 5394 12000
rect 5330 11940 5334 11996
rect 5334 11940 5390 11996
rect 5390 11940 5394 11996
rect 5330 11936 5394 11940
rect 5410 11996 5474 12000
rect 5410 11940 5414 11996
rect 5414 11940 5470 11996
rect 5470 11940 5474 11996
rect 5410 11936 5474 11940
rect 5490 11996 5554 12000
rect 5490 11940 5494 11996
rect 5494 11940 5550 11996
rect 5550 11940 5554 11996
rect 5490 11936 5554 11940
rect 5570 11996 5634 12000
rect 5570 11940 5574 11996
rect 5574 11940 5630 11996
rect 5630 11940 5634 11996
rect 5570 11936 5634 11940
rect 14664 11996 14728 12000
rect 14664 11940 14668 11996
rect 14668 11940 14724 11996
rect 14724 11940 14728 11996
rect 14664 11936 14728 11940
rect 14744 11996 14808 12000
rect 14744 11940 14748 11996
rect 14748 11940 14804 11996
rect 14804 11940 14808 11996
rect 14744 11936 14808 11940
rect 14824 11996 14888 12000
rect 14824 11940 14828 11996
rect 14828 11940 14884 11996
rect 14884 11940 14888 11996
rect 14824 11936 14888 11940
rect 14904 11996 14968 12000
rect 14904 11940 14908 11996
rect 14908 11940 14964 11996
rect 14964 11940 14968 11996
rect 14904 11936 14968 11940
rect 23997 11996 24061 12000
rect 23997 11940 24001 11996
rect 24001 11940 24057 11996
rect 24057 11940 24061 11996
rect 23997 11936 24061 11940
rect 24077 11996 24141 12000
rect 24077 11940 24081 11996
rect 24081 11940 24137 11996
rect 24137 11940 24141 11996
rect 24077 11936 24141 11940
rect 24157 11996 24221 12000
rect 24157 11940 24161 11996
rect 24161 11940 24217 11996
rect 24217 11940 24221 11996
rect 24157 11936 24221 11940
rect 24237 11996 24301 12000
rect 24237 11940 24241 11996
rect 24241 11940 24297 11996
rect 24297 11940 24301 11996
rect 24237 11936 24301 11940
rect 9997 11452 10061 11456
rect 9997 11396 10001 11452
rect 10001 11396 10057 11452
rect 10057 11396 10061 11452
rect 9997 11392 10061 11396
rect 10077 11452 10141 11456
rect 10077 11396 10081 11452
rect 10081 11396 10137 11452
rect 10137 11396 10141 11452
rect 10077 11392 10141 11396
rect 10157 11452 10221 11456
rect 10157 11396 10161 11452
rect 10161 11396 10217 11452
rect 10217 11396 10221 11452
rect 10157 11392 10221 11396
rect 10237 11452 10301 11456
rect 10237 11396 10241 11452
rect 10241 11396 10297 11452
rect 10297 11396 10301 11452
rect 10237 11392 10301 11396
rect 19330 11452 19394 11456
rect 19330 11396 19334 11452
rect 19334 11396 19390 11452
rect 19390 11396 19394 11452
rect 19330 11392 19394 11396
rect 19410 11452 19474 11456
rect 19410 11396 19414 11452
rect 19414 11396 19470 11452
rect 19470 11396 19474 11452
rect 19410 11392 19474 11396
rect 19490 11452 19554 11456
rect 19490 11396 19494 11452
rect 19494 11396 19550 11452
rect 19550 11396 19554 11452
rect 19490 11392 19554 11396
rect 19570 11452 19634 11456
rect 19570 11396 19574 11452
rect 19574 11396 19630 11452
rect 19630 11396 19634 11452
rect 19570 11392 19634 11396
rect 5330 10908 5394 10912
rect 5330 10852 5334 10908
rect 5334 10852 5390 10908
rect 5390 10852 5394 10908
rect 5330 10848 5394 10852
rect 5410 10908 5474 10912
rect 5410 10852 5414 10908
rect 5414 10852 5470 10908
rect 5470 10852 5474 10908
rect 5410 10848 5474 10852
rect 5490 10908 5554 10912
rect 5490 10852 5494 10908
rect 5494 10852 5550 10908
rect 5550 10852 5554 10908
rect 5490 10848 5554 10852
rect 5570 10908 5634 10912
rect 5570 10852 5574 10908
rect 5574 10852 5630 10908
rect 5630 10852 5634 10908
rect 5570 10848 5634 10852
rect 14664 10908 14728 10912
rect 14664 10852 14668 10908
rect 14668 10852 14724 10908
rect 14724 10852 14728 10908
rect 14664 10848 14728 10852
rect 14744 10908 14808 10912
rect 14744 10852 14748 10908
rect 14748 10852 14804 10908
rect 14804 10852 14808 10908
rect 14744 10848 14808 10852
rect 14824 10908 14888 10912
rect 14824 10852 14828 10908
rect 14828 10852 14884 10908
rect 14884 10852 14888 10908
rect 14824 10848 14888 10852
rect 14904 10908 14968 10912
rect 14904 10852 14908 10908
rect 14908 10852 14964 10908
rect 14964 10852 14968 10908
rect 14904 10848 14968 10852
rect 23997 10908 24061 10912
rect 23997 10852 24001 10908
rect 24001 10852 24057 10908
rect 24057 10852 24061 10908
rect 23997 10848 24061 10852
rect 24077 10908 24141 10912
rect 24077 10852 24081 10908
rect 24081 10852 24137 10908
rect 24137 10852 24141 10908
rect 24077 10848 24141 10852
rect 24157 10908 24221 10912
rect 24157 10852 24161 10908
rect 24161 10852 24217 10908
rect 24217 10852 24221 10908
rect 24157 10848 24221 10852
rect 24237 10908 24301 10912
rect 24237 10852 24241 10908
rect 24241 10852 24297 10908
rect 24297 10852 24301 10908
rect 24237 10848 24301 10852
rect 9997 10364 10061 10368
rect 9997 10308 10001 10364
rect 10001 10308 10057 10364
rect 10057 10308 10061 10364
rect 9997 10304 10061 10308
rect 10077 10364 10141 10368
rect 10077 10308 10081 10364
rect 10081 10308 10137 10364
rect 10137 10308 10141 10364
rect 10077 10304 10141 10308
rect 10157 10364 10221 10368
rect 10157 10308 10161 10364
rect 10161 10308 10217 10364
rect 10217 10308 10221 10364
rect 10157 10304 10221 10308
rect 10237 10364 10301 10368
rect 10237 10308 10241 10364
rect 10241 10308 10297 10364
rect 10297 10308 10301 10364
rect 10237 10304 10301 10308
rect 19330 10364 19394 10368
rect 19330 10308 19334 10364
rect 19334 10308 19390 10364
rect 19390 10308 19394 10364
rect 19330 10304 19394 10308
rect 19410 10364 19474 10368
rect 19410 10308 19414 10364
rect 19414 10308 19470 10364
rect 19470 10308 19474 10364
rect 19410 10304 19474 10308
rect 19490 10364 19554 10368
rect 19490 10308 19494 10364
rect 19494 10308 19550 10364
rect 19550 10308 19554 10364
rect 19490 10304 19554 10308
rect 19570 10364 19634 10368
rect 19570 10308 19574 10364
rect 19574 10308 19630 10364
rect 19630 10308 19634 10364
rect 19570 10304 19634 10308
rect 5330 9820 5394 9824
rect 5330 9764 5334 9820
rect 5334 9764 5390 9820
rect 5390 9764 5394 9820
rect 5330 9760 5394 9764
rect 5410 9820 5474 9824
rect 5410 9764 5414 9820
rect 5414 9764 5470 9820
rect 5470 9764 5474 9820
rect 5410 9760 5474 9764
rect 5490 9820 5554 9824
rect 5490 9764 5494 9820
rect 5494 9764 5550 9820
rect 5550 9764 5554 9820
rect 5490 9760 5554 9764
rect 5570 9820 5634 9824
rect 5570 9764 5574 9820
rect 5574 9764 5630 9820
rect 5630 9764 5634 9820
rect 5570 9760 5634 9764
rect 14664 9820 14728 9824
rect 14664 9764 14668 9820
rect 14668 9764 14724 9820
rect 14724 9764 14728 9820
rect 14664 9760 14728 9764
rect 14744 9820 14808 9824
rect 14744 9764 14748 9820
rect 14748 9764 14804 9820
rect 14804 9764 14808 9820
rect 14744 9760 14808 9764
rect 14824 9820 14888 9824
rect 14824 9764 14828 9820
rect 14828 9764 14884 9820
rect 14884 9764 14888 9820
rect 14824 9760 14888 9764
rect 14904 9820 14968 9824
rect 14904 9764 14908 9820
rect 14908 9764 14964 9820
rect 14964 9764 14968 9820
rect 14904 9760 14968 9764
rect 23997 9820 24061 9824
rect 23997 9764 24001 9820
rect 24001 9764 24057 9820
rect 24057 9764 24061 9820
rect 23997 9760 24061 9764
rect 24077 9820 24141 9824
rect 24077 9764 24081 9820
rect 24081 9764 24137 9820
rect 24137 9764 24141 9820
rect 24077 9760 24141 9764
rect 24157 9820 24221 9824
rect 24157 9764 24161 9820
rect 24161 9764 24217 9820
rect 24217 9764 24221 9820
rect 24157 9760 24221 9764
rect 24237 9820 24301 9824
rect 24237 9764 24241 9820
rect 24241 9764 24297 9820
rect 24297 9764 24301 9820
rect 24237 9760 24301 9764
rect 9997 9276 10061 9280
rect 9997 9220 10001 9276
rect 10001 9220 10057 9276
rect 10057 9220 10061 9276
rect 9997 9216 10061 9220
rect 10077 9276 10141 9280
rect 10077 9220 10081 9276
rect 10081 9220 10137 9276
rect 10137 9220 10141 9276
rect 10077 9216 10141 9220
rect 10157 9276 10221 9280
rect 10157 9220 10161 9276
rect 10161 9220 10217 9276
rect 10217 9220 10221 9276
rect 10157 9216 10221 9220
rect 10237 9276 10301 9280
rect 10237 9220 10241 9276
rect 10241 9220 10297 9276
rect 10297 9220 10301 9276
rect 10237 9216 10301 9220
rect 19330 9276 19394 9280
rect 19330 9220 19334 9276
rect 19334 9220 19390 9276
rect 19390 9220 19394 9276
rect 19330 9216 19394 9220
rect 19410 9276 19474 9280
rect 19410 9220 19414 9276
rect 19414 9220 19470 9276
rect 19470 9220 19474 9276
rect 19410 9216 19474 9220
rect 19490 9276 19554 9280
rect 19490 9220 19494 9276
rect 19494 9220 19550 9276
rect 19550 9220 19554 9276
rect 19490 9216 19554 9220
rect 19570 9276 19634 9280
rect 19570 9220 19574 9276
rect 19574 9220 19630 9276
rect 19630 9220 19634 9276
rect 19570 9216 19634 9220
rect 5330 8732 5394 8736
rect 5330 8676 5334 8732
rect 5334 8676 5390 8732
rect 5390 8676 5394 8732
rect 5330 8672 5394 8676
rect 5410 8732 5474 8736
rect 5410 8676 5414 8732
rect 5414 8676 5470 8732
rect 5470 8676 5474 8732
rect 5410 8672 5474 8676
rect 5490 8732 5554 8736
rect 5490 8676 5494 8732
rect 5494 8676 5550 8732
rect 5550 8676 5554 8732
rect 5490 8672 5554 8676
rect 5570 8732 5634 8736
rect 5570 8676 5574 8732
rect 5574 8676 5630 8732
rect 5630 8676 5634 8732
rect 5570 8672 5634 8676
rect 14664 8732 14728 8736
rect 14664 8676 14668 8732
rect 14668 8676 14724 8732
rect 14724 8676 14728 8732
rect 14664 8672 14728 8676
rect 14744 8732 14808 8736
rect 14744 8676 14748 8732
rect 14748 8676 14804 8732
rect 14804 8676 14808 8732
rect 14744 8672 14808 8676
rect 14824 8732 14888 8736
rect 14824 8676 14828 8732
rect 14828 8676 14884 8732
rect 14884 8676 14888 8732
rect 14824 8672 14888 8676
rect 14904 8732 14968 8736
rect 14904 8676 14908 8732
rect 14908 8676 14964 8732
rect 14964 8676 14968 8732
rect 14904 8672 14968 8676
rect 23997 8732 24061 8736
rect 23997 8676 24001 8732
rect 24001 8676 24057 8732
rect 24057 8676 24061 8732
rect 23997 8672 24061 8676
rect 24077 8732 24141 8736
rect 24077 8676 24081 8732
rect 24081 8676 24137 8732
rect 24137 8676 24141 8732
rect 24077 8672 24141 8676
rect 24157 8732 24221 8736
rect 24157 8676 24161 8732
rect 24161 8676 24217 8732
rect 24217 8676 24221 8732
rect 24157 8672 24221 8676
rect 24237 8732 24301 8736
rect 24237 8676 24241 8732
rect 24241 8676 24297 8732
rect 24297 8676 24301 8732
rect 24237 8672 24301 8676
rect 9997 8188 10061 8192
rect 9997 8132 10001 8188
rect 10001 8132 10057 8188
rect 10057 8132 10061 8188
rect 9997 8128 10061 8132
rect 10077 8188 10141 8192
rect 10077 8132 10081 8188
rect 10081 8132 10137 8188
rect 10137 8132 10141 8188
rect 10077 8128 10141 8132
rect 10157 8188 10221 8192
rect 10157 8132 10161 8188
rect 10161 8132 10217 8188
rect 10217 8132 10221 8188
rect 10157 8128 10221 8132
rect 10237 8188 10301 8192
rect 10237 8132 10241 8188
rect 10241 8132 10297 8188
rect 10297 8132 10301 8188
rect 10237 8128 10301 8132
rect 19330 8188 19394 8192
rect 19330 8132 19334 8188
rect 19334 8132 19390 8188
rect 19390 8132 19394 8188
rect 19330 8128 19394 8132
rect 19410 8188 19474 8192
rect 19410 8132 19414 8188
rect 19414 8132 19470 8188
rect 19470 8132 19474 8188
rect 19410 8128 19474 8132
rect 19490 8188 19554 8192
rect 19490 8132 19494 8188
rect 19494 8132 19550 8188
rect 19550 8132 19554 8188
rect 19490 8128 19554 8132
rect 19570 8188 19634 8192
rect 19570 8132 19574 8188
rect 19574 8132 19630 8188
rect 19630 8132 19634 8188
rect 19570 8128 19634 8132
rect 5330 7644 5394 7648
rect 5330 7588 5334 7644
rect 5334 7588 5390 7644
rect 5390 7588 5394 7644
rect 5330 7584 5394 7588
rect 5410 7644 5474 7648
rect 5410 7588 5414 7644
rect 5414 7588 5470 7644
rect 5470 7588 5474 7644
rect 5410 7584 5474 7588
rect 5490 7644 5554 7648
rect 5490 7588 5494 7644
rect 5494 7588 5550 7644
rect 5550 7588 5554 7644
rect 5490 7584 5554 7588
rect 5570 7644 5634 7648
rect 5570 7588 5574 7644
rect 5574 7588 5630 7644
rect 5630 7588 5634 7644
rect 5570 7584 5634 7588
rect 14664 7644 14728 7648
rect 14664 7588 14668 7644
rect 14668 7588 14724 7644
rect 14724 7588 14728 7644
rect 14664 7584 14728 7588
rect 14744 7644 14808 7648
rect 14744 7588 14748 7644
rect 14748 7588 14804 7644
rect 14804 7588 14808 7644
rect 14744 7584 14808 7588
rect 14824 7644 14888 7648
rect 14824 7588 14828 7644
rect 14828 7588 14884 7644
rect 14884 7588 14888 7644
rect 14824 7584 14888 7588
rect 14904 7644 14968 7648
rect 14904 7588 14908 7644
rect 14908 7588 14964 7644
rect 14964 7588 14968 7644
rect 14904 7584 14968 7588
rect 23997 7644 24061 7648
rect 23997 7588 24001 7644
rect 24001 7588 24057 7644
rect 24057 7588 24061 7644
rect 23997 7584 24061 7588
rect 24077 7644 24141 7648
rect 24077 7588 24081 7644
rect 24081 7588 24137 7644
rect 24137 7588 24141 7644
rect 24077 7584 24141 7588
rect 24157 7644 24221 7648
rect 24157 7588 24161 7644
rect 24161 7588 24217 7644
rect 24217 7588 24221 7644
rect 24157 7584 24221 7588
rect 24237 7644 24301 7648
rect 24237 7588 24241 7644
rect 24241 7588 24297 7644
rect 24297 7588 24301 7644
rect 24237 7584 24301 7588
rect 9997 7100 10061 7104
rect 9997 7044 10001 7100
rect 10001 7044 10057 7100
rect 10057 7044 10061 7100
rect 9997 7040 10061 7044
rect 10077 7100 10141 7104
rect 10077 7044 10081 7100
rect 10081 7044 10137 7100
rect 10137 7044 10141 7100
rect 10077 7040 10141 7044
rect 10157 7100 10221 7104
rect 10157 7044 10161 7100
rect 10161 7044 10217 7100
rect 10217 7044 10221 7100
rect 10157 7040 10221 7044
rect 10237 7100 10301 7104
rect 10237 7044 10241 7100
rect 10241 7044 10297 7100
rect 10297 7044 10301 7100
rect 10237 7040 10301 7044
rect 19330 7100 19394 7104
rect 19330 7044 19334 7100
rect 19334 7044 19390 7100
rect 19390 7044 19394 7100
rect 19330 7040 19394 7044
rect 19410 7100 19474 7104
rect 19410 7044 19414 7100
rect 19414 7044 19470 7100
rect 19470 7044 19474 7100
rect 19410 7040 19474 7044
rect 19490 7100 19554 7104
rect 19490 7044 19494 7100
rect 19494 7044 19550 7100
rect 19550 7044 19554 7100
rect 19490 7040 19554 7044
rect 19570 7100 19634 7104
rect 19570 7044 19574 7100
rect 19574 7044 19630 7100
rect 19630 7044 19634 7100
rect 19570 7040 19634 7044
rect 5330 6556 5394 6560
rect 5330 6500 5334 6556
rect 5334 6500 5390 6556
rect 5390 6500 5394 6556
rect 5330 6496 5394 6500
rect 5410 6556 5474 6560
rect 5410 6500 5414 6556
rect 5414 6500 5470 6556
rect 5470 6500 5474 6556
rect 5410 6496 5474 6500
rect 5490 6556 5554 6560
rect 5490 6500 5494 6556
rect 5494 6500 5550 6556
rect 5550 6500 5554 6556
rect 5490 6496 5554 6500
rect 5570 6556 5634 6560
rect 5570 6500 5574 6556
rect 5574 6500 5630 6556
rect 5630 6500 5634 6556
rect 5570 6496 5634 6500
rect 14664 6556 14728 6560
rect 14664 6500 14668 6556
rect 14668 6500 14724 6556
rect 14724 6500 14728 6556
rect 14664 6496 14728 6500
rect 14744 6556 14808 6560
rect 14744 6500 14748 6556
rect 14748 6500 14804 6556
rect 14804 6500 14808 6556
rect 14744 6496 14808 6500
rect 14824 6556 14888 6560
rect 14824 6500 14828 6556
rect 14828 6500 14884 6556
rect 14884 6500 14888 6556
rect 14824 6496 14888 6500
rect 14904 6556 14968 6560
rect 14904 6500 14908 6556
rect 14908 6500 14964 6556
rect 14964 6500 14968 6556
rect 14904 6496 14968 6500
rect 23997 6556 24061 6560
rect 23997 6500 24001 6556
rect 24001 6500 24057 6556
rect 24057 6500 24061 6556
rect 23997 6496 24061 6500
rect 24077 6556 24141 6560
rect 24077 6500 24081 6556
rect 24081 6500 24137 6556
rect 24137 6500 24141 6556
rect 24077 6496 24141 6500
rect 24157 6556 24221 6560
rect 24157 6500 24161 6556
rect 24161 6500 24217 6556
rect 24217 6500 24221 6556
rect 24157 6496 24221 6500
rect 24237 6556 24301 6560
rect 24237 6500 24241 6556
rect 24241 6500 24297 6556
rect 24297 6500 24301 6556
rect 24237 6496 24301 6500
rect 9997 6012 10061 6016
rect 9997 5956 10001 6012
rect 10001 5956 10057 6012
rect 10057 5956 10061 6012
rect 9997 5952 10061 5956
rect 10077 6012 10141 6016
rect 10077 5956 10081 6012
rect 10081 5956 10137 6012
rect 10137 5956 10141 6012
rect 10077 5952 10141 5956
rect 10157 6012 10221 6016
rect 10157 5956 10161 6012
rect 10161 5956 10217 6012
rect 10217 5956 10221 6012
rect 10157 5952 10221 5956
rect 10237 6012 10301 6016
rect 10237 5956 10241 6012
rect 10241 5956 10297 6012
rect 10297 5956 10301 6012
rect 10237 5952 10301 5956
rect 19330 6012 19394 6016
rect 19330 5956 19334 6012
rect 19334 5956 19390 6012
rect 19390 5956 19394 6012
rect 19330 5952 19394 5956
rect 19410 6012 19474 6016
rect 19410 5956 19414 6012
rect 19414 5956 19470 6012
rect 19470 5956 19474 6012
rect 19410 5952 19474 5956
rect 19490 6012 19554 6016
rect 19490 5956 19494 6012
rect 19494 5956 19550 6012
rect 19550 5956 19554 6012
rect 19490 5952 19554 5956
rect 19570 6012 19634 6016
rect 19570 5956 19574 6012
rect 19574 5956 19630 6012
rect 19630 5956 19634 6012
rect 19570 5952 19634 5956
rect 5330 5468 5394 5472
rect 5330 5412 5334 5468
rect 5334 5412 5390 5468
rect 5390 5412 5394 5468
rect 5330 5408 5394 5412
rect 5410 5468 5474 5472
rect 5410 5412 5414 5468
rect 5414 5412 5470 5468
rect 5470 5412 5474 5468
rect 5410 5408 5474 5412
rect 5490 5468 5554 5472
rect 5490 5412 5494 5468
rect 5494 5412 5550 5468
rect 5550 5412 5554 5468
rect 5490 5408 5554 5412
rect 5570 5468 5634 5472
rect 5570 5412 5574 5468
rect 5574 5412 5630 5468
rect 5630 5412 5634 5468
rect 5570 5408 5634 5412
rect 14664 5468 14728 5472
rect 14664 5412 14668 5468
rect 14668 5412 14724 5468
rect 14724 5412 14728 5468
rect 14664 5408 14728 5412
rect 14744 5468 14808 5472
rect 14744 5412 14748 5468
rect 14748 5412 14804 5468
rect 14804 5412 14808 5468
rect 14744 5408 14808 5412
rect 14824 5468 14888 5472
rect 14824 5412 14828 5468
rect 14828 5412 14884 5468
rect 14884 5412 14888 5468
rect 14824 5408 14888 5412
rect 14904 5468 14968 5472
rect 14904 5412 14908 5468
rect 14908 5412 14964 5468
rect 14964 5412 14968 5468
rect 14904 5408 14968 5412
rect 23997 5468 24061 5472
rect 23997 5412 24001 5468
rect 24001 5412 24057 5468
rect 24057 5412 24061 5468
rect 23997 5408 24061 5412
rect 24077 5468 24141 5472
rect 24077 5412 24081 5468
rect 24081 5412 24137 5468
rect 24137 5412 24141 5468
rect 24077 5408 24141 5412
rect 24157 5468 24221 5472
rect 24157 5412 24161 5468
rect 24161 5412 24217 5468
rect 24217 5412 24221 5468
rect 24157 5408 24221 5412
rect 24237 5468 24301 5472
rect 24237 5412 24241 5468
rect 24241 5412 24297 5468
rect 24297 5412 24301 5468
rect 24237 5408 24301 5412
rect 9997 4924 10061 4928
rect 9997 4868 10001 4924
rect 10001 4868 10057 4924
rect 10057 4868 10061 4924
rect 9997 4864 10061 4868
rect 10077 4924 10141 4928
rect 10077 4868 10081 4924
rect 10081 4868 10137 4924
rect 10137 4868 10141 4924
rect 10077 4864 10141 4868
rect 10157 4924 10221 4928
rect 10157 4868 10161 4924
rect 10161 4868 10217 4924
rect 10217 4868 10221 4924
rect 10157 4864 10221 4868
rect 10237 4924 10301 4928
rect 10237 4868 10241 4924
rect 10241 4868 10297 4924
rect 10297 4868 10301 4924
rect 10237 4864 10301 4868
rect 19330 4924 19394 4928
rect 19330 4868 19334 4924
rect 19334 4868 19390 4924
rect 19390 4868 19394 4924
rect 19330 4864 19394 4868
rect 19410 4924 19474 4928
rect 19410 4868 19414 4924
rect 19414 4868 19470 4924
rect 19470 4868 19474 4924
rect 19410 4864 19474 4868
rect 19490 4924 19554 4928
rect 19490 4868 19494 4924
rect 19494 4868 19550 4924
rect 19550 4868 19554 4924
rect 19490 4864 19554 4868
rect 19570 4924 19634 4928
rect 19570 4868 19574 4924
rect 19574 4868 19630 4924
rect 19630 4868 19634 4924
rect 19570 4864 19634 4868
rect 5330 4380 5394 4384
rect 5330 4324 5334 4380
rect 5334 4324 5390 4380
rect 5390 4324 5394 4380
rect 5330 4320 5394 4324
rect 5410 4380 5474 4384
rect 5410 4324 5414 4380
rect 5414 4324 5470 4380
rect 5470 4324 5474 4380
rect 5410 4320 5474 4324
rect 5490 4380 5554 4384
rect 5490 4324 5494 4380
rect 5494 4324 5550 4380
rect 5550 4324 5554 4380
rect 5490 4320 5554 4324
rect 5570 4380 5634 4384
rect 5570 4324 5574 4380
rect 5574 4324 5630 4380
rect 5630 4324 5634 4380
rect 5570 4320 5634 4324
rect 14664 4380 14728 4384
rect 14664 4324 14668 4380
rect 14668 4324 14724 4380
rect 14724 4324 14728 4380
rect 14664 4320 14728 4324
rect 14744 4380 14808 4384
rect 14744 4324 14748 4380
rect 14748 4324 14804 4380
rect 14804 4324 14808 4380
rect 14744 4320 14808 4324
rect 14824 4380 14888 4384
rect 14824 4324 14828 4380
rect 14828 4324 14884 4380
rect 14884 4324 14888 4380
rect 14824 4320 14888 4324
rect 14904 4380 14968 4384
rect 14904 4324 14908 4380
rect 14908 4324 14964 4380
rect 14964 4324 14968 4380
rect 14904 4320 14968 4324
rect 23997 4380 24061 4384
rect 23997 4324 24001 4380
rect 24001 4324 24057 4380
rect 24057 4324 24061 4380
rect 23997 4320 24061 4324
rect 24077 4380 24141 4384
rect 24077 4324 24081 4380
rect 24081 4324 24137 4380
rect 24137 4324 24141 4380
rect 24077 4320 24141 4324
rect 24157 4380 24221 4384
rect 24157 4324 24161 4380
rect 24161 4324 24217 4380
rect 24217 4324 24221 4380
rect 24157 4320 24221 4324
rect 24237 4380 24301 4384
rect 24237 4324 24241 4380
rect 24241 4324 24297 4380
rect 24297 4324 24301 4380
rect 24237 4320 24301 4324
rect 9997 3836 10061 3840
rect 9997 3780 10001 3836
rect 10001 3780 10057 3836
rect 10057 3780 10061 3836
rect 9997 3776 10061 3780
rect 10077 3836 10141 3840
rect 10077 3780 10081 3836
rect 10081 3780 10137 3836
rect 10137 3780 10141 3836
rect 10077 3776 10141 3780
rect 10157 3836 10221 3840
rect 10157 3780 10161 3836
rect 10161 3780 10217 3836
rect 10217 3780 10221 3836
rect 10157 3776 10221 3780
rect 10237 3836 10301 3840
rect 10237 3780 10241 3836
rect 10241 3780 10297 3836
rect 10297 3780 10301 3836
rect 10237 3776 10301 3780
rect 19330 3836 19394 3840
rect 19330 3780 19334 3836
rect 19334 3780 19390 3836
rect 19390 3780 19394 3836
rect 19330 3776 19394 3780
rect 19410 3836 19474 3840
rect 19410 3780 19414 3836
rect 19414 3780 19470 3836
rect 19470 3780 19474 3836
rect 19410 3776 19474 3780
rect 19490 3836 19554 3840
rect 19490 3780 19494 3836
rect 19494 3780 19550 3836
rect 19550 3780 19554 3836
rect 19490 3776 19554 3780
rect 19570 3836 19634 3840
rect 19570 3780 19574 3836
rect 19574 3780 19630 3836
rect 19630 3780 19634 3836
rect 19570 3776 19634 3780
rect 11548 3708 11612 3772
rect 5330 3292 5394 3296
rect 5330 3236 5334 3292
rect 5334 3236 5390 3292
rect 5390 3236 5394 3292
rect 5330 3232 5394 3236
rect 5410 3292 5474 3296
rect 5410 3236 5414 3292
rect 5414 3236 5470 3292
rect 5470 3236 5474 3292
rect 5410 3232 5474 3236
rect 5490 3292 5554 3296
rect 5490 3236 5494 3292
rect 5494 3236 5550 3292
rect 5550 3236 5554 3292
rect 5490 3232 5554 3236
rect 5570 3292 5634 3296
rect 5570 3236 5574 3292
rect 5574 3236 5630 3292
rect 5630 3236 5634 3292
rect 5570 3232 5634 3236
rect 14664 3292 14728 3296
rect 14664 3236 14668 3292
rect 14668 3236 14724 3292
rect 14724 3236 14728 3292
rect 14664 3232 14728 3236
rect 14744 3292 14808 3296
rect 14744 3236 14748 3292
rect 14748 3236 14804 3292
rect 14804 3236 14808 3292
rect 14744 3232 14808 3236
rect 14824 3292 14888 3296
rect 14824 3236 14828 3292
rect 14828 3236 14884 3292
rect 14884 3236 14888 3292
rect 14824 3232 14888 3236
rect 14904 3292 14968 3296
rect 14904 3236 14908 3292
rect 14908 3236 14964 3292
rect 14964 3236 14968 3292
rect 14904 3232 14968 3236
rect 23997 3292 24061 3296
rect 23997 3236 24001 3292
rect 24001 3236 24057 3292
rect 24057 3236 24061 3292
rect 23997 3232 24061 3236
rect 24077 3292 24141 3296
rect 24077 3236 24081 3292
rect 24081 3236 24137 3292
rect 24137 3236 24141 3292
rect 24077 3232 24141 3236
rect 24157 3292 24221 3296
rect 24157 3236 24161 3292
rect 24161 3236 24217 3292
rect 24217 3236 24221 3292
rect 24157 3232 24221 3236
rect 24237 3292 24301 3296
rect 24237 3236 24241 3292
rect 24241 3236 24297 3292
rect 24297 3236 24301 3292
rect 24237 3232 24301 3236
rect 24612 2952 24676 2956
rect 24612 2896 24662 2952
rect 24662 2896 24676 2952
rect 24612 2892 24676 2896
rect 9997 2748 10061 2752
rect 9997 2692 10001 2748
rect 10001 2692 10057 2748
rect 10057 2692 10061 2748
rect 9997 2688 10061 2692
rect 10077 2748 10141 2752
rect 10077 2692 10081 2748
rect 10081 2692 10137 2748
rect 10137 2692 10141 2748
rect 10077 2688 10141 2692
rect 10157 2748 10221 2752
rect 10157 2692 10161 2748
rect 10161 2692 10217 2748
rect 10217 2692 10221 2748
rect 10157 2688 10221 2692
rect 10237 2748 10301 2752
rect 10237 2692 10241 2748
rect 10241 2692 10297 2748
rect 10297 2692 10301 2748
rect 10237 2688 10301 2692
rect 19330 2748 19394 2752
rect 19330 2692 19334 2748
rect 19334 2692 19390 2748
rect 19390 2692 19394 2748
rect 19330 2688 19394 2692
rect 19410 2748 19474 2752
rect 19410 2692 19414 2748
rect 19414 2692 19470 2748
rect 19470 2692 19474 2748
rect 19410 2688 19474 2692
rect 19490 2748 19554 2752
rect 19490 2692 19494 2748
rect 19494 2692 19550 2748
rect 19550 2692 19554 2748
rect 19490 2688 19554 2692
rect 19570 2748 19634 2752
rect 19570 2692 19574 2748
rect 19574 2692 19630 2748
rect 19630 2692 19634 2748
rect 19570 2688 19634 2692
rect 5330 2204 5394 2208
rect 5330 2148 5334 2204
rect 5334 2148 5390 2204
rect 5390 2148 5394 2204
rect 5330 2144 5394 2148
rect 5410 2204 5474 2208
rect 5410 2148 5414 2204
rect 5414 2148 5470 2204
rect 5470 2148 5474 2204
rect 5410 2144 5474 2148
rect 5490 2204 5554 2208
rect 5490 2148 5494 2204
rect 5494 2148 5550 2204
rect 5550 2148 5554 2204
rect 5490 2144 5554 2148
rect 5570 2204 5634 2208
rect 5570 2148 5574 2204
rect 5574 2148 5630 2204
rect 5630 2148 5634 2204
rect 5570 2144 5634 2148
rect 14664 2204 14728 2208
rect 14664 2148 14668 2204
rect 14668 2148 14724 2204
rect 14724 2148 14728 2204
rect 14664 2144 14728 2148
rect 14744 2204 14808 2208
rect 14744 2148 14748 2204
rect 14748 2148 14804 2204
rect 14804 2148 14808 2204
rect 14744 2144 14808 2148
rect 14824 2204 14888 2208
rect 14824 2148 14828 2204
rect 14828 2148 14884 2204
rect 14884 2148 14888 2204
rect 14824 2144 14888 2148
rect 14904 2204 14968 2208
rect 14904 2148 14908 2204
rect 14908 2148 14964 2204
rect 14964 2148 14968 2204
rect 14904 2144 14968 2148
rect 23997 2204 24061 2208
rect 23997 2148 24001 2204
rect 24001 2148 24057 2204
rect 24057 2148 24061 2204
rect 23997 2144 24061 2148
rect 24077 2204 24141 2208
rect 24077 2148 24081 2204
rect 24081 2148 24137 2204
rect 24137 2148 24141 2204
rect 24077 2144 24141 2148
rect 24157 2204 24221 2208
rect 24157 2148 24161 2204
rect 24161 2148 24217 2204
rect 24217 2148 24221 2204
rect 24157 2144 24221 2148
rect 24237 2204 24301 2208
rect 24237 2148 24241 2204
rect 24241 2148 24297 2204
rect 24297 2148 24301 2204
rect 24237 2144 24301 2148
<< metal4 >>
rect 23691 27708 23757 27709
rect 23691 27644 23692 27708
rect 23756 27644 23757 27708
rect 23691 27643 23757 27644
rect 5322 25056 5643 25616
rect 5322 24992 5330 25056
rect 5394 24992 5410 25056
rect 5474 24992 5490 25056
rect 5554 24992 5570 25056
rect 5634 24992 5643 25056
rect 5322 23968 5643 24992
rect 5322 23904 5330 23968
rect 5394 23904 5410 23968
rect 5474 23904 5490 23968
rect 5554 23904 5570 23968
rect 5634 23904 5643 23968
rect 5322 22880 5643 23904
rect 5322 22816 5330 22880
rect 5394 22816 5410 22880
rect 5474 22816 5490 22880
rect 5554 22816 5570 22880
rect 5634 22816 5643 22880
rect 5322 21792 5643 22816
rect 5322 21728 5330 21792
rect 5394 21728 5410 21792
rect 5474 21728 5490 21792
rect 5554 21728 5570 21792
rect 5634 21728 5643 21792
rect 5322 20704 5643 21728
rect 5322 20640 5330 20704
rect 5394 20640 5410 20704
rect 5474 20640 5490 20704
rect 5554 20640 5570 20704
rect 5634 20640 5643 20704
rect 5322 19616 5643 20640
rect 5322 19552 5330 19616
rect 5394 19552 5410 19616
rect 5474 19552 5490 19616
rect 5554 19552 5570 19616
rect 5634 19552 5643 19616
rect 5322 18528 5643 19552
rect 5322 18464 5330 18528
rect 5394 18464 5410 18528
rect 5474 18464 5490 18528
rect 5554 18464 5570 18528
rect 5634 18464 5643 18528
rect 5322 17440 5643 18464
rect 5322 17376 5330 17440
rect 5394 17376 5410 17440
rect 5474 17376 5490 17440
rect 5554 17376 5570 17440
rect 5634 17376 5643 17440
rect 5322 16352 5643 17376
rect 5322 16288 5330 16352
rect 5394 16288 5410 16352
rect 5474 16288 5490 16352
rect 5554 16288 5570 16352
rect 5634 16288 5643 16352
rect 5322 15264 5643 16288
rect 5322 15200 5330 15264
rect 5394 15200 5410 15264
rect 5474 15200 5490 15264
rect 5554 15200 5570 15264
rect 5634 15200 5643 15264
rect 5322 14176 5643 15200
rect 5322 14112 5330 14176
rect 5394 14112 5410 14176
rect 5474 14112 5490 14176
rect 5554 14112 5570 14176
rect 5634 14112 5643 14176
rect 5322 13088 5643 14112
rect 5322 13024 5330 13088
rect 5394 13024 5410 13088
rect 5474 13024 5490 13088
rect 5554 13024 5570 13088
rect 5634 13024 5643 13088
rect 5322 12000 5643 13024
rect 5322 11936 5330 12000
rect 5394 11936 5410 12000
rect 5474 11936 5490 12000
rect 5554 11936 5570 12000
rect 5634 11936 5643 12000
rect 5322 10912 5643 11936
rect 5322 10848 5330 10912
rect 5394 10848 5410 10912
rect 5474 10848 5490 10912
rect 5554 10848 5570 10912
rect 5634 10848 5643 10912
rect 5322 9824 5643 10848
rect 5322 9760 5330 9824
rect 5394 9760 5410 9824
rect 5474 9760 5490 9824
rect 5554 9760 5570 9824
rect 5634 9760 5643 9824
rect 5322 8736 5643 9760
rect 5322 8672 5330 8736
rect 5394 8672 5410 8736
rect 5474 8672 5490 8736
rect 5554 8672 5570 8736
rect 5634 8672 5643 8736
rect 5322 7648 5643 8672
rect 5322 7584 5330 7648
rect 5394 7584 5410 7648
rect 5474 7584 5490 7648
rect 5554 7584 5570 7648
rect 5634 7584 5643 7648
rect 5322 6560 5643 7584
rect 5322 6496 5330 6560
rect 5394 6496 5410 6560
rect 5474 6496 5490 6560
rect 5554 6496 5570 6560
rect 5634 6496 5643 6560
rect 5322 5472 5643 6496
rect 5322 5408 5330 5472
rect 5394 5408 5410 5472
rect 5474 5408 5490 5472
rect 5554 5408 5570 5472
rect 5634 5408 5643 5472
rect 5322 4384 5643 5408
rect 5322 4320 5330 4384
rect 5394 4320 5410 4384
rect 5474 4320 5490 4384
rect 5554 4320 5570 4384
rect 5634 4320 5643 4384
rect 5322 3296 5643 4320
rect 5322 3232 5330 3296
rect 5394 3232 5410 3296
rect 5474 3232 5490 3296
rect 5554 3232 5570 3296
rect 5634 3232 5643 3296
rect 5322 2208 5643 3232
rect 5322 2144 5330 2208
rect 5394 2144 5410 2208
rect 5474 2144 5490 2208
rect 5554 2144 5570 2208
rect 5634 2144 5643 2208
rect 5322 2128 5643 2144
rect 9989 25600 10309 25616
rect 9989 25536 9997 25600
rect 10061 25536 10077 25600
rect 10141 25536 10157 25600
rect 10221 25536 10237 25600
rect 10301 25536 10309 25600
rect 9989 24512 10309 25536
rect 9989 24448 9997 24512
rect 10061 24448 10077 24512
rect 10141 24448 10157 24512
rect 10221 24448 10237 24512
rect 10301 24448 10309 24512
rect 9989 23424 10309 24448
rect 9989 23360 9997 23424
rect 10061 23360 10077 23424
rect 10141 23360 10157 23424
rect 10221 23360 10237 23424
rect 10301 23360 10309 23424
rect 9989 22336 10309 23360
rect 9989 22272 9997 22336
rect 10061 22272 10077 22336
rect 10141 22272 10157 22336
rect 10221 22272 10237 22336
rect 10301 22272 10309 22336
rect 9989 21248 10309 22272
rect 9989 21184 9997 21248
rect 10061 21184 10077 21248
rect 10141 21184 10157 21248
rect 10221 21184 10237 21248
rect 10301 21184 10309 21248
rect 9989 20160 10309 21184
rect 9989 20096 9997 20160
rect 10061 20096 10077 20160
rect 10141 20096 10157 20160
rect 10221 20096 10237 20160
rect 10301 20096 10309 20160
rect 9989 19072 10309 20096
rect 9989 19008 9997 19072
rect 10061 19008 10077 19072
rect 10141 19008 10157 19072
rect 10221 19008 10237 19072
rect 10301 19008 10309 19072
rect 9989 17984 10309 19008
rect 9989 17920 9997 17984
rect 10061 17920 10077 17984
rect 10141 17920 10157 17984
rect 10221 17920 10237 17984
rect 10301 17920 10309 17984
rect 9989 16896 10309 17920
rect 9989 16832 9997 16896
rect 10061 16832 10077 16896
rect 10141 16832 10157 16896
rect 10221 16832 10237 16896
rect 10301 16832 10309 16896
rect 9989 15808 10309 16832
rect 9989 15744 9997 15808
rect 10061 15744 10077 15808
rect 10141 15744 10157 15808
rect 10221 15744 10237 15808
rect 10301 15744 10309 15808
rect 9989 14720 10309 15744
rect 9989 14656 9997 14720
rect 10061 14656 10077 14720
rect 10141 14656 10157 14720
rect 10221 14656 10237 14720
rect 10301 14656 10309 14720
rect 9989 13632 10309 14656
rect 9989 13568 9997 13632
rect 10061 13568 10077 13632
rect 10141 13568 10157 13632
rect 10221 13568 10237 13632
rect 10301 13568 10309 13632
rect 9989 12544 10309 13568
rect 9989 12480 9997 12544
rect 10061 12480 10077 12544
rect 10141 12480 10157 12544
rect 10221 12480 10237 12544
rect 10301 12480 10309 12544
rect 9989 11456 10309 12480
rect 9989 11392 9997 11456
rect 10061 11392 10077 11456
rect 10141 11392 10157 11456
rect 10221 11392 10237 11456
rect 10301 11392 10309 11456
rect 9989 10368 10309 11392
rect 9989 10304 9997 10368
rect 10061 10304 10077 10368
rect 10141 10304 10157 10368
rect 10221 10304 10237 10368
rect 10301 10304 10309 10368
rect 9989 9280 10309 10304
rect 9989 9216 9997 9280
rect 10061 9216 10077 9280
rect 10141 9216 10157 9280
rect 10221 9216 10237 9280
rect 10301 9216 10309 9280
rect 9989 8192 10309 9216
rect 9989 8128 9997 8192
rect 10061 8128 10077 8192
rect 10141 8128 10157 8192
rect 10221 8128 10237 8192
rect 10301 8128 10309 8192
rect 9989 7104 10309 8128
rect 9989 7040 9997 7104
rect 10061 7040 10077 7104
rect 10141 7040 10157 7104
rect 10221 7040 10237 7104
rect 10301 7040 10309 7104
rect 9989 6016 10309 7040
rect 9989 5952 9997 6016
rect 10061 5952 10077 6016
rect 10141 5952 10157 6016
rect 10221 5952 10237 6016
rect 10301 5952 10309 6016
rect 9989 4928 10309 5952
rect 9989 4864 9997 4928
rect 10061 4864 10077 4928
rect 10141 4864 10157 4928
rect 10221 4864 10237 4928
rect 10301 4864 10309 4928
rect 9989 3840 10309 4864
rect 14656 25056 14976 25616
rect 14656 24992 14664 25056
rect 14728 24992 14744 25056
rect 14808 24992 14824 25056
rect 14888 24992 14904 25056
rect 14968 24992 14976 25056
rect 14656 23968 14976 24992
rect 14656 23904 14664 23968
rect 14728 23904 14744 23968
rect 14808 23904 14824 23968
rect 14888 23904 14904 23968
rect 14968 23904 14976 23968
rect 14656 22880 14976 23904
rect 14656 22816 14664 22880
rect 14728 22816 14744 22880
rect 14808 22816 14824 22880
rect 14888 22816 14904 22880
rect 14968 22816 14976 22880
rect 14656 21792 14976 22816
rect 14656 21728 14664 21792
rect 14728 21728 14744 21792
rect 14808 21728 14824 21792
rect 14888 21728 14904 21792
rect 14968 21728 14976 21792
rect 14656 20704 14976 21728
rect 14656 20640 14664 20704
rect 14728 20640 14744 20704
rect 14808 20640 14824 20704
rect 14888 20640 14904 20704
rect 14968 20640 14976 20704
rect 14656 19616 14976 20640
rect 14656 19552 14664 19616
rect 14728 19552 14744 19616
rect 14808 19552 14824 19616
rect 14888 19552 14904 19616
rect 14968 19552 14976 19616
rect 14656 18528 14976 19552
rect 14656 18464 14664 18528
rect 14728 18464 14744 18528
rect 14808 18464 14824 18528
rect 14888 18464 14904 18528
rect 14968 18464 14976 18528
rect 14656 17440 14976 18464
rect 14656 17376 14664 17440
rect 14728 17376 14744 17440
rect 14808 17376 14824 17440
rect 14888 17376 14904 17440
rect 14968 17376 14976 17440
rect 14656 16352 14976 17376
rect 14656 16288 14664 16352
rect 14728 16288 14744 16352
rect 14808 16288 14824 16352
rect 14888 16288 14904 16352
rect 14968 16288 14976 16352
rect 14656 15264 14976 16288
rect 14656 15200 14664 15264
rect 14728 15200 14744 15264
rect 14808 15200 14824 15264
rect 14888 15200 14904 15264
rect 14968 15200 14976 15264
rect 14656 14176 14976 15200
rect 14656 14112 14664 14176
rect 14728 14112 14744 14176
rect 14808 14112 14824 14176
rect 14888 14112 14904 14176
rect 14968 14112 14976 14176
rect 14656 13088 14976 14112
rect 14656 13024 14664 13088
rect 14728 13024 14744 13088
rect 14808 13024 14824 13088
rect 14888 13024 14904 13088
rect 14968 13024 14976 13088
rect 14656 12000 14976 13024
rect 14656 11936 14664 12000
rect 14728 11936 14744 12000
rect 14808 11936 14824 12000
rect 14888 11936 14904 12000
rect 14968 11936 14976 12000
rect 14656 10912 14976 11936
rect 14656 10848 14664 10912
rect 14728 10848 14744 10912
rect 14808 10848 14824 10912
rect 14888 10848 14904 10912
rect 14968 10848 14976 10912
rect 14656 9824 14976 10848
rect 14656 9760 14664 9824
rect 14728 9760 14744 9824
rect 14808 9760 14824 9824
rect 14888 9760 14904 9824
rect 14968 9760 14976 9824
rect 14656 8736 14976 9760
rect 14656 8672 14664 8736
rect 14728 8672 14744 8736
rect 14808 8672 14824 8736
rect 14888 8672 14904 8736
rect 14968 8672 14976 8736
rect 14656 7648 14976 8672
rect 14656 7584 14664 7648
rect 14728 7584 14744 7648
rect 14808 7584 14824 7648
rect 14888 7584 14904 7648
rect 14968 7584 14976 7648
rect 14656 6560 14976 7584
rect 14656 6496 14664 6560
rect 14728 6496 14744 6560
rect 14808 6496 14824 6560
rect 14888 6496 14904 6560
rect 14968 6496 14976 6560
rect 14656 5472 14976 6496
rect 14656 5408 14664 5472
rect 14728 5408 14744 5472
rect 14808 5408 14824 5472
rect 14888 5408 14904 5472
rect 14968 5408 14976 5472
rect 14656 4384 14976 5408
rect 14656 4320 14664 4384
rect 14728 4320 14744 4384
rect 14808 4320 14824 4384
rect 14888 4320 14904 4384
rect 14968 4320 14976 4384
rect 9989 3776 9997 3840
rect 10061 3776 10077 3840
rect 10141 3776 10157 3840
rect 10221 3776 10237 3840
rect 10301 3776 10309 3840
rect 9989 2752 10309 3776
rect 9989 2688 9997 2752
rect 10061 2688 10077 2752
rect 10141 2688 10157 2752
rect 10221 2688 10237 2752
rect 10301 2688 10309 2752
rect 9989 2128 10309 2688
rect 14656 3296 14976 4320
rect 14656 3232 14664 3296
rect 14728 3232 14744 3296
rect 14808 3232 14824 3296
rect 14888 3232 14904 3296
rect 14968 3232 14976 3296
rect 14656 2208 14976 3232
rect 14656 2144 14664 2208
rect 14728 2144 14744 2208
rect 14808 2144 14824 2208
rect 14888 2144 14904 2208
rect 14968 2144 14976 2208
rect 14656 2128 14976 2144
rect 19322 25600 19642 25616
rect 19322 25536 19330 25600
rect 19394 25536 19410 25600
rect 19474 25536 19490 25600
rect 19554 25536 19570 25600
rect 19634 25536 19642 25600
rect 19322 24512 19642 25536
rect 19322 24448 19330 24512
rect 19394 24448 19410 24512
rect 19474 24448 19490 24512
rect 19554 24448 19570 24512
rect 19634 24448 19642 24512
rect 19322 23424 19642 24448
rect 19322 23360 19330 23424
rect 19394 23360 19410 23424
rect 19474 23360 19490 23424
rect 19554 23360 19570 23424
rect 19634 23360 19642 23424
rect 19322 22336 19642 23360
rect 19322 22272 19330 22336
rect 19394 22272 19410 22336
rect 19474 22272 19490 22336
rect 19554 22272 19570 22336
rect 19634 22272 19642 22336
rect 19322 21248 19642 22272
rect 19322 21184 19330 21248
rect 19394 21184 19410 21248
rect 19474 21184 19490 21248
rect 19554 21184 19570 21248
rect 19634 21184 19642 21248
rect 19322 20160 19642 21184
rect 19322 20096 19330 20160
rect 19394 20096 19410 20160
rect 19474 20096 19490 20160
rect 19554 20096 19570 20160
rect 19634 20096 19642 20160
rect 19322 19072 19642 20096
rect 23694 19413 23754 27643
rect 23989 25056 24309 25616
rect 23989 24992 23997 25056
rect 24061 24992 24077 25056
rect 24141 24992 24157 25056
rect 24221 24992 24237 25056
rect 24301 24992 24309 25056
rect 23989 23968 24309 24992
rect 23989 23904 23997 23968
rect 24061 23904 24077 23968
rect 24141 23904 24157 23968
rect 24221 23904 24237 23968
rect 24301 23904 24309 23968
rect 23989 22880 24309 23904
rect 23989 22816 23997 22880
rect 24061 22816 24077 22880
rect 24141 22816 24157 22880
rect 24221 22816 24237 22880
rect 24301 22816 24309 22880
rect 23989 21792 24309 22816
rect 23989 21728 23997 21792
rect 24061 21728 24077 21792
rect 24141 21728 24157 21792
rect 24221 21728 24237 21792
rect 24301 21728 24309 21792
rect 23989 20704 24309 21728
rect 23989 20640 23997 20704
rect 24061 20640 24077 20704
rect 24141 20640 24157 20704
rect 24221 20640 24237 20704
rect 24301 20640 24309 20704
rect 23989 19616 24309 20640
rect 23989 19552 23997 19616
rect 24061 19552 24077 19616
rect 24141 19552 24157 19616
rect 24221 19552 24237 19616
rect 24301 19552 24309 19616
rect 23691 19412 23757 19413
rect 23691 19348 23692 19412
rect 23756 19348 23757 19412
rect 23691 19347 23757 19348
rect 19322 19008 19330 19072
rect 19394 19008 19410 19072
rect 19474 19008 19490 19072
rect 19554 19008 19570 19072
rect 19634 19008 19642 19072
rect 19322 17984 19642 19008
rect 19322 17920 19330 17984
rect 19394 17920 19410 17984
rect 19474 17920 19490 17984
rect 19554 17920 19570 17984
rect 19634 17920 19642 17984
rect 19322 16896 19642 17920
rect 19322 16832 19330 16896
rect 19394 16832 19410 16896
rect 19474 16832 19490 16896
rect 19554 16832 19570 16896
rect 19634 16832 19642 16896
rect 19322 15808 19642 16832
rect 19322 15744 19330 15808
rect 19394 15744 19410 15808
rect 19474 15744 19490 15808
rect 19554 15744 19570 15808
rect 19634 15744 19642 15808
rect 19322 14720 19642 15744
rect 19322 14656 19330 14720
rect 19394 14656 19410 14720
rect 19474 14656 19490 14720
rect 19554 14656 19570 14720
rect 19634 14656 19642 14720
rect 19322 13632 19642 14656
rect 19322 13568 19330 13632
rect 19394 13568 19410 13632
rect 19474 13568 19490 13632
rect 19554 13568 19570 13632
rect 19634 13568 19642 13632
rect 19322 12544 19642 13568
rect 19322 12480 19330 12544
rect 19394 12480 19410 12544
rect 19474 12480 19490 12544
rect 19554 12480 19570 12544
rect 19634 12480 19642 12544
rect 19322 11456 19642 12480
rect 19322 11392 19330 11456
rect 19394 11392 19410 11456
rect 19474 11392 19490 11456
rect 19554 11392 19570 11456
rect 19634 11392 19642 11456
rect 19322 10368 19642 11392
rect 19322 10304 19330 10368
rect 19394 10304 19410 10368
rect 19474 10304 19490 10368
rect 19554 10304 19570 10368
rect 19634 10304 19642 10368
rect 19322 9280 19642 10304
rect 19322 9216 19330 9280
rect 19394 9216 19410 9280
rect 19474 9216 19490 9280
rect 19554 9216 19570 9280
rect 19634 9216 19642 9280
rect 19322 8192 19642 9216
rect 19322 8128 19330 8192
rect 19394 8128 19410 8192
rect 19474 8128 19490 8192
rect 19554 8128 19570 8192
rect 19634 8128 19642 8192
rect 19322 7104 19642 8128
rect 19322 7040 19330 7104
rect 19394 7040 19410 7104
rect 19474 7040 19490 7104
rect 19554 7040 19570 7104
rect 19634 7040 19642 7104
rect 19322 6016 19642 7040
rect 19322 5952 19330 6016
rect 19394 5952 19410 6016
rect 19474 5952 19490 6016
rect 19554 5952 19570 6016
rect 19634 5952 19642 6016
rect 19322 4928 19642 5952
rect 19322 4864 19330 4928
rect 19394 4864 19410 4928
rect 19474 4864 19490 4928
rect 19554 4864 19570 4928
rect 19634 4864 19642 4928
rect 19322 3840 19642 4864
rect 19322 3776 19330 3840
rect 19394 3776 19410 3840
rect 19474 3776 19490 3840
rect 19554 3776 19570 3840
rect 19634 3776 19642 3840
rect 19322 2752 19642 3776
rect 19322 2688 19330 2752
rect 19394 2688 19410 2752
rect 19474 2688 19490 2752
rect 19554 2688 19570 2752
rect 19634 2688 19642 2752
rect 19322 2128 19642 2688
rect 23989 18528 24309 19552
rect 23989 18464 23997 18528
rect 24061 18464 24077 18528
rect 24141 18464 24157 18528
rect 24221 18464 24237 18528
rect 24301 18464 24309 18528
rect 23989 17440 24309 18464
rect 23989 17376 23997 17440
rect 24061 17376 24077 17440
rect 24141 17376 24157 17440
rect 24221 17376 24237 17440
rect 24301 17376 24309 17440
rect 23989 16352 24309 17376
rect 23989 16288 23997 16352
rect 24061 16288 24077 16352
rect 24141 16288 24157 16352
rect 24221 16288 24237 16352
rect 24301 16288 24309 16352
rect 23989 15264 24309 16288
rect 23989 15200 23997 15264
rect 24061 15200 24077 15264
rect 24141 15200 24157 15264
rect 24221 15200 24237 15264
rect 24301 15200 24309 15264
rect 23989 14176 24309 15200
rect 23989 14112 23997 14176
rect 24061 14112 24077 14176
rect 24141 14112 24157 14176
rect 24221 14112 24237 14176
rect 24301 14112 24309 14176
rect 23989 13088 24309 14112
rect 23989 13024 23997 13088
rect 24061 13024 24077 13088
rect 24141 13024 24157 13088
rect 24221 13024 24237 13088
rect 24301 13024 24309 13088
rect 23989 12000 24309 13024
rect 23989 11936 23997 12000
rect 24061 11936 24077 12000
rect 24141 11936 24157 12000
rect 24221 11936 24237 12000
rect 24301 11936 24309 12000
rect 23989 10912 24309 11936
rect 23989 10848 23997 10912
rect 24061 10848 24077 10912
rect 24141 10848 24157 10912
rect 24221 10848 24237 10912
rect 24301 10848 24309 10912
rect 23989 9824 24309 10848
rect 23989 9760 23997 9824
rect 24061 9760 24077 9824
rect 24141 9760 24157 9824
rect 24221 9760 24237 9824
rect 24301 9760 24309 9824
rect 23989 8736 24309 9760
rect 23989 8672 23997 8736
rect 24061 8672 24077 8736
rect 24141 8672 24157 8736
rect 24221 8672 24237 8736
rect 24301 8672 24309 8736
rect 23989 7648 24309 8672
rect 23989 7584 23997 7648
rect 24061 7584 24077 7648
rect 24141 7584 24157 7648
rect 24221 7584 24237 7648
rect 24301 7584 24309 7648
rect 23989 6560 24309 7584
rect 23989 6496 23997 6560
rect 24061 6496 24077 6560
rect 24141 6496 24157 6560
rect 24221 6496 24237 6560
rect 24301 6496 24309 6560
rect 23989 5472 24309 6496
rect 23989 5408 23997 5472
rect 24061 5408 24077 5472
rect 24141 5408 24157 5472
rect 24221 5408 24237 5472
rect 24301 5408 24309 5472
rect 23989 4384 24309 5408
rect 23989 4320 23997 4384
rect 24061 4320 24077 4384
rect 24141 4320 24157 4384
rect 24221 4320 24237 4384
rect 24301 4320 24309 4384
rect 23989 3296 24309 4320
rect 23989 3232 23997 3296
rect 24061 3232 24077 3296
rect 24141 3232 24157 3296
rect 24221 3232 24237 3296
rect 24301 3232 24309 3296
rect 23989 2208 24309 3232
rect 24614 2957 24674 3622
rect 24611 2956 24677 2957
rect 24611 2892 24612 2956
rect 24676 2892 24677 2956
rect 24611 2891 24677 2892
rect 23989 2144 23997 2208
rect 24061 2144 24077 2208
rect 24141 2144 24157 2208
rect 24221 2144 24237 2208
rect 24301 2144 24309 2208
rect 23989 2128 24309 2144
<< via4 >>
rect 11462 3772 11698 3858
rect 11462 3708 11548 3772
rect 11548 3708 11612 3772
rect 11612 3708 11698 3772
rect 11462 3622 11698 3708
rect 24526 3622 24762 3858
<< metal5 >>
rect 11420 3858 24804 3900
rect 11420 3622 11462 3858
rect 11698 3622 24526 3858
rect 24762 3622 24804 3858
rect 11420 3580 24804 3622
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 816 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 816 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1092 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2196 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1092 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2196 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3668 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 3760 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3300 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4404 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6520 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6428 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 4864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5508 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_62
timestamp 1604681595
transform 1 0 6520 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1604681595
transform 1 0 7440 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp 1604681595
transform 1 0 7072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604681595
transform 1 0 6612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7164 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1604681595
transform 1 0 7808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7624 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 7992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7808 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _72_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8176 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_88
timestamp 1604681595
transform 1 0 8912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_84
timestamp 1604681595
transform 1 0 8544 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__90__A
timestamp 1604681595
transform 1 0 8820 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 8728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9372 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1604681595
transform 1 0 9924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1604681595
transform 1 0 9464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 9556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9280 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_111
timestamp 1604681595
transform 1 0 11028 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10660 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_115
timestamp 1604681595
transform 1 0 11396 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12040 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 11856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12224 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1604681595
transform 1 0 12132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12316 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13972 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12408 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13788 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1604681595
transform 1 0 14064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_135
timestamp 1604681595
transform 1 0 13236 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1604681595
transform 1 0 13604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15168 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15076 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148
timestamp 1604681595
transform 1 0 14432 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_162
timestamp 1604681595
transform 1 0 15720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1604681595
transform 1 0 16088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_174
timestamp 1604681595
transform 1 0 16824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1604681595
transform 1 0 16916 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 16456 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1604681595
transform 1 0 17560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1604681595
transform 1 0 17192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1604681595
transform 1 0 17652 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1604681595
transform 1 0 17284 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17652 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17744 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18020 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19676 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1604681595
transform 1 0 19768 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1604681595
transform 1 0 19492 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_207
timestamp 1604681595
transform 1 0 19860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20872 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20228 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 20780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp 1604681595
transform 1 0 20136 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1604681595
transform 1 0 22344 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_230
timestamp 1604681595
transform 1 0 21976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1604681595
transform 1 0 22620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 22712 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 22896 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1604681595
transform 1 0 23540 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_243
timestamp 1604681595
transform 1 0 23172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23080 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23264 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23632 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23356 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23724 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_254
timestamp 1604681595
transform 1 0 24184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1604681595
transform 1 0 24552 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604681595
transform 1 0 24920 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24736 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25104 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 24920 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_266
timestamp 1604681595
transform 1 0 25288 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_269
timestamp 1604681595
transform 1 0 25564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 25288 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_270
timestamp 1604681595
transform 1 0 25656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26576 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604681595
transform 1 0 25932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_274
timestamp 1604681595
transform 1 0 26024 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3668 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 3760 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 4864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 5968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 8176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1604681595
transform 1 0 7072 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1604681595
transform 1 0 7440 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1604681595
transform 1 0 7716 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_79
timestamp 1604681595
transform 1 0 8084 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9372 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9280 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9096 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 8912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11856 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11304 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1604681595
transform 1 0 11120 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1604681595
transform 1 0 11488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_139
timestamp 1604681595
transform 1 0 13604 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1604681595
transform 1 0 14064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14984 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 14892 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1604681595
transform 1 0 15996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_148
timestamp 1604681595
transform 1 0 14432 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1604681595
transform 1 0 15812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16548 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17560 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16364 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1604681595
transform 1 0 16180 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1604681595
transform 1 0 17376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_184
timestamp 1604681595
transform 1 0 17744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18112 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19124 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1604681595
transform 1 0 18940 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_201
timestamp 1604681595
transform 1 0 19308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604681595
transform 1 0 19768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20780 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21792 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20320 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20136 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1604681595
transform 1 0 20596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_226
timestamp 1604681595
transform 1 0 21608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23264 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22528 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_230
timestamp 1604681595
transform 1 0 21976 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_234
timestamp 1604681595
transform 1 0 22344 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_238
timestamp 1604681595
transform 1 0 22712 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25012 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26576 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26116 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26208 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1092 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2196 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3300 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4404 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 6520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6428 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5508 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6244 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7532 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_65
timestamp 1604681595
transform 1 0 6796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_69
timestamp 1604681595
transform 1 0 7164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1604681595
transform 1 0 8360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9096 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1604681595
transform 1 0 8728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1604681595
transform 1 0 9924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1604681595
transform 1 0 10292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 10936 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12132 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12040 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 11488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_107
timestamp 1604681595
transform 1 0 10660 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13880 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13328 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1604681595
transform 1 0 12960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1604681595
transform 1 0 13512 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_161
timestamp 1604681595
transform 1 0 15628 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1604681595
transform 1 0 15996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 16364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17744 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17652 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1604681595
transform 1 0 16180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_173
timestamp 1604681595
transform 1 0 16732 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19584 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1604681595
transform 1 0 18940 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_201
timestamp 1604681595
transform 1 0 19308 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21148 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20964 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20596 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1604681595
transform 1 0 20412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1604681595
transform 1 0 20780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23264 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22160 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22528 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_230
timestamp 1604681595
transform 1 0 21976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_234
timestamp 1604681595
transform 1 0 22344 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1604681595
transform 1 0 22712 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1604681595
transform 1 0 23356 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23908 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 24920 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_260
timestamp 1604681595
transform 1 0 24736 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1604681595
transform 1 0 25104 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26576 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26208 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 816 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3668 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3300 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 3760 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 4864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 5968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 8268 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_68
timestamp 1604681595
transform 1 0 7072 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_74
timestamp 1604681595
transform 1 0 7624 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1604681595
transform 1 0 7900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1604681595
transform 1 0 9372 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 8912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9280 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1604681595
transform 1 0 10016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp 1604681595
transform 1 0 9740 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10108 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_120
timestamp 1604681595
transform 1 0 11856 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1604681595
transform 1 0 12316 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13328 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12684 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_132
timestamp 1604681595
transform 1 0 12960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15628 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 14892 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1604681595
transform 1 0 14984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_158
timestamp 1604681595
transform 1 0 15352 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17192 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_170
timestamp 1604681595
transform 1 0 16456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1604681595
transform 1 0 16824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_187
timestamp 1604681595
transform 1 0 18020 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18572 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_191
timestamp 1604681595
transform 1 0 18388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1604681595
transform 1 0 19584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_208
timestamp 1604681595
transform 1 0 19952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 20596 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21608 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20136 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1604681595
transform 1 0 20320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_218
timestamp 1604681595
transform 1 0 20872 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_223
timestamp 1604681595
transform 1 0 21332 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23172 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22988 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22620 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_235
timestamp 1604681595
transform 1 0 22436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_239
timestamp 1604681595
transform 1 0 22804 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 24736 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24184 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24552 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_252
timestamp 1604681595
transform 1 0 24000 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_256
timestamp 1604681595
transform 1 0 24368 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_264
timestamp 1604681595
transform 1 0 25104 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26576 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_272
timestamp 1604681595
transform 1 0 25840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26208 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 816 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1092 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2196 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3300 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4404 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6428 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5508 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1604681595
transform 1 0 6520 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 7532 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7992 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_70
timestamp 1604681595
transform 1 0 7256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_76
timestamp 1604681595
transform 1 0 7808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_80
timestamp 1604681595
transform 1 0 8176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8544 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1604681595
transform 1 0 9372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1604681595
transform 1 0 9740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1604681595
transform 1 0 10108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12132 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10476 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12040 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11856 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14064 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1604681595
transform 1 0 13880 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15168 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 14616 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1604681595
transform 1 0 14248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_153
timestamp 1604681595
transform 1 0 14892 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17744 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17652 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 16916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 19676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 19308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19124 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1604681595
transform 1 0 18572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1604681595
transform 1 0 18940 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1604681595
transform 1 0 19584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20780 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20596 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_209
timestamp 1604681595
transform 1 0 20044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_213
timestamp 1604681595
transform 1 0 20412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23540 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23264 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23080 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 22712 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22528 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 22896 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_245
timestamp 1604681595
transform 1 0 23356 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 25104 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 25656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24552 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24920 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_256
timestamp 1604681595
transform 1 0 24368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_260
timestamp 1604681595
transform 1 0 24736 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_268
timestamp 1604681595
transform 1 0 25472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26576 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_272
timestamp 1604681595
transform 1 0 25840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26208 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 816 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 816 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1092 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2196 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3668 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3300 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 3760 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3300 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4404 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 4864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 5968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5508 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1604681595
transform 1 0 6520 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_67
timestamp 1604681595
transform 1 0 6980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_68
timestamp 1604681595
transform 1 0 7072 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1604681595
transform 1 0 7716 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 1604681595
transform 1 0 7624 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7900 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7716 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8084 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604681595
transform 1 0 9372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1604681595
transform 1 0 8912 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8544 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9096 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9280 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1604681595
transform 1 0 10200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1604681595
transform 1 0 9832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1604681595
transform 1 0 9740 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9832 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_106
timestamp 1604681595
transform 1 0 10568 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1604681595
transform 1 0 11028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_107
timestamp 1604681595
transform 1 0 10660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 11028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1604681595
transform 1 0 12132 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12040 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12224 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11396 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 1604681595
transform 1 0 13052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_134
timestamp 1604681595
transform 1 0 13144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13236 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_137
timestamp 1604681595
transform 1 0 13420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604681595
transform 1 0 14156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1604681595
transform 1 0 13512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 13880 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13788 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604681595
transform 1 0 14524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 14892 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 14984 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_164
timestamp 1604681595
transform 1 0 15904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1604681595
transform 1 0 15536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_162
timestamp 1604681595
transform 1 0 15720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_157
timestamp 1604681595
transform 1 0 15260 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 15720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15996 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 16916 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_168
timestamp 1604681595
transform 1 0 16272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1604681595
transform 1 0 16824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17008 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 17100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 16548 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1604681595
transform 1 0 17744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17284 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1604681595
transform 1 0 17192 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17376 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17468 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17652 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 17836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 17560 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18940 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 18388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19492 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 19860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1604681595
transform 1 0 19308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_205
timestamp 1604681595
transform 1 0 19676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_189
timestamp 1604681595
transform 1 0 18204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_216
timestamp 1604681595
transform 1 0 20688 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 1604681595
transform 1 0 20044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20320 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_224
timestamp 1604681595
transform 1 0 21424 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1604681595
transform 1 0 21056 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21700 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20596 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604681595
transform 1 0 22528 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_238
timestamp 1604681595
transform 1 0 22712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_234
timestamp 1604681595
transform 1 0 22344 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 22528 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 22712 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_245
timestamp 1604681595
transform 1 0 23356 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 22896 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_242
timestamp 1604681595
transform 1 0 23080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23080 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23264 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23448 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23448 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 25380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1604681595
transform 1 0 25196 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_265
timestamp 1604681595
transform 1 0 25196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_269
timestamp 1604681595
transform 1 0 25564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26576 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26576 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26116 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1604681595
transform 1 0 25932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26208 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_273
timestamp 1604681595
transform 1 0 25932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 816 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3668 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 3760 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 4864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_56
timestamp 1604681595
transform 1 0 5968 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6796 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1604681595
transform 1 0 6704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9372 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1604681595
transform 1 0 8544 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_102
timestamp 1604681595
transform 1 0 10200 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11396 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 11120 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10476 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_107
timestamp 1604681595
transform 1 0 10660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 13880 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1604681595
transform 1 0 13144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1604681595
transform 1 0 13512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 15168 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15536 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 14892 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604681595
transform 1 0 14984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16364 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18848 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19860 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1604681595
transform 1 0 18112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_192
timestamp 1604681595
transform 1 0 18480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1604681595
transform 1 0 19676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20596 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21700 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1604681595
transform 1 0 20044 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_224
timestamp 1604681595
transform 1 0 21424 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_229
timestamp 1604681595
transform 1 0 21884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 22252 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22068 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 24736 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24184 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24552 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_252
timestamp 1604681595
transform 1 0 24000 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_256
timestamp 1604681595
transform 1 0 24368 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_264
timestamp 1604681595
transform 1 0 25104 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26576 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1604681595
transform 1 0 25840 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26208 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 816 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1092 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2196 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3300 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4404 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5508 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6520 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7808 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7624 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1604681595
transform 1 0 9556 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1604681595
transform 1 0 10108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10476 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12040 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1604681595
transform 1 0 12132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12684 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12500 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 15168 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 14984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_148
timestamp 1604681595
transform 1 0 14432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1604681595
transform 1 0 14800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17744 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17652 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17468 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_176
timestamp 1604681595
transform 1 0 17008 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_180
timestamp 1604681595
transform 1 0 17376 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19308 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19124 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1604681595
transform 1 0 18572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1604681595
transform 1 0 18940 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20320 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20688 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_210
timestamp 1604681595
transform 1 0 20136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_214
timestamp 1604681595
transform 1 0 20504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_227
timestamp 1604681595
transform 1 0 21700 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23448 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23264 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23080 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22712 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_231
timestamp 1604681595
transform 1 0 22068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604681595
transform 1 0 22528 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 22896 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_245
timestamp 1604681595
transform 1 0 23356 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 25012 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1604681595
transform 1 0 24736 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 25564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1604681595
transform 1 0 24276 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_259
timestamp 1604681595
transform 1 0 24644 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_262
timestamp 1604681595
transform 1 0 24920 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_267
timestamp 1604681595
transform 1 0 25380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26576 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_271
timestamp 1604681595
transform 1 0 25748 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 816 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 3760 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 4864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 5968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_68
timestamp 1604681595
transform 1 0 7072 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_78
timestamp 1604681595
transform 1 0 7992 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 9372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9280 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1604681595
transform 1 0 9096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp 1604681595
transform 1 0 9648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1604681595
transform 1 0 10384 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10660 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10476 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13144 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_126
timestamp 1604681595
transform 1 0 12408 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_131
timestamp 1604681595
transform 1 0 12868 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_143
timestamp 1604681595
transform 1 0 13972 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14984 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 14892 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1604681595
transform 1 0 14524 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17468 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1604681595
transform 1 0 16732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1604681595
transform 1 0 17100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 19216 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19952 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_190
timestamp 1604681595
transform 1 0 18296 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1604681595
transform 1 0 18664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_198
timestamp 1604681595
transform 1 0 19032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1604681595
transform 1 0 19768 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20596 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20320 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_210
timestamp 1604681595
transform 1 0 20136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23172 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22528 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_234
timestamp 1604681595
transform 1 0 22344 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_238
timestamp 1604681595
transform 1 0 22712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_242
timestamp 1604681595
transform 1 0 23080 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 24736 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24184 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24552 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_252
timestamp 1604681595
transform 1 0 24000 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_256
timestamp 1604681595
transform 1 0 24368 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_264
timestamp 1604681595
transform 1 0 25104 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26576 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_272
timestamp 1604681595
transform 1 0 25840 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26208 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 816 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1092 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2196 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3300 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4404 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6428 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5508 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6520 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7624 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9464 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1604681595
transform 1 0 8728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_90
timestamp 1604681595
transform 1 0 9096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 12132 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12040 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1604681595
transform 1 0 11212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp 1604681595
transform 1 0 11580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 11948 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13512 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13328 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_126
timestamp 1604681595
transform 1 0 12408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_130
timestamp 1604681595
transform 1 0 12776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1604681595
transform 1 0 13144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15168 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_147
timestamp 1604681595
transform 1 0 14340 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1604681595
transform 1 0 14800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17652 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17284 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 17928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_175
timestamp 1604681595
transform 1 0 16916 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1604681595
transform 1 0 17468 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1604681595
transform 1 0 17744 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18572 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_188
timestamp 1604681595
transform 1 0 18112 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21700 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21516 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20596 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_212
timestamp 1604681595
transform 1 0 20320 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1604681595
transform 1 0 20780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_221
timestamp 1604681595
transform 1 0 21148 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23356 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23264 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23080 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604681595
transform 1 0 22528 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 22896 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_264
timestamp 1604681595
transform 1 0 25104 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26208 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 816 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3668 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3300 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 3760 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 4864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 5968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9280 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604681595
transform 1 0 9372 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_101
timestamp 1604681595
transform 1 0 10108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12132 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10568 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_115
timestamp 1604681595
transform 1 0 11396 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_142
timestamp 1604681595
transform 1 0 13880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14984 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 14892 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16088 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_146
timestamp 1604681595
transform 1 0 14248 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_150
timestamp 1604681595
transform 1 0 14616 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_163
timestamp 1604681595
transform 1 0 15812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17284 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 17008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16456 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16824 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_168
timestamp 1604681595
transform 1 0 16272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_172
timestamp 1604681595
transform 1 0 16640 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19216 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_198
timestamp 1604681595
transform 1 0 19032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_202
timestamp 1604681595
transform 1 0 19400 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_207
timestamp 1604681595
transform 1 0 19860 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20596 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21700 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20320 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_211
timestamp 1604681595
transform 1 0 20228 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_224
timestamp 1604681595
transform 1 0 21424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_229
timestamp 1604681595
transform 1 0 21884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23080 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22528 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_233
timestamp 1604681595
transform 1 0 22252 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_238
timestamp 1604681595
transform 1 0 22712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_261
timestamp 1604681595
transform 1 0 24828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1604681595
transform 1 0 25196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26576 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26116 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1604681595
transform 1 0 25932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26208 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 816 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 816 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1092 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2196 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3668 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4404 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3300 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 3760 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6428 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5508 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6520 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 4864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 5968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7624 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9280 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 8728 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 9832 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9372 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 11028 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12040 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_110
timestamp 1604681595
transform 1 0 10936 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11304 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1604681595
transform 1 0 12132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10476 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604681595
transform 1 0 11580 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1604681595
transform 1 0 12684 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_131
timestamp 1604681595
transform 1 0 12868 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_127
timestamp 1604681595
transform 1 0 12500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 12592 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604681595
transform 1 0 14156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1604681595
transform 1 0 13788 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_137
timestamp 1604681595
transform 1 0 13420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 13880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13604 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1604681595
transform 1 0 14984 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604681595
transform 1 0 14524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 14892 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1604681595
transform 1 0 15720 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1604681595
transform 1 0 15352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16088 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15076 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1604681595
transform 1 0 16824 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604681595
transform 1 0 16916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604681595
transform 1 0 17284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_178
timestamp 1604681595
transform 1 0 17192 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1604681595
transform 1 0 17468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 17836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17652 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 17652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17744 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_192
timestamp 1604681595
transform 1 0 18480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1604681595
transform 1 0 18112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_193
timestamp 1604681595
transform 1 0 18572 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18296 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18848 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18848 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_205
timestamp 1604681595
transform 1 0 19676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_204
timestamp 1604681595
transform 1 0 19584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_198
timestamp 1604681595
transform 1 0 19032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 19308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19676 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_215
timestamp 1604681595
transform 1 0 20596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_209
timestamp 1604681595
transform 1 0 20044 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20780 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_226
timestamp 1604681595
transform 1 0 21608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1604681595
transform 1 0 21792 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_224
timestamp 1604681595
transform 1 0 21424 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21792 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_235
timestamp 1604681595
transform 1 0 22436 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_230
timestamp 1604681595
transform 1 0 21976 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22528 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 22712 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 22160 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_240
timestamp 1604681595
transform 1 0 22896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 22896 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23080 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23264 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23356 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23264 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24920 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24736 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_254
timestamp 1604681595
transform 1 0 24184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_258
timestamp 1604681595
transform 1 0 24552 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_268
timestamp 1604681595
transform 1 0 25472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25012 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26576 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26576 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_272
timestamp 1604681595
transform 1 0 25840 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_276
timestamp 1604681595
transform 1 0 26208 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26208 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1092 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2196 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4404 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6428 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5508 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7624 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 8728 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 9832 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12040 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 10936 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12132 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14156 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13604 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13236 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_137
timestamp 1604681595
transform 1 0 13420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1604681595
transform 1 0 13788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16088 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15904 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1604681595
transform 1 0 14984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1604681595
transform 1 0 15352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604681595
transform 1 0 15720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 17744 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17652 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 16916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_187
timestamp 1604681595
transform 1 0 18020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18756 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1604681595
transform 1 0 18388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21700 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20688 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21056 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_214
timestamp 1604681595
transform 1 0 20504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1604681595
transform 1 0 20872 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_222
timestamp 1604681595
transform 1 0 21240 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23356 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23264 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23080 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22712 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604681595
transform 1 0 22528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 22896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1604681595
transform 1 0 25288 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1604681595
transform 1 0 25104 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_268
timestamp 1604681595
transform 1 0 25472 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26208 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 816 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3668 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 3760 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 4864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 5968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9280 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9372 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10476 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604681595
transform 1 0 11580 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13604 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_129
timestamp 1604681595
transform 1 0 12684 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1604681595
transform 1 0 13420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604681595
transform 1 0 14156 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14984 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 14892 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16088 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_160
timestamp 1604681595
transform 1 0 15536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_164
timestamp 1604681595
transform 1 0 15904 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16456 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1604681595
transform 1 0 16272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18940 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18756 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1604681595
transform 1 0 18204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1604681595
transform 1 0 18572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 19768 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20596 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21700 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604681595
transform 1 0 20136 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_224
timestamp 1604681595
transform 1 0 21424 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1604681595
transform 1 0 21884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22252 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 24736 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24184 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_252
timestamp 1604681595
transform 1 0 24000 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_256
timestamp 1604681595
transform 1 0 24368 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_264
timestamp 1604681595
transform 1 0 25104 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26576 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26116 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_272
timestamp 1604681595
transform 1 0 25840 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26208 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 816 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1092 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2196 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3300 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4404 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6428 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5508 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 8728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604681595
transform 1 0 9832 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12040 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 10936 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12132 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604681595
transform 1 0 13236 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15076 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_147
timestamp 1604681595
transform 1 0 14340 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1604681595
transform 1 0 15628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_165
timestamp 1604681595
transform 1 0 15996 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 16640 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17744 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17652 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_171
timestamp 1604681595
transform 1 0 16548 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 16916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19584 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1604681595
transform 1 0 18572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1604681595
transform 1 0 18940 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_201
timestamp 1604681595
transform 1 0 19308 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_223
timestamp 1604681595
transform 1 0 21332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_227
timestamp 1604681595
transform 1 0 21700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 22160 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23356 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23264 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1604681595
transform 1 0 22712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_231
timestamp 1604681595
transform 1 0 22068 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22528 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 22896 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 24920 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24736 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 25472 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_254
timestamp 1604681595
transform 1 0 24184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604681595
transform 1 0 24552 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_266
timestamp 1604681595
transform 1 0 25288 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_270
timestamp 1604681595
transform 1 0 25656 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26576 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_276
timestamp 1604681595
transform 1 0 26208 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3668 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3300 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 3760 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 4864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 5968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9280 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9372 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604681595
transform 1 0 10476 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1604681595
transform 1 0 11580 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1604681595
transform 1 0 12684 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604681595
transform 1 0 13788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 14892 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 14984 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_166
timestamp 1604681595
transform 1 0 16088 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 17652 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16364 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_175
timestamp 1604681595
transform 1 0 16916 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_202
timestamp 1604681595
transform 1 0 19400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_206
timestamp 1604681595
transform 1 0 19768 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20596 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23080 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22528 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22896 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_234
timestamp 1604681595
transform 1 0 22344 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1604681595
transform 1 0 22712 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_261
timestamp 1604681595
transform 1 0 24828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26576 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26116 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1604681595
transform 1 0 25932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26208 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 816 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 816 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1092 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2196 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3668 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3300 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4404 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 3760 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6428 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5508 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6244 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 4864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 5968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7624 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9280 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 8728 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604681595
transform 1 0 9832 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12040 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604681595
transform 1 0 10936 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12132 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604681595
transform 1 0 10476 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604681595
transform 1 0 11580 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1604681595
transform 1 0 13236 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604681595
transform 1 0 12684 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1604681595
transform 1 0 13788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 14892 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1604681595
transform 1 0 14340 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1604681595
transform 1 0 15444 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 14984 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16088 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 17928 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17652 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1604681595
transform 1 0 16548 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1604681595
transform 1 0 17744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17192 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_196
timestamp 1604681595
transform 1 0 18848 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1604681595
transform 1 0 18296 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1604681595
transform 1 0 18572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1604681595
transform 1 0 18204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18940 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18940 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_203
timestamp 1604681595
transform 1 0 19492 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_199
timestamp 1604681595
transform 1 0 19124 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_206
timestamp 1604681595
transform 1 0 19768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 19216 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_211
timestamp 1604681595
transform 1 0 20228 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1604681595
transform 1 0 20136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20596 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20504 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_224
timestamp 1604681595
transform 1 0 21424 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_227
timestamp 1604681595
transform 1 0 21700 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_223
timestamp 1604681595
transform 1 0 21332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_232
timestamp 1604681595
transform 1 0 22160 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_231
timestamp 1604681595
transform 1 0 22068 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22436 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 22252 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_248
timestamp 1604681595
transform 1 0 23632 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_244
timestamp 1604681595
transform 1 0 23264 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 22896 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23264 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23356 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_254
timestamp 1604681595
transform 1 0 24184 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1604681595
transform 1 0 24460 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1604681595
transform 1 0 23908 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 24276 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 24644 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 24276 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_267
timestamp 1604681595
transform 1 0 25380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_263
timestamp 1604681595
transform 1 0 25012 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__89__A
timestamp 1604681595
transform 1 0 25196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604681595
transform 1 0 24644 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26576 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26116 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_275
timestamp 1604681595
transform 1 0 26116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604681595
transform 1 0 25748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26208 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 816 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1092 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2196 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3300 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4404 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6428 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5508 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7624 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 8728 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 9832 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12040 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 10936 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12132 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604681595
transform 1 0 13236 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604681595
transform 1 0 14340 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604681595
transform 1 0 15444 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17652 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604681595
transform 1 0 16548 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_184
timestamp 1604681595
transform 1 0 17744 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18296 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1604681595
transform 1 0 18848 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_200
timestamp 1604681595
transform 1 0 19216 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_208
timestamp 1604681595
transform 1 0 19952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 20136 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 21884 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_213
timestamp 1604681595
transform 1 0 20412 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1604681595
transform 1 0 21516 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23264 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23080 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_232
timestamp 1604681595
transform 1 0 22160 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 22896 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_245
timestamp 1604681595
transform 1 0 23356 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 24276 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 24828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 24092 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_259
timestamp 1604681595
transform 1 0 24644 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_263
timestamp 1604681595
transform 1 0 25012 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_275
timestamp 1604681595
transform 1 0 26116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 816 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3668 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3300 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 3760 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 4864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 5968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9280 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9372 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10476 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11580 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604681595
transform 1 0 13788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 14892 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 14984 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16088 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17192 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18296 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19400 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 20596 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_218
timestamp 1604681595
transform 1 0 20872 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23080 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_230
timestamp 1604681595
transform 1 0 21976 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_248
timestamp 1604681595
transform 1 0 23632 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 24368 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_260
timestamp 1604681595
transform 1 0 24736 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26576 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26116 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_272
timestamp 1604681595
transform 1 0 25840 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26208 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 816 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1092 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2196 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3300 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4404 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6428 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5508 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7624 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 8728 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 9832 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 10936 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12132 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13236 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14340 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15444 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17652 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16548 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 17744 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 18848 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 19952 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21056 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23540 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23264 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_232
timestamp 1604681595
transform 1 0 22160 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 22896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1604681595
transform 1 0 23356 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 24828 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 24368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 25380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_253
timestamp 1604681595
transform 1 0 24092 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_258
timestamp 1604681595
transform 1 0 24552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_265
timestamp 1604681595
transform 1 0 25196 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25564 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26576 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 816 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3668 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3300 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 3760 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 4864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 5968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9280 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9372 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10476 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11580 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12684 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 13788 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 14892 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 14984 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16088 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17192 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18296 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19400 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23080 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_239
timestamp 1604681595
transform 1 0 22804 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_248
timestamp 1604681595
transform 1 0 23632 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 24368 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_260
timestamp 1604681595
transform 1 0 24736 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26576 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26116 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_272
timestamp 1604681595
transform 1 0 25840 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26208 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 816 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1092 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2196 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3300 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4404 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6428 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5508 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6244 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7624 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 8728 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 9832 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12040 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 10936 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12132 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13236 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_147
timestamp 1604681595
transform 1 0 14340 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1604681595
transform 1 0 14892 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1604681595
transform 1 0 15168 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17928 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17652 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_168
timestamp 1604681595
transform 1 0 16272 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1604681595
transform 1 0 17376 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1604681595
transform 1 0 17744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18664 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1604681595
transform 1 0 18480 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 18848 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 19952 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21056 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23264 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22160 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1604681595
transform 1 0 23356 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 24276 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 24828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 24092 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_259
timestamp 1604681595
transform 1 0 24644 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_263
timestamp 1604681595
transform 1 0 25012 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26576 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1604681595
transform 1 0 26116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 816 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 816 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1092 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2196 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3668 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3300 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 3760 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4404 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6428 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 4864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 5968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5508 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9280 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9372 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 8728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1604681595
transform 1 0 9832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_102
timestamp 1604681595
transform 1 0 10200 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12040 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10476 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11580 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1604681595
transform 1 0 11304 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1604681595
transform 1 0 12132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12592 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12684 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 13788 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_127
timestamp 1604681595
transform 1 0 12500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_134
timestamp 1604681595
transform 1 0 13144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_138
timestamp 1604681595
transform 1 0 13512 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14984 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 14892 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 15812 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_160
timestamp 1604681595
transform 1 0 15536 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_150
timestamp 1604681595
transform 1 0 14616 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_162
timestamp 1604681595
transform 1 0 15720 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_165
timestamp 1604681595
transform 1 0 15996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17652 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_172
timestamp 1604681595
transform 1 0 16640 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1604681595
transform 1 0 17744 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_177
timestamp 1604681595
transform 1 0 17100 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 17744 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_196
timestamp 1604681595
transform 1 0 18848 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1604681595
transform 1 0 19952 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 18848 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 19952 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21056 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23264 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 22804 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22160 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1604681595
transform 1 0 23356 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 24276 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 24276 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 24828 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_251
timestamp 1604681595
transform 1 0 23908 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_259
timestamp 1604681595
transform 1 0 24644 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_253
timestamp 1604681595
transform 1 0 24092 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_259
timestamp 1604681595
transform 1 0 24644 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_263
timestamp 1604681595
transform 1 0 25012 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26116 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1604681595
transform 1 0 25748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26208 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_275
timestamp 1604681595
transform 1 0 26116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 816 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3668 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3300 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 3760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 4864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 5968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10016 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9280 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_93
timestamp 1604681595
transform 1 0 9372 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_99
timestamp 1604681595
transform 1 0 9924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_106
timestamp 1604681595
transform 1 0 10568 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_118
timestamp 1604681595
transform 1 0 11672 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_130
timestamp 1604681595
transform 1 0 12776 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_142
timestamp 1604681595
transform 1 0 13880 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 15812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 14892 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1604681595
transform 1 0 14616 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_154
timestamp 1604681595
transform 1 0 14984 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_162
timestamp 1604681595
transform 1 0 15720 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_167
timestamp 1604681595
transform 1 0 16180 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_179
timestamp 1604681595
transform 1 0 17284 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_191
timestamp 1604681595
transform 1 0 18388 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_203
timestamp 1604681595
transform 1 0 19492 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1604681595
transform 1 0 20228 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 22804 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 23908 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25012 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26576 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26116 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26208 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 816 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1092 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2196 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3300 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4404 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6428 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5508 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7624 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 8728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 9832 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12040 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 10936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_112
timestamp 1604681595
transform 1 0 11120 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1604681595
transform 1 0 11856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12132 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13236 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14340 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_161
timestamp 1604681595
transform 1 0 15628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17652 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1604681595
transform 1 0 16732 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1604681595
transform 1 0 17468 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 17744 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 18848 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 19952 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21056 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23356 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23264 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22160 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 24644 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 25196 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24092 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_251
timestamp 1604681595
transform 1 0 23908 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_255
timestamp 1604681595
transform 1 0 24276 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_263
timestamp 1604681595
transform 1 0 25012 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_267
timestamp 1604681595
transform 1 0 25380 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26576 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_275
timestamp 1604681595
transform 1 0 26116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 816 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3668 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 3760 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 4864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 5968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9372 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 10936 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_105
timestamp 1604681595
transform 1 0 10476 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_109
timestamp 1604681595
transform 1 0 10844 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_114
timestamp 1604681595
transform 1 0 11304 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_126
timestamp 1604681595
transform 1 0 12408 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_138
timestamp 1604681595
transform 1 0 13512 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15444 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 14892 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1604681595
transform 1 0 14616 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1604681595
transform 1 0 14984 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_158
timestamp 1604681595
transform 1 0 15352 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1604681595
transform 1 0 15996 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1604681595
transform 1 0 17100 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_189
timestamp 1604681595
transform 1 0 18204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1604681595
transform 1 0 19308 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1604681595
transform 1 0 20412 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 22804 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 23908 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25012 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26576 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26116 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26208 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 816 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1092 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2196 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3300 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4404 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6428 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5508 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6244 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6520 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7624 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 8728 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 9832 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12040 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 10936 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12132 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13236 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14340 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15444 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17652 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16548 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 17744 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 18848 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 19952 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21148 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_220
timestamp 1604681595
transform 1 0 21056 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_223
timestamp 1604681595
transform 1 0 21332 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23264 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1604681595
transform 1 0 22620 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1604681595
transform 1 0 23172 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1604681595
transform 1 0 23356 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 24276 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 24828 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 24092 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_259
timestamp 1604681595
transform 1 0 24644 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_263
timestamp 1604681595
transform 1 0 25012 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26576 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_275
timestamp 1604681595
transform 1 0 26116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 816 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3668 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 3760 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 4864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 5968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9280 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9372 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10476 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12684 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 13788 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 14892 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 14984 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16088 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17192 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18296 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19400 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21148 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1604681595
transform 1 0 20596 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_227
timestamp 1604681595
transform 1 0 21700 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22436 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_241
timestamp 1604681595
transform 1 0 22988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 24276 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1604681595
transform 1 0 24092 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_259
timestamp 1604681595
transform 1 0 24644 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26576 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26116 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1604681595
transform 1 0 25748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26208 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 816 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 816 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1092 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2196 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3668 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3300 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4404 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3300 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 3760 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6428 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5508 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 4864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 5968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7624 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9280 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 8728 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 9832 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9372 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12040 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 10936 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12132 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10476 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11580 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13236 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12684 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 13788 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 14892 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14340 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604681595
transform 1 0 15444 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 14984 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16088 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17652 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16548 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 17744 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17192 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 18848 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 19952 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18296 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19400 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21056 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21700 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_232
timestamp 1604681595
transform 1 0 22160 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_243
timestamp 1604681595
transform 1 0 23172 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1604681595
transform 1 0 22804 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 22896 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23080 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23264 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23264 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 23356 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_250
timestamp 1604681595
transform 1 0 23816 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_249
timestamp 1604681595
transform 1 0 23724 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 24552 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 23908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 24552 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_253
timestamp 1604681595
transform 1 0 24092 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_257
timestamp 1604681595
transform 1 0 24460 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_260
timestamp 1604681595
transform 1 0 24736 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_262
timestamp 1604681595
transform 1 0 24920 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26576 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26576 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26116 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1604681595
transform 1 0 25840 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26208 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26024 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26208 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 816 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1092 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2196 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3300 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4404 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6428 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5508 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6244 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7624 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9464 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_86
timestamp 1604681595
transform 1 0 8728 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_96
timestamp 1604681595
transform 1 0 9648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12040 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_108
timestamp 1604681595
transform 1 0 10752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1604681595
transform 1 0 11856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1604681595
transform 1 0 12132 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_127
timestamp 1604681595
transform 1 0 12500 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1604681595
transform 1 0 13604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14708 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15444 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_157
timestamp 1604681595
transform 1 0 15260 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_161
timestamp 1604681595
transform 1 0 15628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17652 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_173
timestamp 1604681595
transform 1 0 16732 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_181
timestamp 1604681595
transform 1 0 17468 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 17744 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 18848 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 19952 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21056 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23264 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1604681595
transform 1 0 23356 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 24276 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 24828 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 24092 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_259
timestamp 1604681595
transform 1 0 24644 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_263
timestamp 1604681595
transform 1 0 25012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26576 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_275
timestamp 1604681595
transform 1 0 26116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 816 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3668 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3300 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 3760 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 4864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 5968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9464 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9280 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_93
timestamp 1604681595
transform 1 0 9372 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_100
timestamp 1604681595
transform 1 0 10016 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12132 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_112
timestamp 1604681595
transform 1 0 11120 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_120
timestamp 1604681595
transform 1 0 11856 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604681595
transform 1 0 12684 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604681595
transform 1 0 13788 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 14892 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 14984 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604681595
transform 1 0 16088 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604681595
transform 1 0 17192 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604681595
transform 1 0 18296 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19400 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 22804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 24276 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_251
timestamp 1604681595
transform 1 0 23908 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_259
timestamp 1604681595
transform 1 0 24644 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26576 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26116 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1604681595
transform 1 0 25748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26208 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 816 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1092 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2196 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3300 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4404 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6428 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5508 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6244 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7624 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 8728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_98
timestamp 1604681595
transform 1 0 9832 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_104
timestamp 1604681595
transform 1 0 10384 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12040 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 10476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_107
timestamp 1604681595
transform 1 0 10660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_119
timestamp 1604681595
transform 1 0 11764 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12132 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604681595
transform 1 0 13236 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604681595
transform 1 0 14340 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604681595
transform 1 0 15444 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17652 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604681595
transform 1 0 16548 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 17744 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604681595
transform 1 0 18848 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604681595
transform 1 0 19952 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604681595
transform 1 0 21056 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23356 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23264 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23080 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_232
timestamp 1604681595
transform 1 0 22160 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 22896 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 24644 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 24276 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 25196 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1604681595
transform 1 0 23908 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_257
timestamp 1604681595
transform 1 0 24460 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_263
timestamp 1604681595
transform 1 0 25012 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_267
timestamp 1604681595
transform 1 0 25380 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26576 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_275
timestamp 1604681595
transform 1 0 26116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 816 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3668 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3300 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 3760 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 4864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 5968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9280 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9372 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 10476 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1604681595
transform 1 0 10844 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1604681595
transform 1 0 11948 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_133
timestamp 1604681595
transform 1 0 13052 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_145
timestamp 1604681595
transform 1 0 14156 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 14892 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 14984 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16088 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604681595
transform 1 0 17192 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604681595
transform 1 0 18296 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604681595
transform 1 0 19400 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 22804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 24276 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_251
timestamp 1604681595
transform 1 0 23908 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_259
timestamp 1604681595
transform 1 0 24644 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26576 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26116 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1604681595
transform 1 0 25748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26208 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 816 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 816 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1092 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2196 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3668 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4404 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3300 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 3760 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6428 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5508 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6244 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 4864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 5968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7624 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9280 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 8728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 9832 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9372 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12040 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604681595
transform 1 0 10936 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12132 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10476 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11580 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13236 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12684 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 13788 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 14892 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14340 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15444 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 14984 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16088 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17652 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604681595
transform 1 0 16548 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604681595
transform 1 0 17744 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17192 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1604681595
transform 1 0 18848 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1604681595
transform 1 0 19952 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18296 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19400 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1604681595
transform 1 0 21056 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21700 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 23632 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23264 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1604681595
transform 1 0 22160 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604681595
transform 1 0 23356 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_239
timestamp 1604681595
transform 1 0 22804 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_247
timestamp 1604681595
transform 1 0 23540 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 24276 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 24828 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1604681595
transform 1 0 24092 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604681595
transform 1 0 24644 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604681595
transform 1 0 25012 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_252
timestamp 1604681595
transform 1 0 24000 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_264
timestamp 1604681595
transform 1 0 25104 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26576 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26576 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26116 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_272
timestamp 1604681595
transform 1 0 25840 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26208 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 816 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1092 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2196 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4404 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6428 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5508 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6244 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6520 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7624 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 8728 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 9832 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12040 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 10936 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12132 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13236 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14340 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15444 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17652 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16548 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 17744 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 18848 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 19952 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21056 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23264 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22160 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23356 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24460 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25564 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26576 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 816 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1092 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2196 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3668 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3300 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 3760 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6520 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 4864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 5968 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6612 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 7716 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9372 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 8820 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9464 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12224 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10568 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11672 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15076 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14524 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15168 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 17928 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16272 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17376 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18020 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19124 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 20780 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20228 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 20872 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23632 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 21976 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23080 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 23724 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 24828 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26576 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 25932 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 26594 0 26650 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 19234 27520 19290 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 27238 0 27294 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 24846 27520 24902 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 6 0 62 480 6 bottom_left_grid_pin_1_
port 4 nsew default input
rlabel metal2 s 8010 27520 8066 28000 6 ccff_head
port 5 nsew default input
rlabel metal2 s 13622 27520 13678 28000 6 ccff_tail
port 6 nsew default tristate
rlabel metal3 s 27232 4768 27712 4888 6 chanx_right_in[0]
port 7 nsew default input
rlabel metal3 s 27232 10480 27712 10600 6 chanx_right_in[10]
port 8 nsew default input
rlabel metal3 s 27232 11024 27712 11144 6 chanx_right_in[11]
port 9 nsew default input
rlabel metal3 s 27232 11704 27712 11824 6 chanx_right_in[12]
port 10 nsew default input
rlabel metal3 s 27232 12248 27712 12368 6 chanx_right_in[13]
port 11 nsew default input
rlabel metal3 s 27232 12792 27712 12912 6 chanx_right_in[14]
port 12 nsew default input
rlabel metal3 s 27232 13336 27712 13456 6 chanx_right_in[15]
port 13 nsew default input
rlabel metal3 s 27232 13880 27712 14000 6 chanx_right_in[16]
port 14 nsew default input
rlabel metal3 s 27232 14560 27712 14680 6 chanx_right_in[17]
port 15 nsew default input
rlabel metal3 s 27232 15104 27712 15224 6 chanx_right_in[18]
port 16 nsew default input
rlabel metal3 s 27232 15648 27712 15768 6 chanx_right_in[19]
port 17 nsew default input
rlabel metal3 s 27232 5312 27712 5432 6 chanx_right_in[1]
port 18 nsew default input
rlabel metal3 s 27232 5992 27712 6112 6 chanx_right_in[2]
port 19 nsew default input
rlabel metal3 s 27232 6536 27712 6656 6 chanx_right_in[3]
port 20 nsew default input
rlabel metal3 s 27232 7080 27712 7200 6 chanx_right_in[4]
port 21 nsew default input
rlabel metal3 s 27232 7624 27712 7744 6 chanx_right_in[5]
port 22 nsew default input
rlabel metal3 s 27232 8168 27712 8288 6 chanx_right_in[6]
port 23 nsew default input
rlabel metal3 s 27232 8848 27712 8968 6 chanx_right_in[7]
port 24 nsew default input
rlabel metal3 s 27232 9392 27712 9512 6 chanx_right_in[8]
port 25 nsew default input
rlabel metal3 s 27232 9936 27712 10056 6 chanx_right_in[9]
port 26 nsew default input
rlabel metal3 s 27232 16192 27712 16312 6 chanx_right_out[0]
port 27 nsew default tristate
rlabel metal3 s 27232 21904 27712 22024 6 chanx_right_out[10]
port 28 nsew default tristate
rlabel metal3 s 27232 22448 27712 22568 6 chanx_right_out[11]
port 29 nsew default tristate
rlabel metal3 s 27232 23128 27712 23248 6 chanx_right_out[12]
port 30 nsew default tristate
rlabel metal3 s 27232 23672 27712 23792 6 chanx_right_out[13]
port 31 nsew default tristate
rlabel metal3 s 27232 24216 27712 24336 6 chanx_right_out[14]
port 32 nsew default tristate
rlabel metal3 s 27232 24760 27712 24880 6 chanx_right_out[15]
port 33 nsew default tristate
rlabel metal3 s 27232 25304 27712 25424 6 chanx_right_out[16]
port 34 nsew default tristate
rlabel metal3 s 27232 25984 27712 26104 6 chanx_right_out[17]
port 35 nsew default tristate
rlabel metal3 s 27232 26528 27712 26648 6 chanx_right_out[18]
port 36 nsew default tristate
rlabel metal3 s 27232 27072 27712 27192 6 chanx_right_out[19]
port 37 nsew default tristate
rlabel metal3 s 27232 16736 27712 16856 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal3 s 27232 17416 27712 17536 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal3 s 27232 17960 27712 18080 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal3 s 27232 18504 27712 18624 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal3 s 27232 19048 27712 19168 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 27232 19592 27712 19712 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 27232 20272 27712 20392 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 27232 20816 27712 20936 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal3 s 27232 21360 27712 21480 6 chanx_right_out[9]
port 46 nsew default tristate
rlabel metal2 s 650 0 706 480 6 chany_bottom_in[0]
port 47 nsew default input
rlabel metal2 s 7090 0 7146 480 6 chany_bottom_in[10]
port 48 nsew default input
rlabel metal2 s 7734 0 7790 480 6 chany_bottom_in[11]
port 49 nsew default input
rlabel metal2 s 8378 0 8434 480 6 chany_bottom_in[12]
port 50 nsew default input
rlabel metal2 s 9022 0 9078 480 6 chany_bottom_in[13]
port 51 nsew default input
rlabel metal2 s 9758 0 9814 480 6 chany_bottom_in[14]
port 52 nsew default input
rlabel metal2 s 10402 0 10458 480 6 chany_bottom_in[15]
port 53 nsew default input
rlabel metal2 s 11046 0 11102 480 6 chany_bottom_in[16]
port 54 nsew default input
rlabel metal2 s 11690 0 11746 480 6 chany_bottom_in[17]
port 55 nsew default input
rlabel metal2 s 12334 0 12390 480 6 chany_bottom_in[18]
port 56 nsew default input
rlabel metal2 s 12978 0 13034 480 6 chany_bottom_in[19]
port 57 nsew default input
rlabel metal2 s 1294 0 1350 480 6 chany_bottom_in[1]
port 58 nsew default input
rlabel metal2 s 1938 0 1994 480 6 chany_bottom_in[2]
port 59 nsew default input
rlabel metal2 s 2582 0 2638 480 6 chany_bottom_in[3]
port 60 nsew default input
rlabel metal2 s 3226 0 3282 480 6 chany_bottom_in[4]
port 61 nsew default input
rlabel metal2 s 3870 0 3926 480 6 chany_bottom_in[5]
port 62 nsew default input
rlabel metal2 s 4514 0 4570 480 6 chany_bottom_in[6]
port 63 nsew default input
rlabel metal2 s 5158 0 5214 480 6 chany_bottom_in[7]
port 64 nsew default input
rlabel metal2 s 5802 0 5858 480 6 chany_bottom_in[8]
port 65 nsew default input
rlabel metal2 s 6446 0 6502 480 6 chany_bottom_in[9]
port 66 nsew default input
rlabel metal2 s 13622 0 13678 480 6 chany_bottom_out[0]
port 67 nsew default tristate
rlabel metal2 s 20154 0 20210 480 6 chany_bottom_out[10]
port 68 nsew default tristate
rlabel metal2 s 20798 0 20854 480 6 chany_bottom_out[11]
port 69 nsew default tristate
rlabel metal2 s 21442 0 21498 480 6 chany_bottom_out[12]
port 70 nsew default tristate
rlabel metal2 s 22086 0 22142 480 6 chany_bottom_out[13]
port 71 nsew default tristate
rlabel metal2 s 22730 0 22786 480 6 chany_bottom_out[14]
port 72 nsew default tristate
rlabel metal2 s 23374 0 23430 480 6 chany_bottom_out[15]
port 73 nsew default tristate
rlabel metal2 s 24018 0 24074 480 6 chany_bottom_out[16]
port 74 nsew default tristate
rlabel metal2 s 24662 0 24718 480 6 chany_bottom_out[17]
port 75 nsew default tristate
rlabel metal2 s 25306 0 25362 480 6 chany_bottom_out[18]
port 76 nsew default tristate
rlabel metal2 s 25950 0 26006 480 6 chany_bottom_out[19]
port 77 nsew default tristate
rlabel metal2 s 14266 0 14322 480 6 chany_bottom_out[1]
port 78 nsew default tristate
rlabel metal2 s 14910 0 14966 480 6 chany_bottom_out[2]
port 79 nsew default tristate
rlabel metal2 s 15554 0 15610 480 6 chany_bottom_out[3]
port 80 nsew default tristate
rlabel metal2 s 16198 0 16254 480 6 chany_bottom_out[4]
port 81 nsew default tristate
rlabel metal2 s 16842 0 16898 480 6 chany_bottom_out[5]
port 82 nsew default tristate
rlabel metal2 s 17486 0 17542 480 6 chany_bottom_out[6]
port 83 nsew default tristate
rlabel metal2 s 18130 0 18186 480 6 chany_bottom_out[7]
port 84 nsew default tristate
rlabel metal2 s 18866 0 18922 480 6 chany_bottom_out[8]
port 85 nsew default tristate
rlabel metal2 s 19510 0 19566 480 6 chany_bottom_out[9]
port 86 nsew default tristate
rlabel metal2 s 2490 27520 2546 28000 6 prog_clk
port 87 nsew default input
rlabel metal3 s 27232 280 27712 400 6 right_bottom_grid_pin_34_
port 88 nsew default input
rlabel metal3 s 27232 824 27712 944 6 right_bottom_grid_pin_35_
port 89 nsew default input
rlabel metal3 s 27232 1368 27712 1488 6 right_bottom_grid_pin_36_
port 90 nsew default input
rlabel metal3 s 27232 1912 27712 2032 6 right_bottom_grid_pin_37_
port 91 nsew default input
rlabel metal3 s 27232 2456 27712 2576 6 right_bottom_grid_pin_38_
port 92 nsew default input
rlabel metal3 s 27232 3136 27712 3256 6 right_bottom_grid_pin_39_
port 93 nsew default input
rlabel metal3 s 27232 3680 27712 3800 6 right_bottom_grid_pin_40_
port 94 nsew default input
rlabel metal3 s 27232 4224 27712 4344 6 right_bottom_grid_pin_41_
port 95 nsew default input
rlabel metal3 s 27232 27616 27712 27736 6 right_top_grid_pin_1_
port 96 nsew default input
rlabel metal4 s 5323 2128 5643 25616 6 VPWR
port 97 nsew default input
rlabel metal4 s 9989 2128 10309 25616 6 VGND
port 98 nsew default input
<< properties >>
string FIXED_BBOX 1 0 27712 28000
<< end >>
