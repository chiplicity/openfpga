* NGSPICE file created from sb_1__2_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

.subckt sb_1__2_ bottom_left_grid_pin_34_ bottom_left_grid_pin_35_ bottom_left_grid_pin_36_
+ bottom_left_grid_pin_37_ bottom_left_grid_pin_38_ bottom_left_grid_pin_39_ bottom_left_grid_pin_40_
+ bottom_left_grid_pin_41_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_top_grid_pin_1_ prog_clk right_top_grid_pin_1_ vpwr vgnd
Xmem_bottom_track_39.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_39.mux_l1_in_0_/S
+ mux_bottom_track_39.mux_l2_in_0_/S mem_bottom_track_39.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_22_133 vgnd vpwr scs8hd_fill_1
XFILLER_26_85 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_25.scs8hd_buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X _115_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_67 vpwr vgnd scs8hd_fill_2
XFILLER_8_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_25.mux_l3_in_0__A1 mux_left_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_6_107 vpwr vgnd scs8hd_fill_2
XFILLER_6_118 vgnd vpwr scs8hd_decap_4
XFILLER_10_158 vgnd vpwr scs8hd_decap_3
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_87 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 right_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_23_20 vgnd vpwr scs8hd_decap_4
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
X_062_ _062_/HI _062_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_132 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_3__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__D mux_bottom_track_21.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__S mux_bottom_track_7.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_1.mux_l2_in_1_/S mux_left_track_1.mux_l3_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_97 vgnd vpwr scs8hd_decap_4
XFILLER_11_231 vgnd vpwr scs8hd_decap_3
X_045_ _045_/HI _045_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_224 vgnd vpwr scs8hd_fill_1
X_114_ _114_/A chany_bottom_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XFILLER_22_7 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_25.mux_l3_in_0__S mux_bottom_track_25.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_ bottom_left_grid_pin_38_ chanx_right_in[13] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_1__A1 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_20_65 vpwr vgnd scs8hd_fill_2
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D mux_right_track_16.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_29.mux_l2_in_0_ _065_/HI mux_bottom_track_29.mux_l1_in_0_/X mux_bottom_track_29.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_13.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_11.mux_l3_in_0_/S
+ mux_bottom_track_13.mux_l1_in_1_/S mem_bottom_track_13.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_3_271 vgnd vpwr scs8hd_decap_6
XFILLER_6_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l3_in_0__S mux_right_track_16.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.scs8hd_buf_4_0__A mux_left_track_33.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_19.mux_l2_in_0__S mux_bottom_track_19.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_31.mux_l2_in_0_ _067_/HI mux_bottom_track_31.mux_l1_in_0_/X mux_bottom_track_31.mux_l2_in_0_/S
+ mux_bottom_track_31.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_33.scs8hd_buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X _111_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_1_208 vpwr vgnd scs8hd_fill_2
XFILLER_25_142 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vgnd vpwr scs8hd_decap_8
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XFILLER_0_241 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_8
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_33.mux_l3_in_0__A1 mux_left_track_33.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_39.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_37.mux_l2_in_0_/S
+ mux_bottom_track_39.mux_l1_in_0_/S mem_bottom_track_39.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_22_167 vpwr vgnd scs8hd_fill_2
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
XFILLER_22_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_27.scs8hd_buf_4_0__A mux_bottom_track_27.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_116 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_259 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A0 _055_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A1 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_39.mux_l2_in_0__A0 _037_/HI vgnd vpwr scs8hd_diode_2
XFILLER_12_55 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__D mux_bottom_track_7.mux_l1_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_259 vgnd vpwr scs8hd_decap_12
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XFILLER_15_229 vgnd vpwr scs8hd_decap_3
X_061_ _061_/HI _061_/LO vgnd vpwr scs8hd_conb_1
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_9_34 vpwr vgnd scs8hd_fill_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_1.mux_l1_in_1_/S mux_left_track_1.mux_l2_in_1_/S
+ mem_left_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_32 vpwr vgnd scs8hd_fill_2
XFILLER_18_54 vpwr vgnd scs8hd_fill_2
X_113_ _113_/A chany_bottom_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
X_044_ _044_/HI _044_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l3_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_11 vpwr vgnd scs8hd_fill_2
XFILLER_4_206 vgnd vpwr scs8hd_decap_4
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vgnd vpwr scs8hd_fill_1
XFILLER_19_151 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D mux_bottom_track_25.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_15_11 vgnd vpwr scs8hd_decap_3
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_264 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D mux_bottom_track_7.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_29.mux_l1_in_0_ bottom_left_grid_pin_36_ chanx_right_in[11] mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
Xmem_right_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_1_/S
+ mem_right_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_106 vgnd vpwr scs8hd_decap_3
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_31.mux_l1_in_0_ bottom_left_grid_pin_37_ chanx_right_in[7] mux_bottom_track_31.mux_l1_in_0_/S
+ mux_bottom_track_31.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XFILLER_10_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__S mux_bottom_track_23.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_39.mux_l2_in_0__A1 mux_bottom_track_39.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_37_31 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_271 vgnd vpwr scs8hd_decap_4
XFILLER_18_249 vgnd vpwr scs8hd_decap_6
XFILLER_5_131 vpwr vgnd scs8hd_fill_2
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vpwr vgnd scs8hd_fill_2
XFILLER_23_263 vgnd vpwr scs8hd_decap_12
XFILLER_23_66 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_4
X_060_ _060_/HI _060_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_167 vpwr vgnd scs8hd_fill_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
Xmem_left_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l3_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_200 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__D mux_bottom_track_27.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
Xmem_left_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_39.mux_l2_in_0_/S mux_left_track_1.mux_l1_in_1_/S
+ mem_left_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
X_043_ _043_/HI _043_/LO vgnd vpwr scs8hd_conb_1
X_112_ _112_/A chany_bottom_out[15] vgnd vpwr scs8hd_buf_2
Xmem_bottom_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l2_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_4_229 vpwr vgnd scs8hd_fill_2
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_58 vgnd vpwr scs8hd_decap_4
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_174 vpwr vgnd scs8hd_fill_2
XFILLER_19_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D mux_right_track_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_1__A0 _057_/HI vgnd vpwr scs8hd_diode_2
XFILLER_15_56 vpwr vgnd scs8hd_fill_2
XFILLER_15_67 vpwr vgnd scs8hd_fill_2
XFILLER_31_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_25.mux_l2_in_1__S mux_left_track_25.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_276 vgnd vpwr scs8hd_fill_1
XFILLER_0_210 vgnd vpwr scs8hd_fill_1
XFILLER_16_100 vpwr vgnd scs8hd_fill_2
XFILLER_16_144 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_188 vgnd vpwr scs8hd_decap_3
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XFILLER_22_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0__S mux_bottom_track_15.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
Xmem_right_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ mem_right_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_99 vgnd vpwr scs8hd_fill_1
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XFILLER_13_158 vpwr vgnd scs8hd_fill_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A0 mux_bottom_track_13.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.scs8hd_buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _125_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_21.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l2_in_0_/S mem_bottom_track_21.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__D mux_bottom_track_27.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_128 vpwr vgnd scs8hd_fill_2
XFILLER_12_79 vpwr vgnd scs8hd_fill_2
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_37_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XFILLER_23_231 vpwr vgnd scs8hd_fill_2
XFILLER_23_275 vpwr vgnd scs8hd_fill_2
XFILLER_23_56 vpwr vgnd scs8hd_fill_2
XFILLER_23_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_2_179 vgnd vpwr scs8hd_decap_3
XFILLER_2_146 vgnd vpwr scs8hd_fill_1
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_1_/S
+ mem_left_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D mux_right_track_2.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_89 vgnd vpwr scs8hd_decap_3
X_042_ _042_/HI _042_/LO vgnd vpwr scs8hd_conb_1
X_111_ _111_/A chany_bottom_out[16] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_216 vpwr vgnd scs8hd_fill_2
XFILLER_11_245 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_21.mux_l1_in_1__A0 _061_/HI vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_3.mux_l1_in_1_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_109 vgnd vpwr scs8hd_decap_3
XANTENNA__072__A chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_29_11 vgnd vpwr scs8hd_decap_12
XFILLER_20_79 vpwr vgnd scs8hd_fill_2
XFILLER_28_131 vpwr vgnd scs8hd_fill_2
XFILLER_3_263 vpwr vgnd scs8hd_fill_2
XFILLER_3_230 vpwr vgnd scs8hd_fill_2
XFILLER_6_26 vpwr vgnd scs8hd_fill_2
XFILLER_20_7 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_1__A1 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 mux_bottom_track_5.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A0 mux_bottom_track_21.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D mux_left_track_25.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_1_ _054_/HI mux_right_track_8.mux_l1_in_2_/X mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_123 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.scs8hd_buf_4_0_ mux_left_track_9.mux_l3_in_0_/X _083_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_3_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A1 mux_bottom_track_13.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_181 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_21.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/S mem_bottom_track_21.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D mux_right_track_2.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__080__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_2_ chanx_left_in[16] chanx_left_in[6] mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_55 vgnd vpwr scs8hd_decap_6
XFILLER_18_218 vpwr vgnd scs8hd_fill_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_5_144 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_70 vgnd vpwr scs8hd_fill_1
XFILLER_23_243 vgnd vpwr scs8hd_fill_1
XFILLER_23_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_125 vgnd vpwr scs8hd_decap_4
XFILLER_0_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_210 vgnd vpwr scs8hd_fill_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_35.scs8hd_buf_4_0__A mux_bottom_track_35.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_5.mux_l3_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_68 vpwr vgnd scs8hd_fill_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A chany_bottom_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_257 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
X_041_ _041_/HI _041_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_21.mux_l1_in_1__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2__A0 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_23 vgnd vpwr scs8hd_decap_12
XFILLER_20_69 vgnd vpwr scs8hd_fill_1
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_80 vpwr vgnd scs8hd_fill_2
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_25_146 vpwr vgnd scs8hd_fill_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 mux_bottom_track_5.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A1 mux_bottom_track_21.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 _054_/HI vgnd vpwr scs8hd_diode_2
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
XFILLER_22_116 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_29.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/S mem_bottom_track_29.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_142 vpwr vgnd scs8hd_fill_2
XFILLER_8_186 vgnd vpwr scs8hd_decap_3
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XFILLER_12_59 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_1_ chany_bottom_in[16] chany_bottom_in[9] mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__S mux_bottom_track_11.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_112 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_38 vgnd vpwr scs8hd_decap_4
XFILLER_14_233 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_20_247 vgnd vpwr scs8hd_decap_8
XFILLER_20_236 vgnd vpwr scs8hd_decap_8
XFILLER_9_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__D mux_bottom_track_9.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_58 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_203 vgnd vpwr scs8hd_decap_3
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_269 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
X_040_ _040_/HI _040_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__D mux_bottom_track_29.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2__A1 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_35 vgnd vpwr scs8hd_decap_12
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XFILLER_28_144 vpwr vgnd scs8hd_fill_2
XFILLER_19_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D mux_right_track_24.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XFILLER_24_191 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 mux_right_track_8.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_39.scs8hd_buf_4_0_ mux_bottom_track_39.mux_l2_in_0_/X _108_/A vgnd
+ vpwr scs8hd_buf_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_150 vgnd vpwr scs8hd_decap_3
XANTENNA__094__A chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chanx_right_in[19] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_ mux_bottom_track_13.mux_l1_in_1_/X mux_bottom_track_13.mux_l1_in_0_/X
+ mux_bottom_track_13.mux_l2_in_0_/S mux_bottom_track_13.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_3_29 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_29.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/S mem_bottom_track_29.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_194 vgnd vpwr scs8hd_decap_3
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A mux_bottom_track_17.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_0_ chany_bottom_in[2] right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D mux_right_track_8.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_3__A0 _039_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__089__A chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_17_264 vgnd vpwr scs8hd_decap_12
XFILLER_4_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_245 vpwr vgnd scs8hd_fill_2
XFILLER_23_26 vpwr vgnd scs8hd_fill_2
XFILLER_3_7 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_13.mux_l1_in_1_ _057_/HI chanx_left_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.mux_l2_in_1_ _063_/HI chanx_left_in[18] mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_171 vpwr vgnd scs8hd_fill_2
XFILLER_20_204 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S mux_bottom_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XFILLER_18_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_099_ _099_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_47 vgnd vpwr scs8hd_decap_12
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XANTENNA__097__A chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_3_222 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_1_ _040_/HI chanx_left_in[15] mux_bottom_track_9.mux_l2_in_1_/S
+ mux_bottom_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_60 vgnd vpwr scs8hd_decap_4
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
XFILLER_19_178 vgnd vpwr scs8hd_decap_3
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_37.mux_l1_in_0__S mux_bottom_track_37.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l3_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_148 vgnd vpwr scs8hd_decap_4
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 _044_/HI vgnd vpwr scs8hd_diode_2
XFILLER_22_129 vgnd vpwr scs8hd_decap_4
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_72 vpwr vgnd scs8hd_fill_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
XFILLER_21_162 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_140 vgnd vpwr scs8hd_decap_4
XFILLER_12_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_7.mux_l1_in_3__A1 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A mux_bottom_track_5.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_11.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_11.mux_l2_in_1_/S
+ mux_bottom_track_11.mux_l3_in_0_/S mem_bottom_track_11.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_17_221 vpwr vgnd scs8hd_fill_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_4.scs8hd_buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _105_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_4_180 vpwr vgnd scs8hd_fill_2
XFILLER_4_73 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D mux_left_track_1.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_235 vgnd vpwr scs8hd_decap_8
XFILLER_23_16 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_ bottom_left_grid_pin_36_ chanx_right_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_33.mux_l3_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_224 vgnd vpwr scs8hd_decap_3
XFILLER_13_93 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.mux_l2_in_0_ bottom_left_grid_pin_34_ mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S mux_bottom_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l1_in_1__S mux_bottom_track_13.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__D mux_bottom_track_15.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_17.mux_l2_in_1_/S mux_left_track_17.mux_l3_in_0_/S
+ mem_left_track_17.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_29.mux_l2_in_0__S mux_bottom_track_29.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 _052_/HI vgnd vpwr scs8hd_diode_2
X_098_ chanx_left_in[8] chanx_right_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_1_30 vpwr vgnd scs8hd_fill_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__D mux_bottom_track_35.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_102 vgnd vpwr scs8hd_decap_3
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_245 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l2_in_0_ chanx_left_in[8] mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S mux_bottom_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_267 vpwr vgnd scs8hd_fill_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.scs8hd_buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X _121_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_15_39 vpwr vgnd scs8hd_fill_2
XFILLER_0_237 vgnd vpwr scs8hd_decap_4
Xmem_right_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_16.mux_l1_in_1_/S mux_right_track_16.mux_l2_in_1_/S
+ mem_right_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 mux_right_track_32.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_127 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_19.mux_l1_in_1__A0 _060_/HI vgnd vpwr scs8hd_diode_2
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D mux_left_track_3.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_174 vpwr vgnd scs8hd_fill_2
XFILLER_8_101 vpwr vgnd scs8hd_fill_2
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A0 mux_bottom_track_19.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D mux_bottom_track_15.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_148 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_11.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l2_in_1_/S mem_bottom_track_11.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__D mux_bottom_track_35.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_192 vgnd vpwr scs8hd_decap_3
XFILLER_23_214 vgnd vpwr scs8hd_decap_12
XFILLER_23_203 vpwr vgnd scs8hd_fill_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_fill_1
XFILLER_14_236 vpwr vgnd scs8hd_fill_2
XFILLER_13_72 vpwr vgnd scs8hd_fill_2
XFILLER_1_140 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_37.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_37.mux_l1_in_0_/S
+ mux_bottom_track_37.mux_l2_in_0_/S mem_bottom_track_37.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_17.mux_l1_in_1_/S mux_left_track_17.mux_l2_in_1_/S
+ mem_left_track_17.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_8.mux_l1_in_2__S mux_right_track_8.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_8
XFILLER_6_210 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_221 vpwr vgnd scs8hd_fill_2
XFILLER_6_254 vpwr vgnd scs8hd_fill_2
XFILLER_6_265 vgnd vpwr scs8hd_decap_8
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
X_097_ chanx_left_in[9] chanx_right_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_21.scs8hd_buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X _117_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D mux_left_track_3.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l1_in_0_ chanx_right_in[19] chanx_right_in[18] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_147 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_103 vpwr vgnd scs8hd_fill_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_4
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_37.mux_l2_in_0_ _036_/HI mux_bottom_track_37.mux_l1_in_0_/X mux_bottom_track_37.mux_l2_in_0_/S
+ mux_bottom_track_37.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_25_117 vgnd vpwr scs8hd_decap_3
XFILLER_31_17 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_0_249 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_8.mux_l3_in_0_/S mux_right_track_16.mux_l1_in_1_/S
+ mem_right_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_19.mux_l1_in_1__A1 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 right_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_11_8 vpwr vgnd scs8hd_fill_2
XFILLER_30_142 vgnd vpwr scs8hd_decap_8
XFILLER_30_131 vgnd vpwr scs8hd_decap_3
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A0 _064_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D mux_left_track_33.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_197 vgnd vpwr scs8hd_decap_4
XFILLER_21_131 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_34_ chanx_right_in[8] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_16_83 vgnd vpwr scs8hd_decap_8
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_124 vgnd vpwr scs8hd_decap_3
XFILLER_8_146 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A1 mux_bottom_track_19.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_127 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l2_in_1_ _044_/HI chany_bottom_in[14] mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_11.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_9.mux_l3_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/S mem_bottom_track_11.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_17_234 vpwr vgnd scs8hd_fill_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_259 vpwr vgnd scs8hd_fill_2
XFILLER_23_226 vpwr vgnd scs8hd_fill_2
XFILLER_14_259 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
XFILLER_9_230 vpwr vgnd scs8hd_fill_2
XFILLER_13_270 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_37.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_35.mux_l2_in_0_/S
+ mux_bottom_track_37.mux_l1_in_0_/S mem_bottom_track_37.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
Xmem_right_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A mux_bottom_track_25.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_9.mux_l3_in_0_/S mux_left_track_17.mux_l1_in_1_/S
+ mem_left_track_17.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ chanx_left_in[10] chanx_right_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_20_19 vpwr vgnd scs8hd_fill_2
XFILLER_28_148 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.mux_l1_in_1__S mux_bottom_track_7.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_10_41 vgnd vpwr scs8hd_decap_3
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_35.mux_l2_in_0__A0 _035_/HI vgnd vpwr scs8hd_diode_2
X_079_ _079_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_25_129 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_29 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_206 vgnd vpwr scs8hd_decap_4
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_62 vgnd vpwr scs8hd_decap_3
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_140 vpwr vgnd scs8hd_fill_2
XFILLER_15_184 vgnd vpwr scs8hd_fill_1
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__S mux_bottom_track_19.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A1 mux_bottom_track_27.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_154 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_37.mux_l1_in_0_ bottom_left_grid_pin_40_ chanx_right_in[0] mux_bottom_track_37.mux_l1_in_0_/S
+ mux_bottom_track_37.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_62 vgnd vpwr scs8hd_decap_4
XFILLER_16_73 vgnd vpwr scs8hd_fill_1
XFILLER_8_158 vpwr vgnd scs8hd_fill_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l3_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_bottom_track_19.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l2_in_0_/S mem_bottom_track_19.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
Xmem_right_track_24.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l3_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_87 vpwr vgnd scs8hd_fill_2
XFILLER_23_249 vgnd vpwr scs8hd_decap_4
XFILLER_22_271 vgnd vpwr scs8hd_decap_4
XFILLER_13_52 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XFILLER_20_208 vgnd vpwr scs8hd_decap_6
Xmem_right_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_3.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_208 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l2_in_1_ _049_/HI chanx_left_in[17] mux_right_track_16.mux_l2_in_1_/S
+ mux_right_track_16.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
Xmux_right_track_4.mux_l2_in_1_ _053_/HI mux_right_track_4.mux_l1_in_2_/X mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
X_095_ _095_/A chanx_right_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A0 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_259 vpwr vgnd scs8hd_fill_2
XFILLER_3_226 vpwr vgnd scs8hd_fill_2
XFILLER_10_64 vgnd vpwr scs8hd_fill_1
XFILLER_10_97 vgnd vpwr scs8hd_fill_1
XFILLER_27_160 vgnd vpwr scs8hd_decap_12
XFILLER_19_73 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_35.mux_l2_in_0__A1 mux_bottom_track_35.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
X_078_ chanx_right_in[8] chanx_left_out[9] vgnd vpwr scs8hd_buf_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_193 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_2_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_174 vgnd vpwr scs8hd_decap_12
XFILLER_24_163 vpwr vgnd scs8hd_fill_2
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D mux_left_track_17.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_152 vpwr vgnd scs8hd_fill_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
Xmem_left_track_25.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_25.mux_l2_in_1_/S mux_left_track_25.mux_l3_in_0_/S
+ mem_left_track_25.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_32 vpwr vgnd scs8hd_fill_2
XFILLER_7_65 vgnd vpwr scs8hd_decap_4
XFILLER_26_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vpwr vgnd scs8hd_fill_2
XFILLER_12_144 vgnd vpwr scs8hd_fill_1
XFILLER_12_177 vpwr vgnd scs8hd_fill_2
XFILLER_12_199 vgnd vpwr scs8hd_decap_3
XFILLER_16_96 vpwr vgnd scs8hd_fill_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l2_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_bottom_track_19.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l1_in_1_/S mem_bottom_track_19.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_26_247 vgnd vpwr scs8hd_decap_8
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
Xmem_right_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_24.mux_l1_in_1_/S mux_right_track_24.mux_l2_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_184 vpwr vgnd scs8hd_fill_2
XFILLER_4_66 vgnd vpwr scs8hd_decap_4
XFILLER_4_22 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l1_in_1__S mux_right_track_32.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_4
XFILLER_13_31 vpwr vgnd scs8hd_fill_2
XFILLER_13_97 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_3.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_right_track_0.mux_l1_in_1_/S
+ mem_right_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
X_094_ chanx_left_in[12] chanx_right_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A1 mux_left_track_33.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_205 vpwr vgnd scs8hd_fill_2
XFILLER_10_21 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.scs8hd_buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _127_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_172 vgnd vpwr scs8hd_decap_8
XFILLER_19_52 vgnd vpwr scs8hd_decap_6
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2__A0 left_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
X_077_ chanx_right_in[9] chanx_left_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_153 vgnd vpwr scs8hd_decap_12
XFILLER_33_131 vgnd vpwr scs8hd_fill_1
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_ chanx_left_in[8] chany_bottom_in[15] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_ chany_bottom_in[17] chany_bottom_in[10] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_186 vpwr vgnd scs8hd_fill_2
XFILLER_24_131 vpwr vgnd scs8hd_fill_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_86 vgnd vpwr scs8hd_decap_6
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_39.mux_l1_in_0__A0 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
Xmem_left_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_25.mux_l1_in_1_/S mux_left_track_25.mux_l2_in_1_/S
+ mem_left_track_25.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
XFILLER_21_178 vgnd vpwr scs8hd_decap_3
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_21_112 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 _047_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D mux_bottom_track_3.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__S mux_bottom_track_21.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_9.mux_l2_in_1_/S mux_bottom_track_9.mux_l3_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_32_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_32.mux_l2_in_0_/S mux_bottom_track_1.mux_l1_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_37_19 vgnd vpwr scs8hd_decap_12
XFILLER_26_259 vgnd vpwr scs8hd_decap_12
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0__S mux_bottom_track_15.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D mux_right_track_8.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_25_270 vgnd vpwr scs8hd_decap_6
Xmem_right_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_16.mux_l3_in_0_/S mux_right_track_24.mux_l1_in_1_/S
+ mem_right_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_229 vgnd vpwr scs8hd_decap_4
XFILLER_13_65 vgnd vpwr scs8hd_decap_4
XFILLER_1_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 mux_bottom_track_1.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_222 vpwr vgnd scs8hd_fill_2
XFILLER_9_266 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_8.mux_l1_in_1_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_210 vpwr vgnd scs8hd_fill_2
X_093_ chanx_left_in[13] chanx_right_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_6_225 vpwr vgnd scs8hd_fill_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_24 vgnd vpwr scs8hd_decap_4
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_79 vgnd vpwr scs8hd_decap_3
Xmux_left_track_5.scs8hd_buf_4_0_ mux_left_track_5.mux_l3_in_0_/X _085_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__D mux_bottom_track_23.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_107 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l1_in_3_ _038_/HI chanx_left_in[7] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vpwr vgnd scs8hd_fill_2
XFILLER_19_31 vpwr vgnd scs8hd_fill_2
XFILLER_10_88 vgnd vpwr scs8hd_fill_1
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_19_86 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2__A1 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_32_7 vgnd vpwr scs8hd_decap_8
X_076_ chanx_right_in[10] chanx_left_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_140 vpwr vgnd scs8hd_fill_2
XFILLER_33_165 vgnd vpwr scs8hd_decap_12
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_ chany_bottom_in[8] chany_bottom_in[1] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_4.mux_l1_in_0_ chany_bottom_in[3] right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_19.scs8hd_buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X _118_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_39.mux_l1_in_0__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_30_102 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_left_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_1_/S
+ mem_left_track_25.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A mux_bottom_track_33.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_12 vpwr vgnd scs8hd_fill_2
XFILLER_7_45 vpwr vgnd scs8hd_fill_2
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
X_059_ _059_/HI _059_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 mux_left_track_9.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_9.mux_l1_in_0_/S mux_bottom_track_9.mux_l2_in_1_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_34_271 vgnd vpwr scs8hd_decap_4
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_17_238 vgnd vpwr scs8hd_decap_4
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D mux_bottom_track_23.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_230 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__D mux_bottom_track_7.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_44 vpwr vgnd scs8hd_fill_2
XFILLER_1_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmem_right_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_4.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_1_/S
+ mem_right_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 _053_/HI vgnd vpwr scs8hd_diode_2
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
XFILLER_6_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_244 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_27.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/S mem_bottom_track_27.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_6_248 vgnd vpwr scs8hd_decap_4
X_092_ chanx_left_in[14] chanx_right_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_27.scs8hd_buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X _114_/A vgnd
+ vpwr scs8hd_buf_1
Xmux_bottom_track_5.mux_l1_in_2_ chanx_left_in[5] bottom_left_grid_pin_40_ mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_67 vpwr vgnd scs8hd_fill_2
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_075_ _075_/A chanx_left_out[12] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_240 vpwr vgnd scs8hd_fill_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XFILLER_33_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_11 vpwr vgnd scs8hd_fill_2
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XFILLER_30_136 vgnd vpwr scs8hd_decap_3
XFILLER_30_114 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_5.scs8hd_buf_4_0__A mux_left_track_5.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_144 vgnd vpwr scs8hd_fill_1
X_127_ _127_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
X_058_ _058_/HI _058_/LO vgnd vpwr scs8hd_conb_1
XFILLER_21_158 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_19.mux_l2_in_0_ mux_bottom_track_19.mux_l1_in_1_/X mux_bottom_track_19.mux_l1_in_0_/X
+ mux_bottom_track_19.mux_l2_in_0_/S mux_bottom_track_19.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_9.mux_l1_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_125 vpwr vgnd scs8hd_fill_2
XFILLER_12_136 vpwr vgnd scs8hd_fill_2
XFILLER_12_147 vgnd vpwr scs8hd_decap_3
XFILLER_16_66 vgnd vpwr scs8hd_fill_1
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_129 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_21.mux_l2_in_0_ mux_bottom_track_21.mux_l1_in_1_/X mux_bottom_track_21.mux_l1_in_0_/X
+ mux_bottom_track_21.mux_l2_in_0_/S mux_bottom_track_21.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_7_162 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vgnd vpwr scs8hd_fill_1
XFILLER_26_239 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_217 vpwr vgnd scs8hd_fill_2
XFILLER_4_132 vpwr vgnd scs8hd_fill_2
XFILLER_4_36 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_19.mux_l1_in_1_ _060_/HI chanx_left_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_1__A0 _056_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_1__S mux_bottom_track_23.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_33.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_33.mux_l2_in_1_/S ccff_tail
+ mem_left_track_33.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_21.mux_l1_in_1_ _061_/HI chanx_left_in[16] mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_56 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.mux_l1_in_0__S mux_bottom_track_11.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_39.mux_l2_in_0__S mux_bottom_track_39.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_35.scs8hd_buf_4_0_ mux_bottom_track_35.mux_l2_in_0_/X _110_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_091_ _091_/A chanx_right_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_10_234 vpwr vgnd scs8hd_fill_2
XFILLER_10_267 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_27.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/S mem_bottom_track_27.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l3_in_0__A0 mux_bottom_track_11.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A0 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.scs8hd_buf_4_0__A mux_bottom_track_15.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_32.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_32.mux_l1_in_1_/S mux_right_track_32.mux_l2_in_0_/S
+ mem_right_track_32.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_38_ bottom_left_grid_pin_36_
+ mux_bottom_track_5.mux_l1_in_0_/S mux_bottom_track_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_46 vgnd vpwr scs8hd_decap_3
XFILLER_27_153 vgnd vpwr scs8hd_decap_4
XFILLER_19_66 vgnd vpwr scs8hd_fill_1
XFILLER_19_11 vgnd vpwr scs8hd_decap_3
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_074_ chanx_right_in[12] chanx_left_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A0 _066_/HI vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 mux_bottom_track_5.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_167 vpwr vgnd scs8hd_fill_2
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XFILLER_24_101 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.scs8hd_buf_4_0__A mux_right_track_4.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_23 vgnd vpwr scs8hd_decap_4
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_7_69 vgnd vpwr scs8hd_fill_1
X_126_ _126_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_057_ _057_/HI _057_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l3_in_0__S mux_bottom_track_7.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_45 vpwr vgnd scs8hd_fill_2
X_109_ _109_/A chany_bottom_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_4
XFILLER_27_11 vpwr vgnd scs8hd_fill_2
XANTENNA__070__A chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_188 vpwr vgnd scs8hd_fill_2
XFILLER_4_26 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_19.mux_l1_in_0_ bottom_left_grid_pin_39_ chanx_right_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_1__A1 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_1_/S
+ mem_left_track_33.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__D mux_bottom_track_29.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_21.mux_l1_in_0_ bottom_left_grid_pin_40_ chanx_right_in[16] mux_bottom_track_21.mux_l1_in_0_/S
+ mux_bottom_track_21.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_103 vgnd vpwr scs8hd_decap_3
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_33.mux_l2_in_0_ _034_/HI mux_bottom_track_33.mux_l1_in_0_/X mux_bottom_track_33.mux_l2_in_0_/S
+ mux_bottom_track_33.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_236 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_67 vgnd vpwr scs8hd_decap_8
XFILLER_24_56 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_6_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_11.mux_l3_in_0__A1 mux_bottom_track_11.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
X_090_ chanx_left_in[16] chanx_right_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_6_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A1 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_5_261 vpwr vgnd scs8hd_fill_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D mux_right_track_2.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_32.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_24.mux_l3_in_0_/S mux_right_track_32.mux_l1_in_1_/S
+ mem_right_track_32.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_3_209 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_34_ chanx_right_in[5] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_25 vgnd vpwr scs8hd_decap_4
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A mux_bottom_track_3.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_073_ chanx_right_in[13] chanx_left_out[14] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_121 vgnd vpwr scs8hd_decap_8
XFILLER_18_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.scs8hd_buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _107_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_24_135 vgnd vpwr scs8hd_fill_1
XFILLER_24_124 vgnd vpwr scs8hd_decap_4
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA__073__A chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_15_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 mux_right_track_8.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
X_125_ _125_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_30_7 vgnd vpwr scs8hd_decap_12
X_056_ _056_/HI _056_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_21_127 vpwr vgnd scs8hd_fill_2
XFILLER_21_116 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__068__A chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D mux_left_track_25.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
X_108_ _108_/A chany_bottom_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
X_039_ _039_/HI _039_/LO vgnd vpwr scs8hd_conb_1
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
XFILLER_4_101 vpwr vgnd scs8hd_fill_2
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_4_49 vpwr vgnd scs8hd_fill_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
Xmem_left_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ mem_left_track_33.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D mux_right_track_4.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_69 vgnd vpwr scs8hd_fill_1
XANTENNA__081__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_226 vpwr vgnd scs8hd_fill_2
XFILLER_13_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_1__A0 _058_/HI vgnd vpwr scs8hd_diode_2
XFILLER_5_81 vpwr vgnd scs8hd_fill_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XANTENNA__076__A chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_35.mux_l2_in_0__S mux_bottom_track_35.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_35 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_33.mux_l1_in_0_ bottom_left_grid_pin_38_ chanx_right_in[3] mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
X_072_ chanx_right_in[14] chanx_left_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_2_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A0 mux_bottom_track_15.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_7.scs8hd_buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X _124_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_29.mux_l1_in_0__S mux_bottom_track_29.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_144 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_1_ _042_/HI chany_bottom_in[17] mux_left_track_17.mux_l2_in_1_/S
+ mux_left_track_17.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_93 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_191 vgnd vpwr scs8hd_decap_4
X_124_ _124_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_055_ _055_/HI _055_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_16 vpwr vgnd scs8hd_fill_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_3
XFILLER_7_49 vpwr vgnd scs8hd_fill_2
XFILLER_23_7 vgnd vpwr scs8hd_fill_1
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_35.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_35.mux_l1_in_0_/S
+ mux_bottom_track_35.mux_l2_in_0_/S mem_bottom_track_35.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_16_58 vpwr vgnd scs8hd_fill_2
XFILLER_16_69 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_183 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_107_ _107_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_038_ _038_/HI _038_/LO vgnd vpwr scs8hd_conb_1
XFILLER_26_209 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l2_in_1_ _047_/HI mux_left_track_9.mux_l1_in_2_/X mux_left_track_9.mux_l2_in_1_/S
+ mux_left_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_70 vgnd vpwr scs8hd_fill_1
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A0 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_1_ _048_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_1__A0 _062_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_90 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XFILLER_13_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D mux_right_track_16.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_48 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_25.mux_l3_in_0__S mux_left_track_25.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_1__S mux_bottom_track_11.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_205 vpwr vgnd scs8hd_fill_2
XFILLER_13_223 vpwr vgnd scs8hd_fill_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_2_ left_top_grid_pin_1_ chany_bottom_in[16] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_15.mux_l1_in_1__A1 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A0 mux_bottom_track_7.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_ chanx_left_in[12] chanx_left_in[2] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_36 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A0 mux_bottom_track_23.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__D mux_bottom_track_11.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_69 vpwr vgnd scs8hd_fill_2
XFILLER_19_58 vgnd vpwr scs8hd_fill_1
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_071_ _071_/A chanx_left_out[16] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A1 mux_bottom_track_15.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A0 mux_bottom_track_7.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_101 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__D mux_bottom_track_31.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_189 vpwr vgnd scs8hd_fill_2
XFILLER_24_104 vgnd vpwr scs8hd_fill_1
XFILLER_2_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_1_/S mux_left_track_17.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_148 vpwr vgnd scs8hd_fill_2
X_123_ _123_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
X_054_ _054_/HI _054_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 mux_left_track_3.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_35.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_33.mux_l2_in_0_/S
+ mux_bottom_track_35.mux_l1_in_0_/S mem_bottom_track_35.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_23.scs8hd_buf_4_0__A mux_bottom_track_23.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_4
X_106_ _106_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_22_80 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_ chany_bottom_in[10] chany_bottom_in[3] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_037_ _037_/HI _037_/LO vgnd vpwr scs8hd_conb_1
XFILLER_19_240 vgnd vpwr scs8hd_decap_4
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_93 vgnd vpwr scs8hd_fill_1
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_276 vgnd vpwr scs8hd_fill_1
XFILLER_25_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_23.mux_l1_in_1__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_16_210 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_31.mux_l2_in_0__A0 _067_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__D mux_bottom_track_11.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D mux_right_track_8.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_ chany_bottom_in[9] chany_bottom_in[2] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_28_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D mux_bottom_track_31.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A1 mux_bottom_track_7.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_24_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A1 mux_bottom_track_23.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_ chany_bottom_in[19] chany_bottom_in[12] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_48 vgnd vpwr scs8hd_decap_8
XFILLER_10_238 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_24.mux_l2_in_1_ _051_/HI chanx_left_in[18] mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_220 vpwr vgnd scs8hd_fill_2
XFILLER_5_231 vgnd vpwr scs8hd_fill_1
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l2_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_48 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
X_070_ chanx_right_in[16] chanx_left_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_201 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A1 mux_bottom_track_7.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_157 vgnd vpwr scs8hd_decap_6
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_2_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_149 vpwr vgnd scs8hd_fill_2
XFILLER_21_27 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D mux_bottom_track_39.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_31.mux_l2_in_0__S mux_bottom_track_31.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__098__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_23_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
X_122_ _122_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
X_053_ _053_/HI _053_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_182 vpwr vgnd scs8hd_fill_2
XFILLER_37_252 vgnd vpwr scs8hd_decap_3
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_119 vgnd vpwr scs8hd_decap_4
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
X_105_ _105_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_7_112 vpwr vgnd scs8hd_fill_2
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
XFILLER_7_156 vgnd vpwr scs8hd_decap_4
XFILLER_7_189 vpwr vgnd scs8hd_fill_2
X_036_ _036_/HI _036_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_17.mux_l1_in_0_ chanx_right_in[17] chanx_right_in[8] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_83 vpwr vgnd scs8hd_fill_2
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_31.mux_l2_in_0__A1 mux_bottom_track_31.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_247 vgnd vpwr scs8hd_decap_8
XFILLER_22_236 vgnd vpwr scs8hd_decap_8
XFILLER_22_203 vgnd vpwr scs8hd_decap_8
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_3_ _055_/HI chanx_left_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_203 vpwr vgnd scs8hd_fill_2
XFILLER_13_236 vgnd vpwr scs8hd_decap_4
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_8
Xmem_left_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l3_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_3__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_273 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_ chany_bottom_in[5] right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vpwr vgnd scs8hd_fill_2
XFILLER_6_7 vpwr vgnd scs8hd_fill_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_60 vgnd vpwr scs8hd_decap_4
XFILLER_5_265 vpwr vgnd scs8hd_fill_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/S mem_bottom_track_17.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_224 vpwr vgnd scs8hd_fill_2
XFILLER_18_169 vgnd vpwr scs8hd_fill_1
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vpwr vgnd scs8hd_fill_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_128 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_24.mux_l1_in_1_ chanx_left_in[9] chany_bottom_in[14] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_180 vgnd vpwr scs8hd_decap_3
XFILLER_17_191 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_23_161 vpwr vgnd scs8hd_fill_2
X_121_ _121_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A1 chanx_right_in[14] vgnd vpwr scs8hd_diode_2
X_052_ _052_/HI _052_/LO vgnd vpwr scs8hd_conb_1
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_104_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_035_ _035_/HI _035_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_135 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_142 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_8_73 vgnd vpwr scs8hd_fill_1
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A0 _063_/HI vgnd vpwr scs8hd_diode_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D mux_left_track_3.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_105 vpwr vgnd scs8hd_fill_2
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_234 vpwr vgnd scs8hd_fill_2
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_3_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_22_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_108 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_2_ chanx_left_in[1] bottom_left_grid_pin_40_ mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A0 mux_bottom_track_25.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_5.mux_l1_in_2_/S mux_left_track_5.mux_l2_in_1_/S
+ mem_left_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_30 vpwr vgnd scs8hd_fill_2
XFILLER_5_85 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_35.mux_l1_in_0__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__D mux_bottom_track_37.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_7.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l3_in_0_/S
+ mem_bottom_track_7.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_14_83 vpwr vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 _046_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chanx_right_in[18] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l2_in_0_ mux_bottom_track_15.mux_l1_in_1_/X mux_bottom_track_15.mux_l1_in_0_/X
+ mux_bottom_track_15.mux_l2_in_0_/S mux_bottom_track_15.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A1 chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_2_236 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_18_148 vpwr vgnd scs8hd_fill_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_24.mux_l1_in_0_ chany_bottom_in[7] chany_bottom_in[0] mux_right_track_24.mux_l1_in_1_/S
+ mux_right_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D mux_left_track_5.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_195 vgnd vpwr scs8hd_fill_1
X_051_ _051_/HI _051_/LO vgnd vpwr scs8hd_conb_1
X_120_ _120_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_11_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.scs8hd_buf_4_0__A mux_right_track_16.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_1_ _058_/HI chanx_left_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_195 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_187 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_20_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__D mux_bottom_track_17.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l3_in_0_/S mem_bottom_track_25.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _103_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_034_ _034_/HI _034_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_221 vgnd vpwr scs8hd_decap_12
XFILLER_19_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__D mux_bottom_track_37.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.scs8hd_buf_4_0_ mux_left_track_1.mux_l3_in_0_/X _087_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D mux_left_track_33.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__S mux_bottom_track_21.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_257 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_38_ bottom_left_grid_pin_36_
+ mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_31.scs8hd_buf_4_0__A mux_bottom_track_31.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_0_175 vgnd vpwr scs8hd_decap_4
XFILLER_28_93 vgnd vpwr scs8hd_decap_6
Xmem_left_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_3.mux_l3_in_0_/S mux_left_track_5.mux_l1_in_2_/S
+ mem_left_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A1 mux_bottom_track_25.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_242 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.scs8hd_buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X _120_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_35.mux_l1_in_0__A1 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_5_20 vgnd vpwr scs8hd_decap_3
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_7.mux_l1_in_2_/S mux_bottom_track_7.mux_l2_in_1_/S
+ mem_bottom_track_7.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_4
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_149 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_98 vpwr vgnd scs8hd_fill_2
XFILLER_2_76 vpwr vgnd scs8hd_fill_2
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XFILLER_21_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_174 vpwr vgnd scs8hd_fill_2
XFILLER_23_130 vpwr vgnd scs8hd_fill_2
X_050_ _050_/HI _050_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_7.mux_l1_in_2__S mux_bottom_track_7.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XFILLER_11_74 vpwr vgnd scs8hd_fill_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l1_in_0_ bottom_left_grid_pin_37_ chanx_right_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__S mux_bottom_track_25.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_18 vgnd vpwr scs8hd_decap_12
XFILLER_20_122 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_27.mux_l2_in_0_ _064_/HI mux_bottom_track_27.mux_l1_in_0_/X mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0__S mux_bottom_track_13.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 _048_/HI vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l2_in_1_/S mem_bottom_track_25.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_102_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_22_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_19.mux_l1_in_1__S mux_bottom_track_19.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_203 vgnd vpwr scs8hd_decap_12
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_258 vgnd vpwr scs8hd_decap_12
XFILLER_25_236 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D mux_right_track_32.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_62 vgnd vpwr scs8hd_decap_3
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_23.scs8hd_buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X _116_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA__104__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_195 vpwr vgnd scs8hd_fill_2
XFILLER_3_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_34_ chanx_right_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.scs8hd_buf_4_0__A mux_left_track_3.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D mux_left_track_9.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_265 vgnd vpwr scs8hd_decap_8
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XFILLER_24_19 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_7.mux_l1_in_2_/S
+ mem_bottom_track_7.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_224 vgnd vpwr scs8hd_decap_4
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_29.mux_l2_in_0__A0 _065_/HI vgnd vpwr scs8hd_diode_2
XFILLER_4_7 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_1__A0 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_55 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XFILLER_17_172 vpwr vgnd scs8hd_fill_2
XFILLER_17_194 vpwr vgnd scs8hd_fill_2
XFILLER_15_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D mux_left_track_9.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_31 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 mux_left_track_9.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_31.scs8hd_buf_4_0_ mux_bottom_track_31.mux_l2_in_0_/X _112_/A vgnd
+ vpwr scs8hd_buf_1
Xmem_bottom_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S mem_bottom_track_25.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
X_101_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_41 vpwr vgnd scs8hd_fill_2
XFILLER_7_116 vgnd vpwr scs8hd_decap_4
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XFILLER_34_259 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.scs8hd_buf_4_0__A mux_bottom_track_13.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_43 vgnd vpwr scs8hd_fill_1
XFILLER_8_87 vpwr vgnd scs8hd_fill_2
XFILLER_6_193 vpwr vgnd scs8hd_fill_2
XFILLER_25_215 vgnd vpwr scs8hd_decap_12
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_27.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[15] mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.scs8hd_buf_4_0__A mux_right_track_2.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_39.scs8hd_buf_4_0__A mux_bottom_track_39.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_39.mux_l2_in_0_ _037_/HI mux_bottom_track_39.mux_l1_in_0_/X mux_bottom_track_39.mux_l2_in_0_/S
+ mux_bottom_track_39.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_207 vpwr vgnd scs8hd_fill_2
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_37.mux_l2_in_0__A0 _036_/HI vgnd vpwr scs8hd_diode_2
XFILLER_0_144 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_273 vpwr vgnd scs8hd_fill_2
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__D mux_bottom_track_19.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_203 vpwr vgnd scs8hd_fill_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_39.mux_l1_in_0__S mux_bottom_track_39.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_29.mux_l2_in_0__A1 mux_bottom_track_29.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_228 vpwr vgnd scs8hd_fill_2
XFILLER_2_206 vpwr vgnd scs8hd_fill_2
XFILLER_26_173 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XFILLER_25_74 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_1_ _046_/HI mux_left_track_5.mux_l1_in_2_/X mux_left_track_5.mux_l2_in_1_/S
+ mux_left_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XFILLER_14_143 vpwr vgnd scs8hd_fill_2
XFILLER_14_165 vpwr vgnd scs8hd_fill_2
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_102 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_100_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_11_146 vpwr vgnd scs8hd_fill_2
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_2__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_1_ chany_bottom_in[15] mux_left_track_5.mux_l1_in_2_/S
+ mux_left_track_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_8_66 vgnd vpwr scs8hd_decap_4
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_249 vpwr vgnd scs8hd_fill_2
XFILLER_25_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A mux_bottom_track_1.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__S mux_bottom_track_7.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_238 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vpwr vgnd scs8hd_fill_2
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_1__S mux_bottom_track_15.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.scs8hd_buf_4_0__A mux_right_track_24.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_219 vpwr vgnd scs8hd_fill_2
XFILLER_21_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_37.mux_l2_in_0__A1 mux_bottom_track_37.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D mux_right_track_16.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_234 vpwr vgnd scs8hd_fill_2
XFILLER_5_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_10 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_3
XFILLER_14_87 vgnd vpwr scs8hd_decap_3
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_39.mux_l1_in_0_ chanx_left_in[0] bottom_left_grid_pin_41_ mux_bottom_track_39.mux_l1_in_0_/S
+ mux_bottom_track_39.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__126__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_185 vgnd vpwr scs8hd_decap_12
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XFILLER_2_68 vpwr vgnd scs8hd_fill_2
XFILLER_1_273 vgnd vpwr scs8hd_decap_4
XFILLER_17_130 vgnd vpwr scs8hd_fill_1
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_133 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_25.mux_l2_in_1_ _043_/HI chany_bottom_in[18] mux_left_track_25.mux_l2_in_1_/S
+ mux_left_track_25.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__D mux_bottom_track_5.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_122 vgnd vpwr scs8hd_fill_1
XFILLER_14_199 vpwr vgnd scs8hd_fill_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_158 vgnd vpwr scs8hd_decap_4
XFILLER_20_114 vgnd vpwr scs8hd_decap_8
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_76 vpwr vgnd scs8hd_fill_2
XFILLER_7_129 vgnd vpwr scs8hd_decap_4
XFILLER_11_169 vgnd vpwr scs8hd_decap_4
XFILLER_0_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_19_214 vgnd vpwr scs8hd_decap_4
Xmux_left_track_5.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_left_track_5.mux_l1_in_2_/S
+ mux_left_track_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XFILLER_17_21 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_143 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_15_261 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.scs8hd_buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _126_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_179 vgnd vpwr scs8hd_fill_1
XFILLER_8_202 vpwr vgnd scs8hd_fill_2
XFILLER_12_242 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l2_in_0_/S mem_bottom_track_33.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_66 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_5_249 vgnd vpwr scs8hd_fill_1
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_197 vgnd vpwr scs8hd_decap_12
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_35.mux_l1_in_0__S mux_bottom_track_35.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_134 vpwr vgnd scs8hd_fill_2
XFILLER_23_101 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_1_/S mux_left_track_25.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_178 vgnd vpwr scs8hd_decap_4
XFILLER_2_7 vgnd vpwr scs8hd_decap_3
XFILLER_11_78 vpwr vgnd scs8hd_fill_2
XFILLER_14_101 vpwr vgnd scs8hd_fill_2
XFILLER_14_178 vpwr vgnd scs8hd_fill_2
XFILLER_37_248 vpwr vgnd scs8hd_fill_2
XFILLER_9_193 vgnd vpwr scs8hd_decap_4
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 mux_bottom_track_3.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l3_in_0_ mux_bottom_track_11.mux_l2_in_1_/X mux_bottom_track_11.mux_l2_in_0_/X
+ mux_bottom_track_11.mux_l3_in_0_/S mux_bottom_track_11.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_ chanx_right_in[14] chanx_right_in[5] mux_left_track_5.mux_l1_in_2_/S
+ mux_left_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_35 vpwr vgnd scs8hd_fill_2
XFILLER_8_46 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A mux_bottom_track_9.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_left_track_25.mux_l1_in_1_/S
+ mux_left_track_25.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_089_ chanx_left_in[17] chanx_right_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__D mux_bottom_track_25.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D mux_bottom_track_9.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_177 vgnd vpwr scs8hd_decap_4
XFILLER_3_111 vpwr vgnd scs8hd_fill_2
XFILLER_3_199 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A1 mux_bottom_track_11.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l2_in_1_ _056_/HI chanx_left_in[19] mux_bottom_track_11.mux_l2_in_1_/S
+ mux_bottom_track_11.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_232 vgnd vpwr scs8hd_fill_1
XFILLER_0_103 vgnd vpwr scs8hd_decap_3
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_265 vgnd vpwr scs8hd_decap_8
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_31.mux_l2_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/S mem_bottom_track_33.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D mux_right_track_0.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.scs8hd_buf_4_0__A mux_bottom_track_21.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_228 vgnd vpwr scs8hd_fill_1
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_56 vpwr vgnd scs8hd_fill_2
XFILLER_30_99 vgnd vpwr scs8hd_fill_1
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__S mux_bottom_track_27.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_121 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_25_22 vgnd vpwr scs8hd_decap_12
XFILLER_25_11 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_17_176 vpwr vgnd scs8hd_fill_2
XFILLER_17_187 vgnd vpwr scs8hd_decap_4
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_157 vpwr vgnd scs8hd_fill_2
XFILLER_11_35 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_135 vpwr vgnd scs8hd_fill_2
XFILLER_14_157 vpwr vgnd scs8hd_fill_2
XFILLER_28_7 vgnd vpwr scs8hd_decap_12
XFILLER_20_149 vpwr vgnd scs8hd_fill_2
XFILLER_9_161 vpwr vgnd scs8hd_fill_2
XFILLER_36_271 vgnd vpwr scs8hd_decap_4
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 mux_bottom_track_3.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_105 vpwr vgnd scs8hd_fill_2
XFILLER_22_45 vgnd vpwr scs8hd_decap_4
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_19_249 vgnd vpwr scs8hd_decap_4
Xmux_left_track_25.mux_l1_in_0_ chanx_right_in[18] chanx_right_in[9] mux_left_track_25.mux_l1_in_1_/S
+ mux_left_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_193 vpwr vgnd scs8hd_fill_2
X_088_ chanx_left_in[18] chanx_right_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_6_164 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_15.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l2_in_0_/S mem_bottom_track_15.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D mux_right_track_0.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_271 vgnd vpwr scs8hd_decap_4
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_56 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_22 vgnd vpwr scs8hd_decap_12
XFILLER_33_11 vgnd vpwr scs8hd_decap_4
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_7.mux_l1_in_3_ _039_/HI chanx_left_in[11] mux_bottom_track_7.mux_l1_in_2_/S
+ mux_bottom_track_7.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l2_in_0_ chanx_left_in[9] mux_bottom_track_11.mux_l1_in_0_/X
+ mux_bottom_track_11.mux_l2_in_1_/S mux_bottom_track_11.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
Xmux_bottom_track_29.scs8hd_buf_4_0_ mux_bottom_track_29.mux_l2_in_0_/X _113_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_21_222 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_99 vgnd vpwr scs8hd_fill_1
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l3_in_0__S mux_left_track_17.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_148 vgnd vpwr scs8hd_fill_1
XFILLER_12_233 vgnd vpwr scs8hd_fill_1
XFILLER_5_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A0 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_10_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_207 vpwr vgnd scs8hd_fill_2
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D mux_left_track_17.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 right_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
XFILLER_26_133 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_34 vgnd vpwr scs8hd_decap_12
XPHY_45 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_7.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_32.scs8hd_buf_4_0__A mux_right_track_32.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_32_136 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.scs8hd_buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _079_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_17_133 vgnd vpwr scs8hd_decap_3
XFILLER_17_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l1_in_1_ _052_/HI chanx_left_in[10] mux_right_track_32.mux_l1_in_1_/S
+ mux_right_track_32.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vgnd vpwr scs8hd_fill_1
XFILLER_22_180 vgnd vpwr scs8hd_decap_4
XFILLER_14_147 vgnd vpwr scs8hd_decap_6
Xmem_left_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l3_in_0_/S
+ mem_left_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_128 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.mux_l2_in_1_ mux_bottom_track_7.mux_l1_in_3_/X mux_bottom_track_7.mux_l1_in_2_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_31.mux_l1_in_0__S mux_bottom_track_31.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__074__A chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_22_68 vgnd vpwr scs8hd_decap_6
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_087_ _087_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_172 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_15.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l1_in_1_/S mem_bottom_track_15.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_37.scs8hd_buf_4_0_ mux_bottom_track_37.mux_l2_in_0_/X _109_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XANTENNA__069__A chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_34 vgnd vpwr scs8hd_decap_12
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A0 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_2_ chanx_left_in[6] bottom_left_grid_pin_41_ mux_bottom_track_7.mux_l1_in_2_/S
+ mux_bottom_track_7.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_245 vpwr vgnd scs8hd_fill_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_29.scs8hd_buf_4_0__A mux_bottom_track_29.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A0 _038_/HI vgnd vpwr scs8hd_diode_2
XFILLER_8_238 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A1 chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A0 mux_bottom_track_7.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D mux_right_track_4.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_25.scs8hd_buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _075_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_29_142 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[9] mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_252 vgnd vpwr scs8hd_decap_4
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_23.mux_l2_in_0_ mux_bottom_track_23.mux_l1_in_1_/X mux_bottom_track_23.mux_l1_in_0_/X
+ mux_bottom_track_23.mux_l2_in_0_/S mux_bottom_track_23.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA__077__A chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_6
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_46 vgnd vpwr scs8hd_decap_12
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_32_148 vgnd vpwr scs8hd_decap_4
XFILLER_15_90 vgnd vpwr scs8hd_decap_4
XFILLER_23_126 vpwr vgnd scs8hd_fill_2
Xmux_right_track_32.mux_l1_in_0_ chany_bottom_in[13] chany_bottom_in[6] mux_right_track_32.mux_l1_in_1_/S
+ mux_right_track_32.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_23.mux_l2_in_0__S mux_bottom_track_23.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_22_192 vgnd vpwr scs8hd_decap_8
Xmem_left_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_1_/S
+ mem_left_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_130 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_23.mux_l1_in_1_ _062_/HI chanx_left_in[17] mux_bottom_track_23.mux_l1_in_1_/S
+ mux_bottom_track_23.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l3_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_0_7 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_31.mux_l1_in_0__A0 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA__090__A chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
X_086_ _086_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_111 vpwr vgnd scs8hd_fill_2
XFILLER_6_122 vgnd vpwr scs8hd_fill_1
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 _041_/HI vgnd vpwr scs8hd_diode_2
XFILLER_17_25 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_46 vgnd vpwr scs8hd_decap_12
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A1 chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_15_221 vpwr vgnd scs8hd_fill_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_1_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_7.mux_l1_in_2_/S mux_bottom_track_7.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_254 vgnd vpwr scs8hd_decap_4
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_069_ chanx_right_in[17] chanx_left_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
Xmux_left_track_33.scs8hd_buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _071_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_9_81 vpwr vgnd scs8hd_fill_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_8_206 vpwr vgnd scs8hd_fill_2
XFILLER_12_224 vgnd vpwr scs8hd_decap_3
Xmem_right_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_4.mux_l1_in_2_/S mux_right_track_4.mux_l2_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A1 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.scs8hd_buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _106_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A1 mux_bottom_track_7.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D mux_right_track_24.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_154 vgnd vpwr scs8hd_decap_12
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XFILLER_4_264 vgnd vpwr scs8hd_decap_8
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XFILLER_6_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_decap_3
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.scs8hd_buf_4_0__A mux_left_track_17.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_2__D mux_bottom_track_11.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA__088__A chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D mux_right_track_4.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_105 vpwr vgnd scs8hd_fill_2
Xmem_left_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_1.mux_l3_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ mem_left_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_23.mux_l1_in_0_ bottom_left_grid_pin_41_ chanx_right_in[17] mux_bottom_track_23.mux_l1_in_1_/S
+ mux_bottom_track_23.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_9.mux_l1_in_1__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_90 vpwr vgnd scs8hd_fill_2
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vpwr vgnd scs8hd_fill_2
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_35.mux_l2_in_0_ _035_/HI mux_bottom_track_35.mux_l1_in_0_/X mux_bottom_track_35.mux_l2_in_0_/S
+ mux_bottom_track_35.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_5.mux_l1_in_0_/S mux_bottom_track_5.mux_l2_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_bottom_track_11.scs8hd_buf_4_0_ mux_bottom_track_11.mux_l3_in_0_/X _122_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_31.mux_l1_in_0__A1 chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_263 vgnd vpwr scs8hd_decap_12
XFILLER_8_39 vgnd vpwr scs8hd_decap_4
X_085_ _085_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_189 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 _059_/HI vgnd vpwr scs8hd_diode_2
XFILLER_26_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 left_top_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_17_48 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_decap_3
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_266 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[6] mux_bottom_track_7.mux_l1_in_2_/S
+ mux_bottom_track_7.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
X_068_ chanx_right_in[18] chanx_left_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_3
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 mux_bottom_track_17.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_2_/S
+ mem_right_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.scs8hd_buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X _123_/A vgnd
+ vpwr scs8hd_buf_1
Xmux_right_track_16.scs8hd_buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _099_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l2_in_1_ _041_/HI left_top_grid_pin_1_ mux_left_track_1.mux_l2_in_1_/S
+ mux_left_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__D mux_bottom_track_13.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_23.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_23.mux_l1_in_1_/S
+ mux_bottom_track_23.mux_l2_in_0_/S mem_bottom_track_23.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_29_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vgnd vpwr scs8hd_fill_1
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D mux_bottom_track_33.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_125 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_2_19 vpwr vgnd scs8hd_fill_2
XFILLER_1_235 vgnd vpwr scs8hd_decap_3
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_191 vgnd vpwr scs8hd_decap_12
XFILLER_11_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.scs8hd_buf_4_0__A mux_left_track_1.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_139 vpwr vgnd scs8hd_fill_2
XFILLER_26_80 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_5.mux_l1_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D mux_left_track_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_109 vpwr vgnd scs8hd_fill_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_275 vpwr vgnd scs8hd_fill_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
XFILLER_6_102 vgnd vpwr scs8hd_decap_3
X_084_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_4
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 _040_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 _049_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__D mux_bottom_track_13.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0__S mux_bottom_track_13.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_127 vgnd vpwr scs8hd_fill_1
Xmux_right_track_24.scs8hd_buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _095_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_23_70 vpwr vgnd scs8hd_fill_2
X_067_ _067_/HI _067_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_35.mux_l1_in_0_ bottom_left_grid_pin_39_ chanx_right_in[1] mux_bottom_track_35.mux_l1_in_0_/S
+ mux_bottom_track_35.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__D mux_bottom_track_33.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_259 vpwr vgnd scs8hd_fill_2
XFILLER_21_226 vgnd vpwr scs8hd_decap_6
XFILLER_21_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A0 mux_bottom_track_9.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A0 mux_right_track_16.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_81 vgnd vpwr scs8hd_decap_8
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ _119_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S mux_left_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_23.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l1_in_1_/S mem_bottom_track_23.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_29_178 vgnd vpwr scs8hd_decap_4
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_11.scs8hd_buf_4_0__A mux_bottom_track_11.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_6_84 vgnd vpwr scs8hd_decap_4
XPHY_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D mux_left_track_1.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vpwr vgnd scs8hd_fill_2
XFILLER_1_203 vgnd vpwr scs8hd_decap_3
XFILLER_32_129 vgnd vpwr scs8hd_decap_4
XFILLER_17_126 vgnd vpwr scs8hd_decap_4
XFILLER_17_159 vpwr vgnd scs8hd_fill_2
XFILLER_25_181 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_15_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.scs8hd_buf_4_0__A mux_right_track_0.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_118 vgnd vpwr scs8hd_decap_4
XFILLER_16_181 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_37.scs8hd_buf_4_0__A mux_bottom_track_37.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_1_ _050_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l3_in_0__S mux_bottom_track_9.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_118 vgnd vpwr scs8hd_decap_4
XFILLER_22_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l3_in_0__S mux_bottom_track_11.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_140 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A0 _034_/HI vgnd vpwr scs8hd_diode_2
XFILLER_9_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 _051_/HI vgnd vpwr scs8hd_diode_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_32.scs8hd_buf_4_0_ mux_right_track_32.mux_l2_in_0_/X _091_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
X_083_ _083_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_125 vgnd vpwr scs8hd_fill_1
XFILLER_6_158 vgnd vpwr scs8hd_decap_4
XFILLER_10_132 vpwr vgnd scs8hd_fill_2
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
XFILLER_10_176 vpwr vgnd scs8hd_fill_2
XFILLER_12_83 vpwr vgnd scs8hd_fill_2
XFILLER_18_210 vgnd vpwr scs8hd_decap_4
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1__S mux_right_track_8.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_23_93 vpwr vgnd scs8hd_fill_2
XFILLER_23_60 vgnd vpwr scs8hd_fill_1
X_066_ _066_/HI _066_/LO vgnd vpwr scs8hd_conb_1
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_21_249 vgnd vpwr scs8hd_decap_4
XFILLER_12_238 vpwr vgnd scs8hd_fill_2
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A1 mux_bottom_track_9.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A1 mux_right_track_16.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_220 vgnd vpwr scs8hd_decap_4
X_118_ _118_/A chany_bottom_out[9] vgnd vpwr scs8hd_buf_2
X_049_ _049_/HI _049_/LO vgnd vpwr scs8hd_conb_1
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_83 vgnd vpwr scs8hd_decap_8
XFILLER_20_61 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XFILLER_6_30 vgnd vpwr scs8hd_fill_1
XFILLER_6_41 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D mux_left_track_25.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_9_7 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[2] mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_9.scs8hd_buf_4_0__A mux_left_track_9.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_193 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
Xmux_left_track_33.mux_l2_in_1_ _045_/HI chany_bottom_in[19] mux_left_track_33.mux_l2_in_1_/S
+ mux_left_track_33.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_6
XFILLER_9_112 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A1 mux_bottom_track_33.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_178 vgnd vpwr scs8hd_decap_3
XFILLER_3_53 vgnd vpwr scs8hd_decap_4
XFILLER_3_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D mux_left_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_082_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_12_51 vpwr vgnd scs8hd_fill_2
XFILLER_12_62 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_1_ chanx_left_in[4] chany_bottom_in[18] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_222 vpwr vgnd scs8hd_fill_2
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_247 vgnd vpwr scs8hd_decap_8
XFILLER_24_236 vgnd vpwr scs8hd_decap_8
XFILLER_3_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__D mux_bottom_track_19.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.scs8hd_buf_4_0__A mux_left_track_25.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_15_258 vgnd vpwr scs8hd_fill_1
X_065_ _065_/HI _065_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_7 vgnd vpwr scs8hd_decap_8
XFILLER_0_21 vgnd vpwr scs8hd_decap_4
XFILLER_0_32 vgnd vpwr scs8hd_decap_3
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_76 vgnd vpwr scs8hd_decap_3
XFILLER_9_30 vpwr vgnd scs8hd_fill_2
XFILLER_9_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__D mux_bottom_track_39.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_29.mux_l1_in_0__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_21.mux_l1_in_1__S mux_bottom_track_21.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__S mux_bottom_track_7.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_11_261 vpwr vgnd scs8hd_fill_2
X_117_ _117_/A chany_bottom_out[10] vgnd vpwr scs8hd_buf_2
X_048_ _048_/HI _048_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_37.mux_l2_in_0__S mux_bottom_track_37.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_19.scs8hd_buf_4_0__A mux_bottom_track_19.mux_l2_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_64 vgnd vpwr scs8hd_decap_4
XFILLER_25_18 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.scs8hd_buf_4_0__A mux_right_track_8.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA__102__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_260 vpwr vgnd scs8hd_fill_2
XFILLER_31_153 vgnd vpwr scs8hd_decap_12
XFILLER_31_131 vgnd vpwr scs8hd_fill_1
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
Xmux_left_track_33.mux_l2_in_0_ chany_bottom_in[12] mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S mux_left_track_33.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_186 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_31.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_31.mux_l1_in_0_/S
+ mux_bottom_track_31.mux_l2_in_0_/S mem_bottom_track_31.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_9_102 vpwr vgnd scs8hd_fill_2
XFILLER_9_157 vpwr vgnd scs8hd_fill_2
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 _042_/HI vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_3_ _066_/HI chanx_left_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_19 vpwr vgnd scs8hd_fill_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_3__S mux_bottom_track_7.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_081_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_189 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_0_ chany_bottom_in[11] chany_bottom_in[4] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_37.mux_l1_in_0__A0 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_5_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_18 vpwr vgnd scs8hd_fill_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l3_in_0__A0 mux_left_track_17.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_204 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vpwr vgnd scs8hd_fill_2
XFILLER_23_51 vgnd vpwr scs8hd_decap_3
X_064_ _064_/HI _064_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_218 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_29.mux_l1_in_0__A1 chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_229 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D mux_left_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_62 vgnd vpwr scs8hd_decap_4
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _116_/A chany_bottom_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XFILLER_11_273 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
X_047_ _047_/HI _047_/LO vgnd vpwr scs8hd_conb_1
XFILLER_30_19 vgnd vpwr scs8hd_decap_12
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.scs8hd_buf_4_0_ mux_right_track_8.mux_l3_in_0_/X _103_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_20_96 vgnd vpwr scs8hd_decap_6
XFILLER_4_225 vpwr vgnd scs8hd_fill_2
XFILLER_4_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.scs8hd_buf_4_0__A mux_bottom_track_7.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D mux_left_track_17.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D mux_right_track_32.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_129 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_17_118 vgnd vpwr scs8hd_decap_4
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_173 vgnd vpwr scs8hd_decap_8
XFILLER_15_52 vpwr vgnd scs8hd_fill_2
XFILLER_15_96 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_25.mux_l2_in_1__A0 _043_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XFILLER_16_140 vpwr vgnd scs8hd_fill_2
XFILLER_16_173 vgnd vpwr scs8hd_decap_8
XFILLER_31_165 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_3.scs8hd_buf_4_0_ mux_left_track_3.mux_l3_in_0_/X _086_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_6 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_31.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_29.mux_l2_in_0_/S
+ mux_bottom_track_31.mux_l1_in_0_/S mem_bottom_track_31.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_13_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A1 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l1_in_2_ chanx_left_in[3] bottom_left_grid_pin_41_ mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A0 mux_left_track_25.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D mux_bottom_track_1.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_75 vpwr vgnd scs8hd_fill_2
XFILLER_12_97 vgnd vpwr scs8hd_fill_1
Xmux_left_track_33.mux_l1_in_0_ chany_bottom_in[5] chanx_right_in[10] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_17.scs8hd_buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X _119_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_37.mux_l1_in_0__A1 chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A1 mux_left_track_17.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_063_ _063_/HI _063_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S mux_bottom_track_17.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_2_197 vpwr vgnd scs8hd_fill_2
XFILLER_2_175 vpwr vgnd scs8hd_fill_2
XFILLER_2_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_8 vpwr vgnd scs8hd_fill_2
XFILLER_21_208 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_9_98 vpwr vgnd scs8hd_fill_2
XFILLER_28_19 vgnd vpwr scs8hd_decap_12
XFILLER_20_230 vgnd vpwr scs8hd_decap_3
XFILLER_18_41 vpwr vgnd scs8hd_fill_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_3
X_115_ _115_/A chany_bottom_out[12] vgnd vpwr scs8hd_buf_2
X_046_ _046_/HI _046_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_33.mux_l2_in_1__A0 _045_/HI vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_ _059_/HI chanx_left_in[13] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_215 vgnd vpwr scs8hd_fill_1
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_20_53 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_13.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l2_in_0_/S mem_bottom_track_13.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_6_11 vpwr vgnd scs8hd_fill_2
XFILLER_6_22 vpwr vgnd scs8hd_fill_2
XFILLER_6_88 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__D mux_bottom_track_21.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S mux_bottom_track_33.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 _050_/HI vgnd vpwr scs8hd_diode_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_25.mux_l2_in_1__A1 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_31_41 vgnd vpwr scs8hd_decap_12
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XFILLER_31_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_33.mux_l3_in_0__A0 mux_left_track_33.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_27.mux_l1_in_0__S mux_bottom_track_27.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
.ends

