* NGSPICE file created from sb_0__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_0__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_out[0]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_11_
+ top_left_grid_pin_13_ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_
+ top_left_grid_pin_5_ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_
+ vpwr vgnd
XFILLER_39_222 vpwr vgnd scs8hd_fill_2
Xmem_right_track_12.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_104 vgnd vpwr scs8hd_decap_8
XFILLER_36_258 vgnd vpwr scs8hd_decap_12
XFILLER_36_247 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_181 vgnd vpwr scs8hd_fill_1
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_27_258 vgnd vpwr scs8hd_decap_8
XFILLER_27_214 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _202_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_225 vgnd vpwr scs8hd_decap_6
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_24_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_217 vpwr vgnd scs8hd_fill_2
XFILLER_23_261 vgnd vpwr scs8hd_decap_4
X_131_ _129_/X _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_53 vgnd vpwr scs8hd_decap_8
XFILLER_23_86 vgnd vpwr scs8hd_decap_12
XANTENNA__110__C _126_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vgnd vpwr scs8hd_decap_12
XFILLER_14_250 vgnd vpwr scs8hd_decap_3
XANTENNA__119__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_30 vgnd vpwr scs8hd_fill_1
X_114_ _160_/B _130_/B vgnd vpwr scs8hd_buf_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _206_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_8
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _172_/Y mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_172 vpwr vgnd scs8hd_fill_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XANTENNA__116__B _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_40_189 vpwr vgnd scs8hd_fill_2
XFILLER_15_43 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vgnd vpwr scs8hd_decap_4
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_0_274 vgnd vpwr scs8hd_decap_3
XFILLER_31_123 vgnd vpwr scs8hd_decap_4
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_178 vpwr vgnd scs8hd_fill_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vpwr vgnd scs8hd_fill_2
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
Xmem_top_track_4.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_145 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_138 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_193 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_33_218 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vgnd vpwr scs8hd_fill_1
XFILLER_41_240 vgnd vpwr scs8hd_decap_4
XFILLER_5_174 vgnd vpwr scs8hd_decap_3
XFILLER_5_130 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
X_130_ _130_/A _130_/B _130_/C _168_/A _131_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_240 vgnd vpwr scs8hd_decap_4
XFILLER_23_98 vgnd vpwr scs8hd_decap_12
XANTENNA__110__D _171_/A vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_34 vgnd vpwr scs8hd_decap_12
XFILLER_9_89 vgnd vpwr scs8hd_decap_12
XANTENNA__135__A _129_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_243 vgnd vpwr scs8hd_decap_8
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XFILLER_7_225 vpwr vgnd scs8hd_fill_2
XFILLER_11_210 vpwr vgnd scs8hd_fill_2
X_113_ address[2] _160_/B vgnd vpwr scs8hd_inv_8
XFILLER_38_129 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_7 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.tap_buf4_0_.scs8hd_inv_1 mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_8
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_28_195 vgnd vpwr scs8hd_decap_4
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_55 vgnd vpwr scs8hd_decap_6
XFILLER_25_110 vgnd vpwr scs8hd_decap_8
XFILLER_25_154 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_235 vgnd vpwr scs8hd_decap_8
XFILLER_22_168 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_117 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_190 vpwr vgnd scs8hd_fill_2
XFILLER_27_227 vgnd vpwr scs8hd_decap_4
XFILLER_10_138 vpwr vgnd scs8hd_fill_2
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_41_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_197 vgnd vpwr scs8hd_decap_12
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_274 vgnd vpwr scs8hd_fill_1
XFILLER_17_260 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_134 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XFILLER_9_46 vgnd vpwr scs8hd_decap_12
XFILLER_9_79 vgnd vpwr scs8hd_fill_1
XANTENNA__135__B _136_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_204 vgnd vpwr scs8hd_decap_12
XFILLER_7_259 vpwr vgnd scs8hd_fill_2
X_112_ _128_/A _110_/X _112_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_4.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _192_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_29_98 vgnd vpwr scs8hd_decap_12
XFILLER_28_141 vgnd vpwr scs8hd_decap_8
XFILLER_34_133 vgnd vpwr scs8hd_fill_1
XFILLER_19_130 vgnd vpwr scs8hd_decap_3
XFILLER_19_152 vpwr vgnd scs8hd_fill_2
XFILLER_34_188 vgnd vpwr scs8hd_fill_1
XFILLER_40_158 vgnd vpwr scs8hd_decap_12
XFILLER_40_125 vgnd vpwr scs8hd_decap_3
XFILLER_25_177 vgnd vpwr scs8hd_decap_4
XFILLER_16_144 vgnd vpwr scs8hd_decap_3
XFILLER_16_166 vpwr vgnd scs8hd_fill_2
XFILLER_31_169 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _126_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_136 vgnd vpwr scs8hd_decap_3
XFILLER_13_158 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _196_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_206 vgnd vpwr scs8hd_decap_8
XFILLER_36_228 vgnd vpwr scs8hd_decap_4
XANTENNA__138__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_162 vgnd vpwr scs8hd_fill_1
XFILLER_12_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_275 vpwr vgnd scs8hd_fill_2
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__C _153_/C vgnd vpwr scs8hd_diode_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_32_242 vgnd vpwr scs8hd_decap_4
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_45 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_157 vgnd vpwr scs8hd_decap_12
XFILLER_2_146 vgnd vpwr scs8hd_decap_3
XFILLER_9_58 vgnd vpwr scs8hd_decap_3
XFILLER_14_242 vpwr vgnd scs8hd_fill_2
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _200_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_216 vgnd vpwr scs8hd_decap_6
X_111_ _096_/X _110_/X _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_234 vpwr vgnd scs8hd_fill_2
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XFILLER_11_256 vpwr vgnd scs8hd_fill_2
XFILLER_11_267 vpwr vgnd scs8hd_fill_2
XANTENNA__146__B _130_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_260 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_208 vgnd vpwr scs8hd_decap_6
XFILLER_29_33 vgnd vpwr scs8hd_decap_12
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_186 vgnd vpwr scs8hd_decap_6
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_145 vgnd vpwr scs8hd_decap_8
XANTENNA__157__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XFILLER_19_197 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _204_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XFILLER_25_167 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_31_148 vpwr vgnd scs8hd_fill_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _153_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_226 vgnd vpwr scs8hd_fill_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_115 vgnd vpwr scs8hd_decap_6
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_130 vgnd vpwr scs8hd_decap_6
XFILLER_8_174 vgnd vpwr scs8hd_decap_4
XANTENNA__154__B _154_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_251 vgnd vpwr scs8hd_decap_4
XFILLER_26_262 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vpwr vgnd scs8hd_fill_2
XFILLER_5_166 vpwr vgnd scs8hd_fill_2
XANTENNA__140__D _160_/D vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_221 vpwr vgnd scs8hd_fill_2
XANTENNA__165__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_221 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_169 vgnd vpwr scs8hd_decap_12
XFILLER_14_210 vpwr vgnd scs8hd_fill_2
XFILLER_14_232 vgnd vpwr scs8hd_fill_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_180 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_213 vgnd vpwr scs8hd_fill_1
XFILLER_20_224 vpwr vgnd scs8hd_fill_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _115_/A _126_/B _126_/C _171_/A _110_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd
+ vpwr scs8hd_diode_2
X_239_ _239_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _153_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_250 vgnd vpwr scs8hd_fill_1
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
XFILLER_37_154 vgnd vpwr scs8hd_decap_3
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_37_198 vgnd vpwr scs8hd_decap_3
XFILLER_37_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_45 vgnd vpwr scs8hd_decap_12
XFILLER_29_23 vgnd vpwr scs8hd_decap_3
XFILLER_28_154 vgnd vpwr scs8hd_decap_6
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_264 vgnd vpwr scs8hd_decap_12
XFILLER_3_231 vgnd vpwr scs8hd_decap_8
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XFILLER_34_113 vgnd vpwr scs8hd_decap_3
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_113 vgnd vpwr scs8hd_decap_3
XFILLER_16_157 vpwr vgnd scs8hd_fill_2
XFILLER_16_179 vpwr vgnd scs8hd_fill_2
XANTENNA__143__D _149_/D vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_249 vgnd vpwr scs8hd_decap_4
XANTENNA__168__A _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_105 vgnd vpwr scs8hd_fill_1
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__170__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_263 vgnd vpwr scs8hd_decap_12
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_274 vgnd vpwr scs8hd_fill_1
Xmem_right_track_0.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_134 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_4
Xmem_top_track_8.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__C _153_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_274 vgnd vpwr scs8hd_decap_3
XFILLER_32_266 vgnd vpwr scs8hd_decap_8
XFILLER_32_255 vgnd vpwr scs8hd_decap_8
XANTENNA__165__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_200 vgnd vpwr scs8hd_decap_8
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_270 vgnd vpwr scs8hd_decap_6
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_7_229 vpwr vgnd scs8hd_fill_2
XFILLER_11_214 vgnd vpwr scs8hd_decap_3
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_238_ _238_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
X_169_ _168_/A _168_/B _162_/A _169_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__146__D _160_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_57 vgnd vpwr scs8hd_decap_4
XFILLER_3_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__157__C _153_/C vgnd vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_8
XFILLER_25_136 vpwr vgnd scs8hd_fill_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _190_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_150 vgnd vpwr scs8hd_fill_1
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_14.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_161 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_172 vpwr vgnd scs8hd_fill_2
XFILLER_12_194 vpwr vgnd scs8hd_fill_2
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_8
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XANTENNA__149__D _149_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _194_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vgnd vpwr scs8hd_decap_3
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_14_256 vgnd vpwr scs8hd_decap_8
XFILLER_14_267 vgnd vpwr scs8hd_decap_8
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
X_237_ _237_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_168_ _168_/A _168_/B _161_/A _168_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
X_099_ address[4] address[5] _130_/C vgnd vpwr scs8hd_or2_4
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_3
XFILLER_1_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_8
XFILLER_19_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__157__D _149_/D vgnd vpwr scs8hd_diode_2
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_218 vpwr vgnd scs8hd_fill_2
XANTENNA__168__C _161_/A vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_173 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _202_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_195 vpwr vgnd scs8hd_fill_2
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_151 vpwr vgnd scs8hd_fill_2
XFILLER_35_243 vgnd vpwr scs8hd_fill_1
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_213 vgnd vpwr scs8hd_decap_12
XFILLER_41_202 vpwr vgnd scs8hd_fill_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_232 vgnd vpwr scs8hd_fill_1
XFILLER_23_213 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XFILLER_23_49 vpwr vgnd scs8hd_fill_2
XFILLER_23_257 vpwr vgnd scs8hd_fill_2
XFILLER_23_268 vgnd vpwr scs8hd_decap_8
XFILLER_2_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
XFILLER_14_246 vpwr vgnd scs8hd_fill_2
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_4.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_238 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_236_ _236_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_167_ _166_/X _168_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_242 vgnd vpwr scs8hd_decap_8
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
X_098_ address[2] _126_/B vgnd vpwr scs8hd_buf_1
XFILLER_37_135 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_8
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_8
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_160 vpwr vgnd scs8hd_fill_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_105 vgnd vpwr scs8hd_decap_8
XFILLER_16_127 vgnd vpwr scs8hd_decap_6
XFILLER_16_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_193 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
XFILLER_30_185 vgnd vpwr scs8hd_decap_6
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_263 vgnd vpwr scs8hd_decap_12
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_145 vgnd vpwr scs8hd_decap_8
XFILLER_8_178 vgnd vpwr scs8hd_fill_1
XFILLER_12_163 vgnd vpwr scs8hd_decap_3
XFILLER_35_222 vpwr vgnd scs8hd_fill_2
XFILLER_35_211 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_41_236 vpwr vgnd scs8hd_fill_2
XFILLER_41_225 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_26_211 vgnd vpwr scs8hd_fill_1
Xmem_top_track_10.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_225 vgnd vpwr scs8hd_decap_4
XFILLER_17_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XFILLER_23_39 vgnd vpwr scs8hd_decap_6
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_151 vgnd vpwr scs8hd_decap_3
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_235_ _235_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ address[3] _115_/A vgnd vpwr scs8hd_buf_1
X_166_ address[3] address[2] address[4] _138_/B _166_/X vgnd vpwr scs8hd_or4_4
XFILLER_34_6 vgnd vpwr scs8hd_decap_12
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_191 vgnd vpwr scs8hd_decap_4
XFILLER_10_84 vgnd vpwr scs8hd_decap_8
XFILLER_19_114 vgnd vpwr scs8hd_decap_4
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ address[3] _130_/B _153_/C _149_/D _150_/B vgnd vpwr scs8hd_or4_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_275 vpwr vgnd scs8hd_fill_2
XFILLER_29_231 vgnd vpwr scs8hd_fill_1
XFILLER_12_131 vgnd vpwr scs8hd_decap_8
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_201 vpwr vgnd scs8hd_fill_2
XFILLER_41_259 vpwr vgnd scs8hd_fill_2
XFILLER_26_245 vgnd vpwr scs8hd_decap_4
XFILLER_5_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_4
XFILLER_32_215 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _130_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_241 vgnd vpwr scs8hd_fill_1
XFILLER_20_207 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _192_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
X_234_ _234_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_165_ _162_/A _164_/B _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _152_/A _096_/X vgnd vpwr scs8hd_buf_1
XFILLER_37_159 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_126 vpwr vgnd scs8hd_fill_2
XFILLER_19_148 vpwr vgnd scs8hd_fill_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_4
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
X_148_ _151_/A _148_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_15_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_181 vpwr vgnd scs8hd_fill_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_33_195 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vpwr vgnd scs8hd_fill_2
XFILLER_33_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vgnd vpwr scs8hd_decap_8
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XFILLER_30_154 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_38_243 vgnd vpwr scs8hd_fill_1
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_210 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_176 vpwr vgnd scs8hd_fill_2
XFILLER_8_158 vpwr vgnd scs8hd_fill_2
XFILLER_12_198 vgnd vpwr scs8hd_decap_3
XANTENNA__103__A _160_/D vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_238 vpwr vgnd scs8hd_fill_2
XFILLER_17_224 vgnd vpwr scs8hd_decap_8
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _200_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
Xmem_right_track_14.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_18 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_164_ _161_/A _164_/B _164_/Y vgnd vpwr scs8hd_nor2_4
X_233_ _233_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_095_ address[0] _152_/A vgnd vpwr scs8hd_inv_8
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_29 vpwr vgnd scs8hd_fill_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XFILLER_28_149 vpwr vgnd scs8hd_fill_2
XFILLER_34_119 vgnd vpwr scs8hd_decap_8
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
X_147_ _129_/X _148_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_270 vgnd vpwr scs8hd_decap_4
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_171 vgnd vpwr scs8hd_decap_3
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _188_/A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_144 vgnd vpwr scs8hd_decap_6
XFILLER_30_133 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_199 vpwr vgnd scs8hd_fill_2
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XFILLER_8_126 vpwr vgnd scs8hd_fill_2
XFILLER_41_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_40 vgnd vpwr scs8hd_decap_12
XFILLER_17_236 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _160_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_228 vpwr vgnd scs8hd_fill_2
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_110 vgnd vpwr scs8hd_decap_4
XFILLER_1_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _149_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_276 vgnd vpwr scs8hd_fill_1
X_232_ _232_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_163_ _121_/Y _160_/B _160_/C _149_/D _164_/B vgnd vpwr scs8hd_or4_4
XANTENNA__111__B _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_139 vgnd vpwr scs8hd_decap_4
XFILLER_37_128 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_76 vgnd vpwr scs8hd_fill_1
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_194 vgnd vpwr scs8hd_decap_3
XFILLER_27_161 vpwr vgnd scs8hd_fill_2
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_19_106 vgnd vpwr scs8hd_decap_3
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
X_146_ address[3] _130_/B _153_/C _160_/D _148_/B vgnd vpwr scs8hd_or4_4
XANTENNA__122__A _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_175 vpwr vgnd scs8hd_fill_2
XFILLER_18_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_197 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_86 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_164 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
X_129_ _152_/A _129_/X vgnd vpwr scs8hd_buf_1
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
XFILLER_29_234 vpwr vgnd scs8hd_fill_2
XFILLER_29_201 vgnd vpwr scs8hd_decap_4
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_145 vgnd vpwr scs8hd_decap_4
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_52 vgnd vpwr scs8hd_decap_8
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_25_270 vgnd vpwr scs8hd_decap_6
XFILLER_4_196 vgnd vpwr scs8hd_decap_12
XFILLER_4_185 vpwr vgnd scs8hd_fill_2
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_240 vpwr vgnd scs8hd_fill_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_22_262 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_233 vgnd vpwr scs8hd_decap_8
XFILLER_9_255 vpwr vgnd scs8hd_fill_2
XFILLER_9_266 vpwr vgnd scs8hd_fill_2
XFILLER_13_273 vgnd vpwr scs8hd_decap_4
Xmem_top_track_14.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__A _128_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
X_231_ _231_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_162_ _162_/A _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_221 vgnd vpwr scs8hd_decap_4
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmem_right_track_10.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_195 vgnd vpwr scs8hd_fill_1
XFILLER_3_239 vgnd vpwr scs8hd_decap_3
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_118 vgnd vpwr scs8hd_fill_1
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_8
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _190_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _151_/A _145_/B _145_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_6
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_132 vpwr vgnd scs8hd_fill_2
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_165 vpwr vgnd scs8hd_fill_2
XFILLER_24_176 vgnd vpwr scs8hd_decap_6
XFILLER_21_98 vgnd vpwr scs8hd_decap_8
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _151_/A vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_235 vgnd vpwr scs8hd_decap_8
XFILLER_38_224 vgnd vpwr scs8hd_decap_3
XFILLER_38_213 vgnd vpwr scs8hd_fill_1
Xmux_top_track_10.tap_buf4_0_.scs8hd_inv_1 mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_168 vpwr vgnd scs8hd_fill_2
XFILLER_20_190 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_205 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_205 vgnd vpwr scs8hd_decap_4
XFILLER_4_175 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA__130__B _130_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_230 vgnd vpwr scs8hd_fill_1
XFILLER_22_252 vgnd vpwr scs8hd_fill_1
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_3
XFILLER_1_156 vgnd vpwr scs8hd_decap_12
Xmem_right_track_6.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_212 vpwr vgnd scs8hd_fill_2
XFILLER_9_245 vgnd vpwr scs8hd_fill_1
XFILLER_13_241 vgnd vpwr scs8hd_fill_1
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_193 vgnd vpwr scs8hd_decap_4
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
X_230_ _230_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_161_ _161_/A _162_/B _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_174 vgnd vpwr scs8hd_decap_8
XFILLER_3_207 vgnd vpwr scs8hd_decap_12
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_98 vgnd vpwr scs8hd_decap_8
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_174 vgnd vpwr scs8hd_decap_8
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _129_/X _145_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_33_199 vpwr vgnd scs8hd_fill_2
XFILLER_33_155 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_158 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
X_127_ _096_/X _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_247 vgnd vpwr scs8hd_decap_8
XFILLER_29_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_239 vpwr vgnd scs8hd_fill_2
XANTENNA__144__A _129_/X vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vgnd vpwr scs8hd_decap_8
XFILLER_26_228 vgnd vpwr scs8hd_decap_8
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _186_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_98 vgnd vpwr scs8hd_decap_12
XANTENNA__130__C _130_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_231 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_272 vgnd vpwr scs8hd_decap_3
XFILLER_1_135 vpwr vgnd scs8hd_fill_2
XFILLER_1_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__141__B _140_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_227 vgnd vpwr scs8hd_decap_4
XFILLER_10_245 vpwr vgnd scs8hd_fill_2
X_160_ _121_/Y _160_/B _160_/C _160_/D _162_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B _136_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _152_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_10.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_219 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_8
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
X_143_ _115_/A _126_/B _153_/C _149_/D _145_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
XFILLER_18_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__147__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_134 vpwr vgnd scs8hd_fill_2
X_126_ _130_/A _126_/B _126_/C _171_/A _127_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_37_270 vgnd vpwr scs8hd_decap_6
XFILLER_29_259 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_35_218 vpwr vgnd scs8hd_fill_2
XFILLER_35_207 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_270 vgnd vpwr scs8hd_decap_4
XANTENNA__144__B _145_/B vgnd vpwr scs8hd_diode_2
X_109_ _149_/D _171_/A vgnd vpwr scs8hd_buf_1
XANTENNA__160__A _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_40_243 vgnd vpwr scs8hd_fill_1
XANTENNA__130__D _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_276 vgnd vpwr scs8hd_fill_1
XFILLER_31_254 vpwr vgnd scs8hd_fill_2
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_114 vgnd vpwr scs8hd_fill_1
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_203 vgnd vpwr scs8hd_decap_6
XFILLER_9_225 vpwr vgnd scs8hd_fill_2
XFILLER_13_221 vpwr vgnd scs8hd_fill_2
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XFILLER_13_265 vpwr vgnd scs8hd_fill_2
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_39_151 vpwr vgnd scs8hd_fill_2
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_272 vgnd vpwr scs8hd_decap_4
XFILLER_5_261 vgnd vpwr scs8hd_decap_4
XFILLER_36_198 vpwr vgnd scs8hd_fill_2
Xmem_right_track_2.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_110 vgnd vpwr scs8hd_decap_8
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
X_142_ _151_/A _140_/X _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_253 vpwr vgnd scs8hd_fill_2
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
XANTENNA__147__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_198 vgnd vpwr scs8hd_decap_8
XFILLER_41_190 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _121_/Y vgnd vpwr scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_15_102 vgnd vpwr scs8hd_fill_1
XFILLER_15_168 vpwr vgnd scs8hd_fill_2
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_125_ _128_/A _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_38_205 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_138 vgnd vpwr scs8hd_decap_4
XFILLER_29_227 vgnd vpwr scs8hd_decap_4
XFILLER_29_238 vgnd vpwr scs8hd_decap_6
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_127 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
X_108_ address[1] enable _149_/D vgnd vpwr scs8hd_nand2_4
XFILLER_11_160 vpwr vgnd scs8hd_fill_2
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _160_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XFILLER_27_12 vpwr vgnd scs8hd_fill_2
XFILLER_40_211 vgnd vpwr scs8hd_decap_3
XFILLER_40_200 vgnd vpwr scs8hd_decap_8
XFILLER_4_189 vgnd vpwr scs8hd_decap_4
XFILLER_4_167 vgnd vpwr scs8hd_decap_8
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_16_230 vgnd vpwr scs8hd_decap_8
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_266 vpwr vgnd scs8hd_fill_2
XFILLER_31_200 vpwr vgnd scs8hd_fill_2
XANTENNA__171__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_233 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_259 vgnd vpwr scs8hd_decap_4
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_163 vpwr vgnd scs8hd_fill_2
XFILLER_39_130 vgnd vpwr scs8hd_fill_1
XFILLER_10_225 vgnd vpwr scs8hd_fill_1
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_27_133 vgnd vpwr scs8hd_decap_12
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _129_/X _140_/X _141_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _180_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_33_136 vpwr vgnd scs8hd_fill_2
XFILLER_18_177 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _160_/B vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_136 vgnd vpwr scs8hd_decap_6
XFILLER_24_169 vpwr vgnd scs8hd_fill_2
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
X_124_ _096_/X _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_91 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_6 vgnd vpwr scs8hd_decap_12
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_117 vgnd vpwr scs8hd_fill_1
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_139 vgnd vpwr scs8hd_fill_1
XFILLER_20_150 vgnd vpwr scs8hd_decap_3
XFILLER_20_161 vpwr vgnd scs8hd_fill_2
XFILLER_7_165 vgnd vpwr scs8hd_fill_1
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_110 vgnd vpwr scs8hd_decap_6
X_107_ _128_/A _104_/X _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__160__C _160_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__169__A _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_135 vgnd vpwr scs8hd_fill_1
XFILLER_16_253 vpwr vgnd scs8hd_fill_2
XFILLER_16_264 vgnd vpwr scs8hd_decap_8
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__171__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_22_245 vgnd vpwr scs8hd_decap_4
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _184_/A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vgnd vpwr scs8hd_decap_4
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_4
XFILLER_10_237 vgnd vpwr scs8hd_decap_8
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_241 vgnd vpwr scs8hd_fill_1
XFILLER_36_145 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_145 vgnd vpwr scs8hd_fill_1
XFILLER_27_123 vgnd vpwr scs8hd_fill_1
X_140_ _115_/A _126_/B _153_/C _160_/D _140_/X vgnd vpwr scs8hd_or4_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _188_/Y mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_167 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
Xmem_top_track_6.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_129 vpwr vgnd scs8hd_fill_2
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
X_123_ _130_/A _126_/B _126_/C _168_/A _124_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_229 vgnd vpwr scs8hd_decap_3
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__160__D _160_/D vgnd vpwr scs8hd_diode_2
X_106_ address[0] _128_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_80 vgnd vpwr scs8hd_decap_12
XANTENNA__169__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_262 vgnd vpwr scs8hd_decap_12
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_82 vgnd vpwr scs8hd_decap_8
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_221 vgnd vpwr scs8hd_fill_1
XFILLER_40_235 vgnd vpwr scs8hd_decap_8
XFILLER_40_224 vgnd vpwr scs8hd_decap_8
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_25_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__C _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_22_224 vgnd vpwr scs8hd_decap_6
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_117 vpwr vgnd scs8hd_fill_2
XFILLER_1_139 vgnd vpwr scs8hd_decap_12
XFILLER_13_202 vpwr vgnd scs8hd_fill_2
XFILLER_13_235 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_249 vgnd vpwr scs8hd_fill_1
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XFILLER_36_157 vgnd vpwr scs8hd_decap_6
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_113 vgnd vpwr scs8hd_decap_3
XFILLER_18_146 vgnd vpwr scs8hd_fill_1
XFILLER_41_171 vgnd vpwr scs8hd_fill_1
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__163__D _149_/D vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XFILLER_32_171 vgnd vpwr scs8hd_decap_4
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_138 vgnd vpwr scs8hd_decap_3
X_122_ _121_/Y _130_/A vgnd vpwr scs8hd_buf_1
XFILLER_21_108 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_10.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_274 vgnd vpwr scs8hd_fill_1
XFILLER_28_241 vgnd vpwr scs8hd_decap_8
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
X_105_ _096_/X _104_/X _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_200 vgnd vpwr scs8hd_decap_3
XANTENNA__169__C _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_274 vgnd vpwr scs8hd_decap_3
XFILLER_34_255 vgnd vpwr scs8hd_decap_8
XFILLER_34_211 vgnd vpwr scs8hd_fill_1
XFILLER_25_200 vpwr vgnd scs8hd_fill_2
XFILLER_25_255 vpwr vgnd scs8hd_fill_2
XFILLER_25_266 vpwr vgnd scs8hd_fill_2
XFILLER_40_247 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_258 vgnd vpwr scs8hd_decap_4
XFILLER_31_236 vpwr vgnd scs8hd_fill_2
XFILLER_31_225 vgnd vpwr scs8hd_decap_4
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_192 vgnd vpwr scs8hd_fill_1
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_225 vgnd vpwr scs8hd_decap_8
XFILLER_13_258 vgnd vpwr scs8hd_decap_4
XFILLER_9_229 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vpwr vgnd scs8hd_fill_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XANTENNA__166__D _138_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_5_51 vgnd vpwr scs8hd_decap_8
XFILLER_39_155 vpwr vgnd scs8hd_fill_2
XFILLER_39_199 vgnd vpwr scs8hd_decap_8
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_221 vgnd vpwr scs8hd_decap_8
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XFILLER_26_180 vgnd vpwr scs8hd_decap_6
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XFILLER_41_194 vgnd vpwr scs8hd_decap_4
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XFILLER_32_150 vgnd vpwr scs8hd_fill_1
XFILLER_24_117 vgnd vpwr scs8hd_decap_4
Xmem_right_track_6.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
X_121_ address[3] _121_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_194 vpwr vgnd scs8hd_fill_2
XFILLER_38_209 vgnd vpwr scs8hd_decap_4
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_172 vgnd vpwr scs8hd_decap_4
XFILLER_14_183 vpwr vgnd scs8hd_fill_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _178_/A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
Xmem_top_track_2.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_153 vgnd vpwr scs8hd_fill_1
XFILLER_11_164 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vpwr vgnd scs8hd_fill_2
X_104_ _115_/A _126_/B _126_/C _168_/A _104_/X vgnd vpwr scs8hd_or4_4
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_267 vgnd vpwr scs8hd_decap_8
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_16 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_fill_1
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_149 vgnd vpwr scs8hd_decap_4
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_204 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_182 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_167 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_4
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _182_/A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_233 vpwr vgnd scs8hd_fill_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_35_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vgnd vpwr scs8hd_decap_4
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_140 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_23_140 vgnd vpwr scs8hd_fill_1
X_120_ _128_/A _118_/X _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_162 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_fill_1
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _186_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_254 vpwr vgnd scs8hd_fill_2
XFILLER_16_18 vgnd vpwr scs8hd_decap_12
XFILLER_20_132 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vgnd vpwr scs8hd_decap_4
XFILLER_20_165 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
X_103_ _160_/D _168_/A vgnd vpwr scs8hd_buf_1
XFILLER_19_221 vpwr vgnd scs8hd_fill_2
XFILLER_19_254 vpwr vgnd scs8hd_fill_2
XFILLER_6_180 vgnd vpwr scs8hd_fill_1
XFILLER_27_28 vgnd vpwr scs8hd_decap_12
XFILLER_25_213 vpwr vgnd scs8hd_fill_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_249 vgnd vpwr scs8hd_fill_1
XFILLER_30_271 vgnd vpwr scs8hd_decap_4
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_9_209 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_242 vgnd vpwr scs8hd_decap_4
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vpwr vgnd scs8hd_fill_2
XFILLER_39_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_245 vgnd vpwr scs8hd_decap_3
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_4_6 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_105 vgnd vpwr scs8hd_decap_8
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_17_160 vpwr vgnd scs8hd_fill_2
XFILLER_32_185 vpwr vgnd scs8hd_fill_2
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_6
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_163 vgnd vpwr scs8hd_decap_3
XFILLER_14_196 vpwr vgnd scs8hd_fill_2
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_266 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
X_102_ address[1] _101_/Y _160_/D vgnd vpwr scs8hd_or2_4
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_225 vpwr vgnd scs8hd_fill_2
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_4_129 vgnd vpwr scs8hd_decap_6
XFILLER_16_247 vgnd vpwr scs8hd_decap_4
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_50 vgnd vpwr scs8hd_decap_8
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_195 vgnd vpwr scs8hd_decap_12
XFILLER_3_184 vgnd vpwr scs8hd_decap_8
XFILLER_3_162 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_8
XFILLER_13_206 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_40_18 vgnd vpwr scs8hd_decap_12
XFILLER_5_268 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vpwr vgnd scs8hd_fill_2
XFILLER_36_139 vgnd vpwr scs8hd_decap_3
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XFILLER_2_205 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_175 vgnd vpwr scs8hd_decap_8
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XPHY_51 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_175 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_14_120 vgnd vpwr scs8hd_decap_3
Xmux_top_track_4.tap_buf4_0_.scs8hd_inv_1 mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XANTENNA__107__A _128_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_234 vgnd vpwr scs8hd_decap_4
XFILLER_37_212 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_145 vgnd vpwr scs8hd_decap_3
XFILLER_20_178 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_201 vpwr vgnd scs8hd_fill_2
XFILLER_7_127 vgnd vpwr scs8hd_decap_3
XFILLER_7_116 vgnd vpwr scs8hd_fill_1
X_101_ enable _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_156 vgnd vpwr scs8hd_fill_1
XFILLER_19_201 vgnd vpwr scs8hd_decap_4
XFILLER_34_215 vgnd vpwr scs8hd_decap_3
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _176_/A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vpwr vgnd scs8hd_fill_2
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
XANTENNA__104__B _126_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _128_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_12_273 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _180_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_50 vgnd vpwr scs8hd_decap_8
XFILLER_36_129 vgnd vpwr scs8hd_decap_8
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vpwr vgnd scs8hd_fill_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vpwr vgnd scs8hd_fill_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_198 vgnd vpwr scs8hd_fill_1
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XANTENNA__112__B _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_140 vgnd vpwr scs8hd_fill_1
XFILLER_17_173 vgnd vpwr scs8hd_decap_4
XFILLER_23_110 vgnd vpwr scs8hd_decap_6
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XFILLER_23_143 vpwr vgnd scs8hd_fill_2
XFILLER_23_198 vgnd vpwr scs8hd_decap_4
XANTENNA__107__B _104_/X vgnd vpwr scs8hd_diode_2
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__123__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_224 vgnd vpwr scs8hd_decap_8
X_100_ _130_/C _126_/C vgnd vpwr scs8hd_buf_1
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XFILLER_34_205 vgnd vpwr scs8hd_decap_6
XFILLER_42_271 vgnd vpwr scs8hd_decap_6
XFILLER_34_238 vgnd vpwr scs8hd_decap_8
XFILLER_34_227 vgnd vpwr scs8hd_decap_8
XANTENNA__118__A _115_/A vgnd vpwr scs8hd_diode_2
X_229_ _229_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_172 vgnd vpwr scs8hd_decap_8
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_208 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _184_/Y mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_12.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_4
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_142 vgnd vpwr scs8hd_decap_4
XANTENNA__104__C _126_/C vgnd vpwr scs8hd_diode_2
Xmem_top_track_6.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_252 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_263 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_134 vgnd vpwr scs8hd_decap_8
XFILLER_0_145 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XANTENNA__115__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_127 vgnd vpwr scs8hd_fill_1
XANTENNA__131__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_182 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_237 vgnd vpwr scs8hd_decap_4
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
Xmux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_163 vpwr vgnd scs8hd_fill_2
XFILLER_35_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_163 vpwr vgnd scs8hd_fill_2
XFILLER_26_152 vgnd vpwr scs8hd_fill_1
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_86 vgnd vpwr scs8hd_decap_12
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_258 vgnd vpwr scs8hd_decap_4
XFILLER_9_181 vpwr vgnd scs8hd_fill_2
XFILLER_28_258 vgnd vpwr scs8hd_decap_12
XFILLER_11_103 vgnd vpwr scs8hd_decap_6
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_12.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_19_258 vpwr vgnd scs8hd_fill_2
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _130_/B vgnd vpwr scs8hd_diode_2
X_228_ _228_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
X_159_ _162_/A _159_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_217 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_31 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vgnd vpwr scs8hd_decap_4
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vgnd vpwr scs8hd_decap_4
XFILLER_3_110 vgnd vpwr scs8hd_decap_8
XANTENNA__104__D _168_/A vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _152_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_242 vpwr vgnd scs8hd_fill_2
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA__115__C _126_/C vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_139 vgnd vpwr scs8hd_decap_8
XFILLER_39_117 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _126_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vgnd vpwr scs8hd_fill_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_98 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_189 vpwr vgnd scs8hd_fill_2
XFILLER_32_167 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_134 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _126_/C vgnd vpwr scs8hd_diode_2
XFILLER_28_6 vgnd vpwr scs8hd_decap_12
XFILLER_9_193 vgnd vpwr scs8hd_decap_4
XFILLER_36_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_119 vgnd vpwr scs8hd_decap_3
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
X_227_ _227_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XANTENNA__118__C _126_/C vgnd vpwr scs8hd_diode_2
X_158_ _161_/A _159_/B _158_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_163 vgnd vpwr scs8hd_decap_3
XFILLER_10_192 vgnd vpwr scs8hd_decap_4
XANTENNA__134__B _130_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_240 vpwr vgnd scs8hd_fill_2
XFILLER_25_229 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_30_243 vgnd vpwr scs8hd_decap_3
XANTENNA__145__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _174_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_254 vpwr vgnd scs8hd_fill_2
XFILLER_12_265 vgnd vpwr scs8hd_decap_8
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA__115__D _168_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_2.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_140 vgnd vpwr scs8hd_decap_4
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_250 vpwr vgnd scs8hd_fill_2
XANTENNA__142__B _140_/X vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _126_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_261 vgnd vpwr scs8hd_decap_12
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_253 vpwr vgnd scs8hd_fill_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_143 vpwr vgnd scs8hd_fill_2
XFILLER_32_146 vgnd vpwr scs8hd_decap_4
XANTENNA__153__A _130_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _178_/Y mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
X_243_ _243_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_14_168 vpwr vgnd scs8hd_fill_2
XFILLER_14_179 vpwr vgnd scs8hd_fill_2
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__D _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_216 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_149 vgnd vpwr scs8hd_decap_4
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_205 vgnd vpwr scs8hd_fill_1
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_226_ _226_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__118__D _171_/A vgnd vpwr scs8hd_diode_2
X_157_ _130_/A address[2] _153_/C _149_/D _159_/B vgnd vpwr scs8hd_or4_4
XANTENNA__134__C _130_/C vgnd vpwr scs8hd_diode_2
XFILLER_40_6 vgnd vpwr scs8hd_decap_12
XANTENNA__150__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_208 vgnd vpwr scs8hd_decap_3
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_178 vgnd vpwr scs8hd_decap_4
XFILLER_30_200 vgnd vpwr scs8hd_decap_12
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_233 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_211 vgnd vpwr scs8hd_fill_1
Xmux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _182_/Y mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_248 vpwr vgnd scs8hd_fill_2
XFILLER_8_259 vgnd vpwr scs8hd_decap_12
XFILLER_5_59 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_229 vpwr vgnd scs8hd_fill_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_39_10 vpwr vgnd scs8hd_fill_2
Xmux_top_track_12.tap_buf4_0_.scs8hd_inv_1 mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_141 vgnd vpwr scs8hd_decap_8
XANTENNA__126__D _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_273 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_188 vpwr vgnd scs8hd_fill_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_136 vgnd vpwr scs8hd_decap_4
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_242_ _242_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__148__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_117 vpwr vgnd scs8hd_fill_2
XFILLER_20_128 vpwr vgnd scs8hd_fill_2
XANTENNA__164__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_173 vpwr vgnd scs8hd_fill_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_8
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_22_68 vgnd vpwr scs8hd_decap_12
XFILLER_19_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__134__D _171_/A vgnd vpwr scs8hd_diode_2
X_156_ _162_/A _154_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__159__A _162_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_242 vpwr vgnd scs8hd_fill_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_146 vgnd vpwr scs8hd_fill_1
XANTENNA__161__B _162_/B vgnd vpwr scs8hd_diode_2
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
X_139_ _160_/C _153_/C vgnd vpwr scs8hd_buf_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_212 vpwr vgnd scs8hd_fill_2
XFILLER_21_245 vgnd vpwr scs8hd_decap_3
XFILLER_21_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_205 vgnd vpwr scs8hd_decap_8
XFILLER_8_227 vgnd vpwr scs8hd_decap_4
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _154_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_186 vpwr vgnd scs8hd_fill_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_197 vpwr vgnd scs8hd_fill_2
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_164 vpwr vgnd scs8hd_fill_2
XFILLER_35_167 vpwr vgnd scs8hd_fill_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_4
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _166_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_189 vgnd vpwr scs8hd_fill_1
XFILLER_26_167 vgnd vpwr scs8hd_decap_4
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XFILLER_17_156 vpwr vgnd scs8hd_fill_2
XFILLER_40_170 vgnd vpwr scs8hd_decap_4
XANTENNA__153__C _153_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _198_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_115 vgnd vpwr scs8hd_decap_3
X_241_ _241_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_229 vgnd vpwr scs8hd_decap_3
XANTENNA__164__B _164_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_152 vpwr vgnd scs8hd_fill_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
XFILLER_12_80 vpwr vgnd scs8hd_fill_2
X_155_ address[0] _162_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_7 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_265 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_46 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_158 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_221 vpwr vgnd scs8hd_fill_2
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_224 vpwr vgnd scs8hd_fill_2
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_265 vpwr vgnd scs8hd_fill_2
X_138_ address[4] _138_/B _160_/C vgnd vpwr scs8hd_nand2_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_70 vgnd vpwr scs8hd_decap_3
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
Xmem_right_track_12.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_165 vgnd vpwr scs8hd_decap_8
XFILLER_38_154 vgnd vpwr scs8hd_decap_8
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_209 vgnd vpwr scs8hd_decap_12
XFILLER_29_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _206_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_6
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _172_/A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_113 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_1_245 vgnd vpwr scs8hd_decap_8
XFILLER_17_102 vgnd vpwr scs8hd_fill_1
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XFILLER_40_193 vgnd vpwr scs8hd_decap_4
XANTENNA__153__D _160_/D vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_138 vgnd vpwr scs8hd_decap_4
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
X_171_ _171_/A _168_/B _162_/A _171_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_274 vgnd vpwr scs8hd_fill_1
XFILLER_36_241 vgnd vpwr scs8hd_decap_4
Xmux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _176_/Y mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_130 vgnd vpwr scs8hd_decap_8
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
XFILLER_10_196 vgnd vpwr scs8hd_fill_1
X_154_ _161_/A _154_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_233 vgnd vpwr scs8hd_decap_4
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_decap_3
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_8.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
X_137_ address[5] _138_/B vgnd vpwr scs8hd_inv_8
XFILLER_2_181 vgnd vpwr scs8hd_decap_12
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_203 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _152_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_258 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr scs8hd_diode_2
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_38_144 vgnd vpwr scs8hd_fill_1
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_136 vgnd vpwr scs8hd_decap_12
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vgnd vpwr scs8hd_decap_4
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
X_170_ _171_/A _168_/B _161_/A _170_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_121 vgnd vpwr scs8hd_fill_1
XFILLER_9_165 vgnd vpwr scs8hd_decap_6
XFILLER_13_194 vpwr vgnd scs8hd_fill_2
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_231 vgnd vpwr scs8hd_fill_1
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_175 vpwr vgnd scs8hd_fill_2
X_153_ _130_/A address[2] _153_/C _160_/D _154_/B vgnd vpwr scs8hd_or4_4
XFILLER_6_168 vpwr vgnd scs8hd_fill_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_231 vgnd vpwr scs8hd_fill_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_3
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_24_223 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
XFILLER_15_201 vpwr vgnd scs8hd_fill_2
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_259 vgnd vpwr scs8hd_decap_12
XFILLER_30_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
X_136_ _151_/A _136_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_193 vgnd vpwr scs8hd_decap_12
XFILLER_0_30 vgnd vpwr scs8hd_fill_1
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_21_259 vpwr vgnd scs8hd_fill_2
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XFILLER_12_237 vgnd vpwr scs8hd_decap_8
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_263 vgnd vpwr scs8hd_decap_12
X_119_ _096_/X _118_/X _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_12.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_14 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_148 vgnd vpwr scs8hd_decap_4
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XFILLER_40_151 vpwr vgnd scs8hd_fill_2
XFILLER_31_140 vgnd vpwr scs8hd_decap_6
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_4
XFILLER_31_173 vgnd vpwr scs8hd_decap_3
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_107 vgnd vpwr scs8hd_decap_8
XFILLER_22_140 vpwr vgnd scs8hd_fill_2
XFILLER_22_195 vgnd vpwr scs8hd_decap_8
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_144 vgnd vpwr scs8hd_decap_6
XFILLER_9_177 vpwr vgnd scs8hd_fill_2
XFILLER_9_199 vpwr vgnd scs8hd_fill_2
XFILLER_13_162 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vgnd vpwr scs8hd_fill_1
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_210 vpwr vgnd scs8hd_fill_2
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
X_152_ _152_/A _161_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _196_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_210 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_246 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_135_ _129_/X _136_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_62 vgnd vpwr scs8hd_decap_8
XFILLER_21_216 vpwr vgnd scs8hd_fill_2
XFILLER_21_238 vpwr vgnd scs8hd_fill_2
XFILLER_12_227 vgnd vpwr scs8hd_fill_1
XFILLER_20_260 vgnd vpwr scs8hd_decap_12
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_11_260 vgnd vpwr scs8hd_decap_4
XFILLER_11_271 vgnd vpwr scs8hd_decap_6
XFILLER_7_275 vpwr vgnd scs8hd_fill_2
X_118_ _115_/A _130_/B _126_/C _171_/A _118_/X vgnd vpwr scs8hd_or4_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
Xmem_right_track_4.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_26 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_168 vpwr vgnd scs8hd_fill_2
XFILLER_26_105 vgnd vpwr scs8hd_decap_8
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_34_171 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_152 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _204_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_163 vgnd vpwr scs8hd_decap_3
XFILLER_22_174 vgnd vpwr scs8hd_decap_8
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_101 vgnd vpwr scs8hd_fill_1
XFILLER_9_112 vgnd vpwr scs8hd_decap_3
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XFILLER_13_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_111 vgnd vpwr scs8hd_decap_8
XFILLER_10_188 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vgnd vpwr scs8hd_decap_8
X_151_ _151_/A _150_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_214 vpwr vgnd scs8hd_fill_2
XFILLER_5_170 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_203 vgnd vpwr scs8hd_fill_1
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_228 vgnd vpwr scs8hd_decap_4
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _174_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_15_258 vpwr vgnd scs8hd_fill_2
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
X_134_ _130_/A _130_/B _130_/C _171_/A _136_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_151 vpwr vgnd scs8hd_fill_2
XFILLER_0_10 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_272 vgnd vpwr scs8hd_decap_3
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
X_117_ _128_/A _115_/X _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_147 vgnd vpwr scs8hd_decap_6
XFILLER_38_125 vgnd vpwr scs8hd_fill_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_38 vgnd vpwr scs8hd_decap_12
XFILLER_37_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_183 vgnd vpwr scs8hd_decap_3
XFILLER_40_131 vgnd vpwr scs8hd_decap_12
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_150 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_161 vgnd vpwr scs8hd_decap_3
XFILLER_16_183 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vpwr vgnd scs8hd_fill_2
XFILLER_27_234 vgnd vpwr scs8hd_decap_8
XFILLER_42_259 vgnd vpwr scs8hd_decap_12
XFILLER_10_101 vgnd vpwr scs8hd_fill_1
X_150_ _129_/X _150_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_149 vgnd vpwr scs8hd_decap_4
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_167 vgnd vpwr scs8hd_decap_8
XFILLER_33_259 vgnd vpwr scs8hd_decap_4
XFILLER_33_237 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_234 vgnd vpwr scs8hd_decap_12
XFILLER_18_256 vgnd vpwr scs8hd_decap_8
XFILLER_18_267 vgnd vpwr scs8hd_decap_8
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_8
XFILLER_24_259 vpwr vgnd scs8hd_fill_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
X_133_ _151_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_22 vgnd vpwr scs8hd_decap_8
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _115_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_229 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XFILLER_28_18 vgnd vpwr scs8hd_decap_12
XFILLER_12_207 vgnd vpwr scs8hd_decap_4
X_116_ _096_/X _115_/X _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_137 vpwr vgnd scs8hd_fill_2
XFILLER_4_247 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_143 vgnd vpwr scs8hd_decap_8
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_25_140 vgnd vpwr scs8hd_decap_8
XFILLER_25_173 vpwr vgnd scs8hd_fill_2
XFILLER_25_184 vgnd vpwr scs8hd_decap_3
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XANTENNA__102__B _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_132 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vgnd vpwr scs8hd_decap_6
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_13_198 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_224 vpwr vgnd scs8hd_fill_2
XFILLER_36_202 vgnd vpwr scs8hd_fill_1
XFILLER_3_55 vgnd vpwr scs8hd_decap_6
XFILLER_42_249 vgnd vpwr scs8hd_decap_6
XFILLER_6_117 vgnd vpwr scs8hd_decap_8
XFILLER_6_128 vgnd vpwr scs8hd_decap_8
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_246 vgnd vpwr scs8hd_fill_1
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_227 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_205 vgnd vpwr scs8hd_decap_3
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
X_132_ address[0] _151_/A vgnd vpwr scs8hd_buf_1
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XANTENNA__110__B _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_10 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _194_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_219 vgnd vpwr scs8hd_decap_8
XFILLER_11_230 vpwr vgnd scs8hd_fill_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_3
XANTENNA__105__B _104_/X vgnd vpwr scs8hd_diode_2
X_115_ _115_/A _130_/B _126_/C _168_/A _115_/X vgnd vpwr scs8hd_or4_4
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_193 vgnd vpwr scs8hd_decap_3
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_28_182 vpwr vgnd scs8hd_fill_2
XFILLER_28_171 vgnd vpwr scs8hd_decap_8
XANTENNA__116__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_26_119 vgnd vpwr scs8hd_decap_8
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_160 vpwr vgnd scs8hd_fill_2
XFILLER_19_171 vpwr vgnd scs8hd_fill_2
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _198_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_177 vgnd vpwr scs8hd_decap_8
XFILLER_15_31 vgnd vpwr scs8hd_decap_12
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_25_196 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_262 vgnd vpwr scs8hd_decap_12
XFILLER_16_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_188 vgnd vpwr scs8hd_fill_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

